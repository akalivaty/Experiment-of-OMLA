//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  XOR2_X1   g000(.A(KEYINPUT71), .B(G217), .Z(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  OR3_X1    g004(.A1(new_n190), .A2(KEYINPUT72), .A3(G128), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT72), .B1(new_n190), .B2(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(G128), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT24), .B(G110), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n197), .B(G119), .C1(KEYINPUT73), .C2(KEYINPUT23), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n193), .A2(KEYINPUT23), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT73), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n200), .B1(new_n190), .B2(G128), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n198), .B1(new_n199), .B2(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n196), .B1(G110), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT16), .ZN(new_n205));
  INV_X1    g019(.A(G140), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G125), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G140), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT74), .ZN(new_n210));
  OR3_X1    g024(.A1(new_n208), .A2(KEYINPUT74), .A3(G140), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n205), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n207), .A2(KEYINPUT16), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n204), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n213), .ZN(new_n215));
  NOR3_X1   g029(.A1(new_n208), .A2(KEYINPUT74), .A3(G140), .ZN(new_n216));
  XNOR2_X1  g030(.A(G125), .B(G140), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(KEYINPUT74), .ZN(new_n218));
  OAI211_X1 g032(.A(G146), .B(new_n215), .C1(new_n218), .C2(new_n205), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT75), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n214), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n210), .A2(new_n211), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n213), .B1(new_n222), .B2(KEYINPUT16), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT75), .B1(new_n223), .B2(G146), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n203), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n194), .A2(new_n195), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n226), .B1(new_n202), .B2(G110), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n217), .A2(new_n204), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n219), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G953), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(G221), .A3(G234), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n232), .B(KEYINPUT22), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n233), .B(G137), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n225), .A2(new_n229), .A3(new_n234), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT25), .ZN(new_n238));
  OR2_X1    g052(.A1(new_n238), .A2(KEYINPUT76), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(KEYINPUT76), .ZN(new_n240));
  AOI21_X1  g054(.A(G902), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n236), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n225), .A2(new_n229), .A3(new_n234), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n234), .B1(new_n225), .B2(new_n229), .ZN(new_n244));
  NOR3_X1   g058(.A1(new_n243), .A2(new_n244), .A3(G902), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n189), .B(new_n242), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n189), .A2(G902), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT77), .ZN(new_n249));
  NOR3_X1   g063(.A1(new_n243), .A2(new_n244), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(KEYINPUT77), .B1(new_n236), .B2(new_n237), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT78), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n247), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n253), .B1(new_n247), .B2(new_n252), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT9), .B(G234), .ZN(new_n257));
  OAI21_X1  g071(.A(G221), .B1(new_n257), .B2(G902), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G469), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(new_n188), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT11), .ZN(new_n262));
  INV_X1    g076(.A(G134), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n262), .B1(new_n263), .B2(G137), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(G137), .ZN(new_n265));
  INV_X1    g079(.A(G137), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT11), .A3(G134), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G131), .ZN(new_n269));
  INV_X1    g083(.A(G131), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n264), .A2(new_n267), .A3(new_n270), .A4(new_n265), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT10), .ZN(new_n273));
  INV_X1    g087(.A(G104), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT3), .B1(new_n274), .B2(G107), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT3), .ZN(new_n276));
  INV_X1    g090(.A(G107), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n277), .A3(G104), .ZN(new_n278));
  INV_X1    g092(.A(G101), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(G107), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n275), .A2(new_n278), .A3(new_n279), .A4(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n274), .A2(G107), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n277), .A2(G104), .ZN(new_n283));
  OAI21_X1  g097(.A(G101), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT65), .ZN(new_n287));
  XNOR2_X1  g101(.A(G143), .B(G146), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n204), .A2(G143), .ZN(new_n291));
  INV_X1    g105(.A(G143), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G146), .ZN(new_n293));
  AND4_X1   g107(.A1(new_n287), .A2(new_n289), .A3(new_n291), .A4(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(KEYINPUT1), .B1(new_n292), .B2(G146), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n197), .B1(new_n296), .B2(KEYINPUT81), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT81), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n291), .A2(new_n298), .A3(KEYINPUT1), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n288), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n286), .B1(new_n295), .B2(new_n300), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n296), .A2(G128), .B1(new_n291), .B2(new_n293), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n289), .A2(new_n291), .A3(new_n293), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT65), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n288), .A2(new_n287), .A3(new_n289), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n302), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(new_n273), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n273), .A2(new_n301), .B1(new_n307), .B2(new_n286), .ZN(new_n308));
  AND2_X1   g122(.A1(KEYINPUT0), .A2(G128), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n291), .A2(new_n293), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT0), .B(G128), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n310), .B1(new_n288), .B2(new_n311), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n281), .A2(KEYINPUT4), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n275), .A2(new_n278), .A3(new_n280), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G101), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n312), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT4), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n314), .A2(new_n317), .A3(G101), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT80), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT80), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n314), .A2(new_n320), .A3(new_n317), .A4(G101), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n272), .B1(new_n308), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n297), .A2(new_n299), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n291), .A2(new_n293), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n325), .A2(new_n326), .B1(new_n304), .B2(new_n305), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n273), .B1(new_n327), .B2(new_n285), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n296), .A2(G128), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n326), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n330), .B1(new_n290), .B2(new_n294), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT10), .A3(new_n286), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n323), .A2(new_n328), .A3(new_n272), .A4(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(G110), .B(G140), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(KEYINPUT79), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n231), .A2(G227), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n324), .A2(new_n334), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT12), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n304), .A2(new_n305), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(new_n330), .A3(new_n285), .ZN(new_n343));
  AOI211_X1 g157(.A(new_n341), .B(new_n272), .C1(new_n301), .C2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n343), .B1(new_n327), .B2(new_n285), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n269), .A2(new_n271), .ZN(new_n346));
  AOI21_X1  g160(.A(KEYINPUT12), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n333), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT82), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT82), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n350), .B(new_n333), .C1(new_n344), .C2(new_n347), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n340), .B1(new_n352), .B2(new_n339), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n261), .B1(new_n353), .B2(G469), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT83), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n339), .B1(new_n324), .B2(new_n334), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n338), .B(new_n333), .C1(new_n344), .C2(new_n347), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n357), .A2(new_n355), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n260), .B(new_n188), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n259), .B1(new_n354), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n312), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n346), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT64), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n364), .B1(new_n266), .B2(G134), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n266), .A2(G134), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n263), .A2(KEYINPUT64), .A3(G137), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G131), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n271), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n363), .B(KEYINPUT30), .C1(new_n306), .C2(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(G116), .A2(G119), .ZN(new_n372));
  NOR2_X1   g186(.A1(G116), .A2(G119), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT67), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OR2_X1    g190(.A1(KEYINPUT2), .A2(G113), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT2), .A2(G113), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n374), .A3(new_n375), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n371), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT66), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n369), .A2(new_n271), .ZN(new_n386));
  AOI22_X1  g200(.A1(new_n386), .A2(new_n331), .B1(new_n346), .B2(new_n362), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n385), .B1(new_n387), .B2(KEYINPUT30), .ZN(new_n388));
  OAI22_X1  g202(.A1(new_n272), .A2(new_n312), .B1(new_n306), .B2(new_n370), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT30), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(KEYINPUT66), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n384), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(G237), .A2(G953), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G210), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT27), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n394), .B(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT26), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n394), .B(KEYINPUT27), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(KEYINPUT26), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n279), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(KEYINPUT26), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n396), .A2(new_n397), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(G101), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n383), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n387), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT31), .B1(new_n392), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n401), .A2(new_n404), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n383), .B1(new_n389), .B2(KEYINPUT68), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT68), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n387), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT28), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT28), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n389), .A2(new_n383), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n415), .B1(new_n407), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n410), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n406), .B1(new_n387), .B2(KEYINPUT30), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n387), .A2(new_n385), .A3(KEYINPUT30), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT66), .B1(new_n389), .B2(new_n390), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT31), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n389), .A2(new_n383), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n410), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n422), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n409), .A2(new_n418), .A3(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(G472), .A2(G902), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(KEYINPUT32), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT70), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n410), .B1(new_n392), .B2(new_n424), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT29), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n406), .B1(new_n387), .B2(new_n412), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n389), .A2(KEYINPUT68), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n415), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n386), .A2(new_n331), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n406), .B1(new_n437), .B2(new_n363), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT28), .B1(new_n424), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n436), .A2(new_n405), .A3(new_n439), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n432), .A2(new_n433), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n188), .B1(new_n440), .B2(new_n433), .ZN(new_n442));
  OAI21_X1  g256(.A(G472), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n427), .A2(new_n428), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT69), .B(KEYINPUT32), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n427), .A2(KEYINPUT70), .A3(KEYINPUT32), .A4(new_n428), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n431), .A2(new_n443), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(G214), .B1(G237), .B2(G902), .ZN(new_n449));
  XNOR2_X1  g263(.A(G110), .B(G122), .ZN(new_n450));
  XOR2_X1   g264(.A(new_n450), .B(KEYINPUT8), .Z(new_n451));
  OAI211_X1 g265(.A(new_n377), .B(new_n378), .C1(new_n372), .C2(new_n373), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT5), .ZN(new_n453));
  INV_X1    g267(.A(new_n373), .ZN(new_n454));
  NAND2_X1  g268(.A1(G116), .A2(G119), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(new_n190), .A3(G116), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G113), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n452), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n285), .ZN(new_n460));
  OAI211_X1 g274(.A(G113), .B(new_n457), .C1(new_n374), .C2(new_n453), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n461), .A2(new_n281), .A3(new_n284), .A4(new_n452), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n451), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT84), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(new_n312), .B2(G125), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n342), .A2(new_n208), .A3(new_n330), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n312), .A2(new_n464), .A3(G125), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G224), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(G953), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT85), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n471), .B1(new_n472), .B2(KEYINPUT7), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n473), .B1(new_n472), .B2(KEYINPUT7), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n463), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n319), .A2(new_n321), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n315), .A2(KEYINPUT4), .A3(new_n281), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n383), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n450), .B(new_n462), .C1(new_n476), .C2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n468), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(new_n465), .ZN(new_n481));
  INV_X1    g295(.A(new_n471), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n481), .A2(KEYINPUT7), .A3(new_n482), .A4(new_n467), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n475), .A2(new_n479), .A3(new_n483), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n484), .A2(new_n188), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n459), .A2(new_n285), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n313), .A2(new_n315), .B1(new_n381), .B2(new_n382), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n487), .B1(new_n488), .B2(new_n322), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n486), .B1(new_n489), .B2(new_n450), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n462), .B1(new_n476), .B2(new_n478), .ZN(new_n491));
  INV_X1    g305(.A(new_n450), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n469), .B(new_n471), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n491), .A2(new_n486), .A3(new_n492), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(G210), .B1(G237), .B2(G902), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n485), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n498), .B1(new_n485), .B2(new_n497), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n449), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT20), .ZN(new_n502));
  XNOR2_X1  g316(.A(G113), .B(G122), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(new_n274), .ZN(new_n504));
  AOI21_X1  g318(.A(G143), .B1(new_n393), .B2(G214), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n393), .A2(G143), .A3(G214), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(KEYINPUT18), .A3(G131), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n228), .B1(new_n222), .B2(new_n204), .ZN(new_n510));
  NAND2_X1  g324(.A1(KEYINPUT18), .A2(G131), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n506), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n219), .A2(new_n220), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n223), .A2(KEYINPUT75), .A3(G146), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n515), .A3(new_n214), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n508), .A2(KEYINPUT17), .A3(G131), .ZN(new_n517));
  INV_X1    g331(.A(new_n507), .ZN(new_n518));
  OAI21_X1  g332(.A(G131), .B1(new_n518), .B2(new_n505), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n506), .A2(new_n270), .A3(new_n507), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n517), .B1(new_n521), .B2(KEYINPUT17), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n504), .B(new_n513), .C1(new_n516), .C2(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n217), .A2(KEYINPUT19), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n524), .B1(new_n222), .B2(KEYINPUT19), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n521), .B(new_n219), .C1(new_n525), .C2(G146), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n513), .ZN(new_n527));
  INV_X1    g341(.A(new_n504), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n523), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(G475), .A2(G902), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n502), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n531), .ZN(new_n533));
  AOI211_X1 g347(.A(KEYINPUT20), .B(new_n533), .C1(new_n523), .C2(new_n529), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n513), .B1(new_n516), .B2(new_n522), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n528), .ZN(new_n536));
  AOI21_X1  g350(.A(G902), .B1(new_n536), .B2(new_n523), .ZN(new_n537));
  INV_X1    g351(.A(G475), .ZN(new_n538));
  OAI22_X1  g352(.A1(new_n532), .A2(new_n534), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G478), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(KEYINPUT15), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT86), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n292), .A2(G128), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n292), .A2(G128), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT13), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n543), .B(new_n544), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n197), .A2(G143), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n197), .A2(G143), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n548), .B1(KEYINPUT13), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT86), .B1(new_n544), .B2(new_n546), .ZN(new_n551));
  OAI211_X1 g365(.A(G134), .B(new_n547), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT87), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n543), .B1(new_n548), .B2(KEYINPUT13), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n263), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(KEYINPUT87), .A3(new_n547), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n548), .A2(new_n545), .A3(G134), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G116), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n562), .A2(G122), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(G122), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n564), .A3(new_n277), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n277), .B1(new_n563), .B2(new_n564), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n561), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n559), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n263), .B1(new_n544), .B2(new_n549), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n565), .B1(new_n560), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n564), .A2(KEYINPUT88), .A3(KEYINPUT14), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT88), .B1(new_n564), .B2(KEYINPUT14), .ZN(new_n575));
  OAI221_X1 g389(.A(new_n563), .B1(KEYINPUT14), .B2(new_n564), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n572), .B1(new_n576), .B2(G107), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n187), .A2(G953), .A3(new_n257), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n570), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n579), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n568), .B1(new_n554), .B2(new_n558), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n581), .B1(new_n582), .B2(new_n577), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n542), .B1(new_n584), .B2(new_n188), .ZN(new_n585));
  AOI211_X1 g399(.A(G902), .B(new_n541), .C1(new_n580), .C2(new_n583), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(G952), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n588), .A2(KEYINPUT89), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(KEYINPUT89), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n231), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(G234), .B2(G237), .ZN(new_n592));
  NAND2_X1  g406(.A1(G234), .A2(G237), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(G902), .A3(G953), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(KEYINPUT90), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT21), .B(G898), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n587), .A2(new_n598), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n501), .A2(new_n539), .A3(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n256), .A2(new_n361), .A3(new_n448), .A4(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G101), .ZN(G3));
  OAI211_X1 g416(.A(new_n449), .B(new_n598), .C1(new_n499), .C2(new_n500), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT91), .B1(new_n582), .B2(new_n577), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT33), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n584), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n580), .A2(new_n583), .A3(new_n604), .A4(KEYINPUT33), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n606), .A2(G478), .A3(new_n607), .A4(new_n188), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n584), .A2(new_n188), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n540), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n539), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n603), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n427), .A2(new_n188), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n614), .A2(G472), .B1(new_n428), .B2(new_n427), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n361), .A2(new_n256), .A3(new_n613), .A4(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT34), .B(G104), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  NAND2_X1  g432(.A1(new_n530), .A2(new_n531), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT20), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n530), .A2(new_n502), .A3(new_n531), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(KEYINPUT92), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT92), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n532), .B2(new_n534), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n585), .A2(new_n586), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n536), .A2(new_n523), .ZN(new_n626));
  OAI21_X1  g440(.A(G475), .B1(new_n626), .B2(G902), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n622), .A2(new_n624), .A3(new_n625), .A4(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n603), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n361), .A2(new_n256), .A3(new_n629), .A4(new_n615), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT35), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NOR2_X1   g448(.A1(new_n235), .A2(KEYINPUT36), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n230), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n248), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n247), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n361), .A2(new_n600), .A3(new_n615), .A4(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT37), .B(G110), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G12));
  INV_X1    g455(.A(G900), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n595), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n592), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n628), .A2(new_n501), .A3(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n645), .A2(new_n361), .A3(new_n448), .A4(new_n638), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G128), .ZN(G30));
  XOR2_X1   g461(.A(new_n644), .B(KEYINPUT39), .Z(new_n648));
  NAND2_X1  g462(.A1(new_n361), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT40), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n485), .A2(new_n497), .ZN(new_n652));
  INV_X1    g466(.A(new_n498), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n485), .A2(new_n497), .A3(new_n498), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT38), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n539), .A2(new_n625), .ZN(new_n658));
  INV_X1    g472(.A(new_n449), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n638), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n392), .A2(new_n424), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n410), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n410), .A2(new_n407), .A3(new_n416), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n188), .ZN(new_n665));
  OAI21_X1  g479(.A(G472), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n431), .A2(new_n446), .A3(new_n447), .A4(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT95), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n661), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n651), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(KEYINPUT96), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT96), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n651), .A2(new_n674), .A3(new_n671), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n292), .ZN(G45));
  OAI211_X1 g491(.A(new_n539), .B(new_n611), .C1(new_n592), .C2(new_n643), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n501), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n361), .A2(new_n448), .A3(new_n638), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  OAI21_X1  g495(.A(new_n188), .B1(new_n358), .B2(new_n359), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(G469), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(new_n258), .A3(new_n360), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n685), .A2(new_n448), .A3(new_n256), .A4(new_n613), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT41), .B(G113), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT97), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n686), .B(new_n688), .ZN(G15));
  NAND4_X1  g503(.A1(new_n685), .A2(new_n448), .A3(new_n256), .A4(new_n629), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT98), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n562), .ZN(G18));
  AOI21_X1  g506(.A(new_n659), .B1(new_n654), .B2(new_n655), .ZN(new_n693));
  AND4_X1   g507(.A1(new_n258), .A2(new_n683), .A3(new_n693), .A4(new_n360), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n599), .A2(new_n539), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n694), .A2(new_n448), .A3(new_n695), .A4(new_n638), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  AND2_X1   g511(.A1(new_n683), .A2(new_n360), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n501), .A2(new_n658), .A3(new_n597), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(new_n699), .A3(new_n258), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n247), .A2(new_n252), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n614), .A2(G472), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n428), .B(KEYINPUT99), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n427), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT100), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n427), .A2(KEYINPUT100), .A3(new_n704), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n702), .A2(new_n703), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(KEYINPUT101), .B1(new_n700), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n620), .A2(new_n621), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n587), .B1(new_n711), .B2(new_n627), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n712), .A2(new_n656), .A3(new_n449), .A4(new_n598), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n684), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n709), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT101), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n710), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G122), .ZN(G24));
  NAND4_X1  g533(.A1(new_n703), .A2(new_n707), .A3(new_n638), .A4(new_n708), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n678), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n694), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G125), .ZN(G27));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n678), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n443), .A2(new_n429), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT32), .B1(new_n427), .B2(new_n428), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n725), .B(new_n702), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n345), .A2(new_n346), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n341), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n345), .A2(KEYINPUT12), .A3(new_n346), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n350), .B1(new_n732), .B2(new_n333), .ZN(new_n733));
  INV_X1    g547(.A(new_n351), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n339), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n340), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(G469), .A3(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n261), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n360), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n499), .A2(new_n500), .A3(new_n659), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n258), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n728), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n361), .A2(new_n448), .A3(new_n256), .A4(new_n740), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n724), .B1(new_n744), .B2(new_n678), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G131), .ZN(G33));
  AND2_X1   g561(.A1(new_n448), .A2(new_n256), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n628), .A2(new_n644), .ZN(new_n749));
  INV_X1    g563(.A(new_n741), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  INV_X1    g566(.A(KEYINPUT46), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n261), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n735), .A2(KEYINPUT45), .A3(new_n736), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n338), .B1(new_n349), .B2(new_n351), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n757), .B1(new_n758), .B2(new_n340), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n756), .A2(new_n759), .A3(G469), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT102), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n260), .B1(new_n353), .B2(KEYINPUT45), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(KEYINPUT102), .A3(new_n759), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n755), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n360), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT103), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT102), .B1(new_n763), .B2(new_n759), .ZN(new_n768));
  AND4_X1   g582(.A1(KEYINPUT102), .A2(new_n756), .A3(new_n759), .A4(G469), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n754), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT103), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(new_n771), .A3(new_n360), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n738), .B1(new_n768), .B2(new_n769), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n753), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n767), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n258), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n615), .ZN(new_n778));
  INV_X1    g592(.A(new_n611), .ZN(new_n779));
  OAI21_X1  g593(.A(KEYINPUT43), .B1(new_n779), .B2(new_n539), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n539), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT43), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AND4_X1   g597(.A1(new_n778), .A2(new_n780), .A3(new_n638), .A4(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n784), .A2(KEYINPUT44), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(KEYINPUT44), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n654), .A2(new_n449), .A3(new_n655), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n777), .A2(new_n648), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G137), .ZN(G39));
  NAND2_X1  g604(.A1(new_n776), .A2(KEYINPUT47), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT47), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n775), .A2(new_n792), .A3(new_n258), .ZN(new_n793));
  NOR4_X1   g607(.A1(new_n448), .A2(new_n256), .A3(new_n678), .A4(new_n787), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n791), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G140), .ZN(G42));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n361), .A2(new_n448), .A3(new_n638), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n622), .A2(new_n624), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n585), .A2(new_n586), .A3(new_n644), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n800), .A2(new_n627), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n740), .A2(new_n799), .A3(KEYINPUT109), .A4(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT109), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n622), .A2(new_n624), .A3(new_n800), .A4(new_n627), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n803), .B1(new_n804), .B2(new_n787), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n798), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT110), .B1(new_n721), .B2(new_n750), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT110), .ZN(new_n809));
  NOR4_X1   g623(.A1(new_n741), .A2(new_n720), .A3(new_n809), .A4(new_n678), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n807), .B(new_n751), .C1(new_n808), .C2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n678), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n748), .A2(new_n812), .A3(new_n750), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n742), .B1(new_n813), .B2(new_n724), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n601), .A2(new_n616), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT107), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT107), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n601), .A2(new_n616), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT108), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n701), .A2(KEYINPUT78), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n247), .A2(new_n252), .A3(new_n253), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n615), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n739), .A2(new_n258), .ZN(new_n824));
  INV_X1    g638(.A(new_n539), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n693), .A2(new_n825), .A3(new_n598), .A4(new_n625), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n823), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n693), .A2(new_n695), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n703), .A2(new_n444), .A3(new_n638), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n824), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n820), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n825), .A2(new_n625), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n603), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n361), .A2(new_n256), .A3(new_n833), .A4(new_n615), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(new_n639), .A3(KEYINPUT108), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n817), .A2(new_n819), .B1(new_n831), .B2(new_n835), .ZN(new_n836));
  NOR4_X1   g650(.A1(new_n709), .A2(new_n684), .A3(new_n713), .A4(KEYINPUT101), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n716), .B1(new_n714), .B2(new_n715), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n696), .A2(new_n686), .A3(new_n690), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT106), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT106), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n748), .B(new_n685), .C1(new_n613), .C2(new_n629), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n718), .A2(new_n842), .A3(new_n696), .A4(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n815), .A2(new_n836), .A3(new_n841), .A4(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n501), .A2(new_n658), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n644), .B(KEYINPUT111), .Z(new_n847));
  NOR2_X1   g661(.A1(new_n638), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n361), .A2(new_n667), .A3(new_n846), .A4(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n722), .A2(new_n680), .A3(new_n646), .A4(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT52), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n797), .B1(new_n845), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n721), .A2(new_n750), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n809), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n721), .A2(new_n750), .A3(KEYINPUT110), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n744), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n858), .A2(new_n749), .B1(new_n798), .B2(new_n806), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n746), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n819), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n818), .B1(new_n601), .B2(new_n616), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n834), .A2(new_n639), .A3(KEYINPUT108), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT108), .B1(new_n834), .B2(new_n639), .ZN(new_n864));
  OAI22_X1  g678(.A1(new_n861), .A2(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n718), .A2(new_n696), .A3(new_n843), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT112), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n850), .B(KEYINPUT52), .Z(new_n870));
  AOI21_X1  g684(.A(new_n797), .B1(new_n867), .B2(new_n868), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n866), .A2(new_n869), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n852), .A2(new_n853), .A3(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n841), .A2(new_n844), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n866), .A3(new_n870), .A4(KEYINPUT53), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n853), .B1(new_n852), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT113), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n852), .A2(new_n875), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT54), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT113), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n852), .A2(new_n853), .A3(new_n872), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT51), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n783), .A2(new_n592), .A3(new_n780), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n709), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n740), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n791), .A2(new_n793), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n698), .A2(new_n259), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT114), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n886), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n657), .A2(new_n449), .A3(new_n684), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n885), .A2(new_n891), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n892), .A2(KEYINPUT50), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(KEYINPUT50), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n669), .A2(new_n670), .ZN(new_n896));
  AND4_X1   g710(.A1(new_n256), .A2(new_n685), .A3(new_n592), .A4(new_n740), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n896), .A2(new_n825), .A3(new_n897), .A4(new_n779), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n685), .A2(new_n740), .ZN(new_n899));
  OR3_X1    g713(.A1(new_n899), .A2(new_n720), .A3(new_n884), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n895), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n883), .B1(new_n890), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT115), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n775), .A2(new_n792), .A3(new_n258), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n792), .B1(new_n775), .B2(new_n258), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n888), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n886), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(KEYINPUT51), .A3(new_n902), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n899), .A2(new_n884), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n726), .A2(new_n727), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(new_n701), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT48), .Z(new_n916));
  AOI21_X1  g730(.A(new_n591), .B1(new_n885), .B2(new_n694), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n896), .A2(new_n897), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n917), .B1(new_n918), .B2(new_n612), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n904), .A2(new_n905), .A3(new_n911), .A4(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n922));
  INV_X1    g736(.A(new_n901), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n923), .B(KEYINPUT51), .C1(new_n894), .C2(new_n893), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n920), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n889), .B1(new_n906), .B2(new_n907), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n909), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT51), .B1(new_n927), .B2(new_n902), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT115), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n877), .A2(new_n882), .A3(new_n921), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n588), .A2(new_n231), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n683), .A2(new_n360), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(KEYINPUT49), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT105), .Z(new_n935));
  AOI21_X1  g749(.A(new_n657), .B1(KEYINPUT49), .B2(new_n933), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n781), .A2(new_n702), .A3(new_n258), .A4(new_n449), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT104), .Z(new_n938));
  NAND4_X1  g752(.A1(new_n935), .A2(new_n896), .A3(new_n936), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n932), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT116), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n932), .A2(KEYINPUT116), .A3(new_n939), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(G75));
  NOR2_X1   g758(.A1(new_n231), .A2(G952), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n188), .B1(new_n852), .B2(new_n872), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT56), .B1(new_n947), .B2(G210), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n494), .A2(new_n496), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(new_n495), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT55), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n946), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n948), .B2(new_n951), .ZN(G51));
  NAND2_X1  g767(.A1(new_n852), .A2(new_n872), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(new_n853), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n261), .B(KEYINPUT57), .Z(new_n956));
  OAI22_X1  g770(.A1(new_n955), .A2(new_n956), .B1(new_n358), .B2(new_n359), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n947), .A2(new_n762), .A3(new_n764), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n945), .B1(new_n957), .B2(new_n958), .ZN(G54));
  AND3_X1   g773(.A1(new_n947), .A2(KEYINPUT58), .A3(G475), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n530), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n961), .A2(KEYINPUT117), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n961), .A2(KEYINPUT117), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n946), .B1(new_n960), .B2(new_n530), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(G60));
  AND2_X1   g779(.A1(new_n606), .A2(new_n607), .ZN(new_n966));
  NAND2_X1  g780(.A1(G478), .A2(G902), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT59), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n946), .B1(new_n955), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT118), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n877), .A2(new_n882), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n966), .B1(new_n972), .B2(new_n968), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n971), .A2(new_n973), .ZN(G63));
  NAND2_X1  g788(.A1(G217), .A2(G902), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT119), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT60), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n954), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n250), .A2(new_n251), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n954), .A2(new_n636), .A3(new_n977), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n980), .A2(new_n946), .A3(new_n981), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g797(.A(G953), .B1(new_n596), .B2(new_n470), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT120), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n874), .A2(new_n836), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n985), .B1(new_n986), .B2(G953), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n949), .B1(G898), .B2(new_n231), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(G69));
  OAI21_X1  g803(.A(new_n371), .B1(new_n420), .B2(new_n421), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT121), .Z(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(new_n525), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n722), .A2(new_n680), .A3(new_n646), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n673), .A2(new_n675), .A3(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT62), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n673), .A2(KEYINPUT62), .A3(new_n675), .A4(new_n993), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n787), .B1(new_n832), .B2(new_n612), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n748), .A2(new_n361), .A3(new_n648), .A4(new_n999), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n789), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n998), .A2(new_n1001), .A3(new_n795), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n992), .B1(new_n1002), .B2(new_n231), .ZN(new_n1003));
  OR2_X1    g817(.A1(new_n1003), .A2(KEYINPUT122), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(KEYINPUT122), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n777), .A2(new_n648), .A3(new_n846), .A4(new_n914), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n746), .A2(new_n751), .A3(new_n993), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n1006), .A2(new_n789), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(G953), .B1(new_n1008), .B2(new_n795), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n231), .A2(G900), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1010), .B(KEYINPUT123), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n992), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1004), .A2(new_n1005), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n231), .B1(G227), .B2(G900), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1013), .B(new_n1014), .ZN(G72));
  NAND4_X1  g829(.A1(new_n998), .A2(new_n1001), .A3(new_n795), .A4(new_n986), .ZN(new_n1016));
  XOR2_X1   g830(.A(KEYINPUT124), .B(KEYINPUT63), .Z(new_n1017));
  NAND2_X1  g831(.A1(G472), .A2(G902), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(KEYINPUT125), .B1(new_n1020), .B2(new_n663), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT125), .ZN(new_n1022));
  INV_X1    g836(.A(new_n663), .ZN(new_n1023));
  AOI211_X1 g837(.A(new_n1022), .B(new_n1023), .C1(new_n1016), .C2(new_n1019), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(KEYINPUT127), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1008), .A2(new_n986), .A3(new_n795), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(new_n1019), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT126), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1028), .A2(KEYINPUT126), .A3(new_n1019), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n662), .A2(new_n410), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1033), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1031), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  AND3_X1   g849(.A1(new_n1023), .A2(new_n1019), .A3(new_n1033), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n945), .B1(new_n878), .B2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g851(.A1(new_n1026), .A2(new_n1027), .A3(new_n1035), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1039));
  OAI21_X1  g853(.A(KEYINPUT127), .B1(new_n1039), .B2(new_n1025), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1038), .A2(new_n1040), .ZN(G57));
endmodule


