//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937;
  INV_X1    g000(.A(KEYINPUT76), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT3), .B1(new_n188), .B2(G107), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G104), .ZN(new_n192));
  INV_X1    g006(.A(G101), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n188), .A2(G107), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n189), .A2(new_n192), .A3(new_n193), .A4(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n191), .A2(G104), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n188), .A2(G107), .ZN(new_n197));
  OAI21_X1  g011(.A(G101), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n187), .B1(new_n195), .B2(new_n198), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n198), .A2(new_n187), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G128), .ZN(new_n208));
  OR2_X1    g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  OR2_X1    g023(.A1(new_n203), .A2(G128), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n202), .A2(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(new_n208), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n201), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT10), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT11), .ZN(new_n217));
  INV_X1    g031(.A(G134), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(G137), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(G137), .ZN(new_n220));
  INV_X1    g034(.A(G137), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(KEYINPUT11), .A3(G134), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G131), .ZN(new_n224));
  INV_X1    g038(.A(G131), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n219), .A2(new_n222), .A3(new_n225), .A4(new_n220), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n201), .A2(KEYINPUT10), .A3(new_n213), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n189), .A2(new_n192), .A3(new_n194), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G101), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(KEYINPUT4), .A3(new_n195), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n204), .A2(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  OAI22_X1  g050(.A1(new_n233), .A2(new_n211), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n203), .A2(new_n205), .A3(new_n234), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n230), .A2(new_n240), .A3(G101), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n232), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n216), .A2(new_n228), .A3(new_n229), .A4(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(G110), .B(G140), .ZN(new_n244));
  INV_X1    g058(.A(G227), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(G953), .ZN(new_n246));
  XOR2_X1   g060(.A(new_n244), .B(new_n246), .Z(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT79), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT78), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n195), .A2(new_n198), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT76), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n198), .A2(new_n187), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n213), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n228), .B1(new_n257), .B2(new_n214), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(KEYINPUT12), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT12), .ZN(new_n260));
  AOI211_X1 g074(.A(new_n260), .B(new_n228), .C1(new_n257), .C2(new_n214), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n251), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n255), .A2(new_n256), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n201), .A2(new_n213), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n227), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n260), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n258), .A2(KEYINPUT12), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(KEYINPUT78), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n243), .A2(KEYINPUT79), .A3(new_n247), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n250), .A2(new_n262), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n247), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n216), .A2(new_n242), .ZN(new_n272));
  INV_X1    g086(.A(new_n229), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n227), .A2(KEYINPUT77), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n275), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n272), .A2(new_n277), .A3(new_n273), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n271), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n270), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G469), .ZN(new_n281));
  INV_X1    g095(.A(G902), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n281), .A2(new_n282), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  OR3_X1    g099(.A1(new_n276), .A2(new_n278), .A3(new_n271), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n243), .B1(new_n259), .B2(new_n261), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n271), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n283), .B(new_n285), .C1(new_n281), .C2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT80), .ZN(new_n291));
  INV_X1    g105(.A(G221), .ZN(new_n292));
  XOR2_X1   g106(.A(KEYINPUT9), .B(G234), .Z(new_n293));
  AOI21_X1  g107(.A(new_n292), .B1(new_n293), .B2(new_n282), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n290), .A2(new_n291), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n291), .B1(new_n290), .B2(new_n295), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(KEYINPUT69), .A2(G237), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(KEYINPUT69), .A2(G237), .ZN(new_n301));
  AOI21_X1  g115(.A(G953), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(G143), .B1(new_n302), .B2(G214), .ZN(new_n303));
  INV_X1    g117(.A(G953), .ZN(new_n304));
  INV_X1    g118(.A(new_n301), .ZN(new_n305));
  OAI211_X1 g119(.A(G214), .B(new_n304), .C1(new_n305), .C2(new_n299), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(new_n204), .ZN(new_n307));
  OAI21_X1  g121(.A(G131), .B1(new_n303), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n302), .A2(G143), .A3(G214), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n306), .A2(new_n204), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n225), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT16), .ZN(new_n313));
  INV_X1    g127(.A(G140), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(G125), .ZN(new_n315));
  INV_X1    g129(.A(G125), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n314), .ZN(new_n317));
  NAND2_X1  g131(.A1(G125), .A2(G140), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n315), .B1(new_n320), .B2(new_n313), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(new_n202), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n320), .A2(KEYINPUT19), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT84), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n317), .A2(KEYINPUT84), .A3(new_n318), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n323), .B1(new_n327), .B2(KEYINPUT19), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n322), .B1(new_n328), .B2(new_n202), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n303), .A2(new_n307), .ZN(new_n330));
  NAND2_X1  g144(.A1(KEYINPUT18), .A2(G131), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(G146), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n319), .A2(new_n202), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n330), .A2(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n225), .B1(new_n309), .B2(new_n310), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT18), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n312), .A2(new_n329), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(G113), .B(G122), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(new_n188), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT85), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n329), .A2(new_n312), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n334), .A2(new_n336), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT85), .ZN(new_n344));
  INV_X1    g158(.A(new_n339), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n321), .B(G146), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n335), .A2(KEYINPUT17), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n347), .B(new_n348), .C1(new_n312), .C2(KEYINPUT17), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n339), .A3(new_n342), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n340), .A2(new_n346), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G475), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(new_n282), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT20), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT20), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n351), .A2(new_n355), .A3(new_n352), .A4(new_n282), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n350), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n339), .B1(new_n349), .B2(new_n342), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n282), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT86), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n361), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(G475), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n357), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(G128), .B(G143), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n366), .B(new_n218), .ZN(new_n367));
  INV_X1    g181(.A(G122), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G116), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n368), .A2(G116), .ZN(new_n371));
  OR3_X1    g185(.A1(new_n370), .A2(G107), .A3(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(KEYINPUT88), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT14), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n369), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT89), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n375), .B(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n377), .B1(new_n374), .B2(new_n371), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n367), .B(new_n373), .C1(new_n378), .C2(new_n191), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n218), .B1(new_n366), .B2(KEYINPUT13), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n204), .A2(G128), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n380), .B1(KEYINPUT13), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(KEYINPUT87), .ZN(new_n383));
  OAI21_X1  g197(.A(G107), .B1(new_n370), .B2(new_n371), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n372), .A2(new_n384), .B1(new_n218), .B2(new_n366), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n379), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT75), .B(G217), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n293), .A2(new_n304), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT90), .ZN(new_n391));
  INV_X1    g205(.A(new_n389), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n379), .A2(new_n392), .A3(new_n386), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n387), .A2(KEYINPUT90), .A3(new_n389), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n282), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G478), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n397), .A2(KEYINPUT15), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n396), .B(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G952), .ZN(new_n400));
  AOI211_X1 g214(.A(G953), .B(new_n400), .C1(G234), .C2(G237), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT21), .B(G898), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n402), .B(KEYINPUT91), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AOI211_X1 g218(.A(new_n282), .B(new_n304), .C1(G234), .C2(G237), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n401), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n365), .A2(new_n399), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G119), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G116), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT66), .ZN(new_n411));
  INV_X1    g225(.A(G116), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n411), .B1(new_n412), .B2(G119), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n409), .A2(KEYINPUT66), .A3(G116), .ZN(new_n414));
  OAI211_X1 g228(.A(KEYINPUT5), .B(new_n410), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n410), .A2(KEYINPUT5), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(G113), .A3(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT2), .B(G113), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n419), .B(new_n410), .C1(new_n414), .C2(new_n413), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n253), .A2(new_n417), .A3(new_n420), .A4(new_n254), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT81), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT81), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n201), .A2(new_n423), .A3(new_n420), .A4(new_n417), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n410), .B1(new_n413), .B2(new_n414), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n418), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n241), .A3(new_n232), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n422), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  XOR2_X1   g243(.A(G110), .B(G122), .Z(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT82), .ZN(new_n432));
  INV_X1    g246(.A(new_n430), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n422), .A2(new_n424), .A3(new_n433), .A4(new_n428), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT6), .A4(new_n434), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n431), .A2(KEYINPUT6), .A3(new_n434), .ZN(new_n436));
  OAI21_X1  g250(.A(KEYINPUT82), .B1(new_n431), .B2(KEYINPUT6), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n239), .A2(G125), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n439), .B1(new_n256), .B2(G125), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n304), .A2(G224), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n440), .B(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT83), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n441), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n442), .B1(KEYINPUT7), .B2(new_n446), .ZN(new_n447));
  XOR2_X1   g261(.A(new_n430), .B(KEYINPUT8), .Z(new_n448));
  AOI21_X1  g262(.A(new_n201), .B1(new_n420), .B2(new_n417), .ZN(new_n449));
  INV_X1    g263(.A(new_n421), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OR3_X1    g265(.A1(new_n440), .A2(KEYINPUT7), .A3(new_n446), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n447), .A2(new_n451), .A3(new_n434), .A4(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n453), .A2(new_n282), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n438), .A2(KEYINPUT83), .A3(new_n442), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n445), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G210), .B1(G237), .B2(G902), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n445), .A2(new_n457), .A3(new_n454), .A4(new_n455), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G214), .B1(G237), .B2(G902), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n298), .A2(new_n408), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT32), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT31), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT65), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n221), .A2(G134), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n220), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n467), .B1(new_n469), .B2(G131), .ZN(new_n470));
  AOI211_X1 g284(.A(KEYINPUT65), .B(new_n225), .C1(new_n220), .C2(new_n468), .ZN(new_n471));
  OAI211_X1 g285(.A(KEYINPUT68), .B(new_n226), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(G134), .B(G137), .ZN(new_n474));
  OAI21_X1  g288(.A(KEYINPUT65), .B1(new_n474), .B2(new_n225), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n469), .A2(new_n467), .A3(G131), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT68), .B1(new_n477), .B2(new_n226), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n213), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT67), .ZN(new_n480));
  AOI221_X4 g294(.A(new_n480), .B1(new_n237), .B2(new_n238), .C1(new_n224), .C2(new_n226), .ZN(new_n481));
  AOI21_X1  g295(.A(KEYINPUT67), .B1(new_n227), .B2(new_n239), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n479), .A2(new_n483), .A3(KEYINPUT30), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n227), .A2(new_n239), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT64), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n213), .A2(new_n226), .A3(new_n477), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT64), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n227), .A2(new_n488), .A3(new_n239), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT30), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n484), .A2(new_n492), .A3(new_n427), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(G101), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n302), .A2(G210), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n495), .B(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n427), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n479), .A2(new_n483), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n493), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT70), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT70), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n493), .A2(new_n502), .A3(new_n497), .A4(new_n499), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n466), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n479), .A2(new_n485), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT71), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n479), .A2(KEYINPUT71), .A3(new_n485), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n498), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT28), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n490), .A2(new_n427), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n499), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT28), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n497), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n500), .A2(KEYINPUT31), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n504), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(G472), .A2(G902), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n465), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n501), .A2(new_n503), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT31), .ZN(new_n522));
  INV_X1    g336(.A(new_n515), .ZN(new_n523));
  INV_X1    g337(.A(new_n516), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(KEYINPUT32), .A3(new_n518), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT72), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n520), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n518), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(KEYINPUT72), .A3(new_n465), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n479), .A2(new_n483), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n427), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT74), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XOR2_X1   g348(.A(new_n499), .B(KEYINPUT73), .Z(new_n535));
  AOI21_X1  g349(.A(new_n510), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n511), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(KEYINPUT29), .A3(new_n497), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n493), .A2(new_n499), .ZN(new_n540));
  INV_X1    g354(.A(new_n497), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n543), .A2(KEYINPUT29), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n511), .A2(new_n497), .A3(new_n514), .ZN(new_n545));
  AOI21_X1  g359(.A(G902), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n539), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n528), .A2(new_n530), .B1(G472), .B2(new_n547), .ZN(new_n548));
  OR3_X1    g362(.A1(new_n409), .A2(KEYINPUT23), .A3(G128), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT23), .B1(new_n409), .B2(G128), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n549), .A2(new_n550), .B1(new_n409), .B2(G128), .ZN(new_n551));
  INV_X1    g365(.A(G110), .ZN(new_n552));
  XOR2_X1   g366(.A(G119), .B(G128), .Z(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT24), .B(G110), .ZN(new_n554));
  OAI22_X1  g368(.A1(new_n551), .A2(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n551), .A2(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n333), .B1(new_n321), .B2(new_n202), .ZN(new_n557));
  OAI22_X1  g371(.A1(new_n347), .A2(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n304), .A2(G221), .A3(G234), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT22), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(G137), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n558), .B(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  OR3_X1    g377(.A1(new_n563), .A2(KEYINPUT25), .A3(G902), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n282), .A2(G234), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT25), .B1(new_n563), .B2(G902), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n564), .A2(new_n565), .A3(new_n388), .A4(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(G902), .B1(new_n388), .B2(new_n565), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n548), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n464), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(G101), .ZN(G3));
  OAI21_X1  g388(.A(G472), .B1(new_n517), .B2(G902), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n529), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n298), .A2(new_n571), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT92), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT93), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n461), .B2(new_n462), .ZN(new_n580));
  INV_X1    g394(.A(new_n462), .ZN(new_n581));
  AOI211_X1 g395(.A(KEYINPUT93), .B(new_n581), .C1(new_n459), .C2(new_n460), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n396), .A2(new_n397), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n390), .A2(KEYINPUT33), .A3(new_n393), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n394), .A2(new_n395), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n584), .B1(new_n585), .B2(KEYINPUT33), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n282), .A2(G478), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n583), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n365), .A2(new_n588), .ZN(new_n589));
  NOR4_X1   g403(.A1(new_n580), .A2(new_n582), .A3(new_n406), .A4(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n578), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT34), .B(G104), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(G6));
  NOR2_X1   g408(.A1(new_n580), .A2(new_n582), .ZN(new_n595));
  INV_X1    g409(.A(new_n406), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n354), .A2(KEYINPUT94), .A3(new_n356), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT94), .B1(new_n354), .B2(new_n356), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n364), .B(new_n399), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n595), .A2(new_n596), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n578), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT35), .B(G107), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G9));
  INV_X1    g419(.A(new_n576), .ZN(new_n606));
  INV_X1    g420(.A(new_n561), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n607), .A2(KEYINPUT36), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n558), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n568), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n567), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n464), .A2(new_n606), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT37), .B(G110), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G12));
  INV_X1    g430(.A(KEYINPUT97), .ZN(new_n617));
  INV_X1    g431(.A(G900), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n405), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n401), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n617), .B1(new_n600), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n398), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n396), .B(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT94), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n357), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n625), .B1(new_n627), .B2(new_n597), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n628), .A2(KEYINPUT97), .A3(new_n364), .A4(new_n621), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n611), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n528), .A2(new_n530), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n547), .A2(G472), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n298), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n595), .A2(new_n630), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT98), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n548), .A2(new_n298), .A3(new_n631), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT98), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n638), .A2(new_n639), .A3(new_n595), .A4(new_n630), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G128), .ZN(G30));
  XOR2_X1   g456(.A(new_n621), .B(KEYINPUT39), .Z(new_n643));
  OR2_X1    g457(.A1(new_n298), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT100), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT40), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n581), .ZN(new_n648));
  INV_X1    g462(.A(new_n365), .ZN(new_n649));
  AOI211_X1 g463(.A(new_n649), .B(new_n625), .C1(new_n645), .C2(new_n646), .ZN(new_n650));
  INV_X1    g464(.A(new_n521), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n497), .B1(new_n534), .B2(new_n535), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n282), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(G472), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n632), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(new_n611), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n461), .B(KEYINPUT99), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT38), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n648), .A2(new_n650), .A3(new_n657), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G143), .ZN(G45));
  NOR2_X1   g476(.A1(new_n589), .A2(new_n622), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n595), .A2(new_n634), .A3(new_n635), .A4(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n638), .A2(KEYINPUT101), .A3(new_n595), .A4(new_n663), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G146), .ZN(G48));
  INV_X1    g483(.A(new_n283), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n281), .B1(new_n280), .B2(new_n282), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n295), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n548), .A2(new_n673), .A3(new_n571), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n590), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT41), .B(G113), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G15));
  NAND4_X1  g491(.A1(new_n674), .A2(new_n596), .A3(new_n595), .A4(new_n601), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G116), .ZN(G18));
  INV_X1    g493(.A(new_n673), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT102), .B1(new_n595), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n682));
  NOR4_X1   g496(.A1(new_n580), .A2(new_n582), .A3(new_n682), .A4(new_n673), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n407), .B(new_n634), .C1(new_n681), .C2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G119), .ZN(G21));
  NOR2_X1   g499(.A1(new_n504), .A2(new_n516), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(new_n538), .B2(new_n497), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n518), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n575), .ZN(new_n689));
  OAI21_X1  g503(.A(KEYINPUT103), .B1(new_n689), .B2(new_n571), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n688), .A2(new_n575), .A3(new_n691), .A4(new_n570), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n649), .A2(new_n625), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n673), .A2(new_n406), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n693), .A2(new_n595), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G122), .ZN(G24));
  INV_X1    g511(.A(new_n663), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n698), .A2(new_n631), .A3(new_n689), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n699), .B1(new_n681), .B2(new_n683), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G125), .ZN(G27));
  NAND3_X1  g515(.A1(new_n633), .A2(new_n520), .A3(new_n526), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n702), .A2(new_n570), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n288), .B(KEYINPUT104), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n704), .A2(new_n286), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G469), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n283), .A2(new_n285), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n294), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n461), .A2(new_n581), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n703), .A2(new_n663), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n708), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n711), .A2(new_n548), .A3(new_n571), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n698), .A2(KEYINPUT42), .ZN(new_n713));
  AOI22_X1  g527(.A1(new_n710), .A2(KEYINPUT42), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G131), .ZN(G33));
  NAND2_X1  g529(.A1(new_n712), .A2(new_n630), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT105), .B(G134), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G36));
  AND2_X1   g532(.A1(new_n705), .A2(KEYINPUT45), .ZN(new_n719));
  OR2_X1    g533(.A1(new_n719), .A2(KEYINPUT106), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n281), .B1(new_n289), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n719), .A2(KEYINPUT106), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n720), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n285), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT46), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n724), .A2(KEYINPUT46), .A3(new_n285), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n283), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n295), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n643), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n649), .A2(new_n588), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT43), .ZN(new_n733));
  OR3_X1    g547(.A1(new_n733), .A2(new_n606), .A3(new_n631), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT107), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n734), .A2(new_n735), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n731), .A2(new_n737), .A3(new_n709), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G137), .ZN(G39));
  INV_X1    g554(.A(KEYINPUT47), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n730), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n729), .A2(KEYINPUT47), .A3(new_n295), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n698), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(new_n548), .A3(new_n571), .A4(new_n709), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G140), .ZN(G42));
  AND2_X1   g560(.A1(new_n595), .A2(new_n694), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n708), .A2(new_n631), .A3(new_n621), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT110), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n748), .A2(KEYINPUT110), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n747), .A2(new_n655), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n641), .A2(new_n668), .A3(new_n700), .A4(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n640), .A2(new_n637), .B1(new_n666), .B2(new_n667), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n755), .A2(KEYINPUT52), .A3(new_n700), .A4(new_n751), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n627), .A2(new_n597), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n758), .A2(new_n364), .A3(new_n625), .A4(new_n621), .ZN(new_n759));
  NOR4_X1   g573(.A1(new_n548), .A2(new_n298), .A3(new_n631), .A4(new_n759), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n699), .A2(new_n708), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n709), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n714), .A2(new_n762), .A3(new_n716), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n463), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n589), .B1(new_n365), .B2(new_n625), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n577), .A2(new_n596), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n573), .A3(new_n612), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n769));
  INV_X1    g583(.A(new_n634), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n463), .A2(KEYINPUT93), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n461), .A2(new_n579), .A3(new_n462), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n680), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n682), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n595), .A2(KEYINPUT102), .A3(new_n680), .ZN(new_n775));
  AOI211_X1 g589(.A(new_n408), .B(new_n770), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n675), .A2(new_n678), .A3(new_n696), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n769), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n693), .A2(new_n595), .A3(new_n694), .ZN(new_n779));
  AOI22_X1  g593(.A1(new_n779), .A2(new_n695), .B1(new_n590), .B2(new_n674), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n780), .A2(new_n684), .A3(KEYINPUT109), .A4(new_n678), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n768), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n757), .A2(KEYINPUT53), .A3(new_n764), .A4(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n786));
  INV_X1    g600(.A(new_n757), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n778), .A2(new_n781), .ZN(new_n788));
  INV_X1    g602(.A(new_n768), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n764), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n786), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  AOI211_X1 g605(.A(new_n768), .B(new_n763), .C1(new_n778), .C2(new_n781), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n792), .A2(KEYINPUT111), .A3(KEYINPUT53), .A4(new_n757), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n785), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT54), .ZN(new_n795));
  AOI211_X1 g609(.A(new_n776), .B(new_n777), .C1(new_n754), .C2(new_n756), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(KEYINPUT53), .A3(new_n764), .A4(new_n789), .ZN(new_n797));
  XOR2_X1   g611(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n797), .A2(new_n791), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n795), .A2(KEYINPUT113), .A3(new_n800), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n709), .A2(new_n680), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT116), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n806), .A2(new_n570), .A3(new_n401), .A4(new_n656), .ZN(new_n807));
  OAI211_X1 g621(.A(G952), .B(new_n304), .C1(new_n807), .C2(new_n589), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n774), .A2(new_n775), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n733), .A2(new_n620), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n810), .A2(new_n693), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n808), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT118), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n806), .A2(new_n810), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n703), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT48), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n807), .A2(new_n365), .A3(new_n588), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n818), .B(KEYINPUT117), .Z(new_n819));
  AND4_X1   g633(.A1(new_n581), .A2(new_n659), .A3(new_n680), .A4(new_n811), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n821), .A2(KEYINPUT115), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n823), .B1(KEYINPUT115), .B2(new_n821), .ZN(new_n824));
  XOR2_X1   g638(.A(new_n672), .B(KEYINPUT114), .Z(new_n825));
  OAI211_X1 g639(.A(new_n742), .B(new_n743), .C1(new_n295), .C2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n709), .A3(new_n811), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n820), .A2(new_n822), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n819), .A2(new_n824), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n814), .A2(new_n575), .A3(new_n611), .A4(new_n688), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  OR3_X1    g645(.A1(new_n829), .A2(KEYINPUT51), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT51), .B1(new_n829), .B2(new_n831), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n817), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n803), .A2(new_n804), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n400), .A2(new_n304), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n803), .A2(KEYINPUT119), .A3(new_n804), .A4(new_n834), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n672), .B(KEYINPUT49), .ZN(new_n841));
  NOR4_X1   g655(.A1(new_n732), .A2(new_n571), .A3(new_n294), .A4(new_n581), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT108), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n659), .A2(new_n656), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n840), .A2(new_n844), .ZN(G75));
  INV_X1    g659(.A(KEYINPUT56), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n797), .A2(new_n791), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(G902), .ZN(new_n848));
  INV_X1    g662(.A(G210), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n438), .B(new_n442), .ZN(new_n851));
  XOR2_X1   g665(.A(new_n851), .B(KEYINPUT55), .Z(new_n852));
  OAI21_X1  g666(.A(new_n852), .B1(KEYINPUT120), .B2(KEYINPUT56), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n304), .A2(G952), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n853), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n846), .B(new_n857), .C1(new_n848), .C2(new_n849), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n854), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT121), .ZN(G51));
  NAND2_X1  g674(.A1(new_n847), .A2(new_n798), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n800), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n862), .B1(new_n863), .B2(new_n284), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n285), .A2(KEYINPUT57), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n280), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n848), .A2(new_n724), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n855), .B1(new_n866), .B2(new_n867), .ZN(G54));
  NAND4_X1  g682(.A1(new_n847), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n869));
  INV_X1    g683(.A(new_n351), .ZN(new_n870));
  OR3_X1    g684(.A1(new_n869), .A2(KEYINPUT122), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n855), .B1(new_n869), .B2(new_n870), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT122), .B1(new_n869), .B2(new_n870), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT123), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n871), .A2(new_n876), .A3(new_n872), .A4(new_n873), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n875), .A2(new_n877), .ZN(G60));
  NAND2_X1  g692(.A1(G478), .A2(G902), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT59), .Z(new_n880));
  AOI211_X1 g694(.A(new_n586), .B(new_n880), .C1(new_n861), .C2(new_n800), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n803), .A2(new_n804), .ZN(new_n882));
  INV_X1    g696(.A(new_n880), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI211_X1 g698(.A(new_n855), .B(new_n881), .C1(new_n884), .C2(new_n586), .ZN(G63));
  NAND2_X1  g699(.A1(G217), .A2(G902), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT60), .Z(new_n887));
  NAND2_X1  g701(.A1(new_n847), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n847), .A2(KEYINPUT124), .A3(new_n887), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n609), .B(KEYINPUT125), .Z(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n890), .A2(new_n563), .A3(new_n891), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n856), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n894), .A2(KEYINPUT61), .A3(new_n856), .A4(new_n895), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(G66));
  INV_X1    g714(.A(G224), .ZN(new_n901));
  OAI21_X1  g715(.A(G953), .B1(new_n404), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n902), .B1(new_n782), .B2(G953), .ZN(new_n903));
  INV_X1    g717(.A(new_n438), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(G898), .B2(new_n304), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n903), .B(new_n905), .ZN(G69));
  NAND2_X1  g720(.A1(new_n484), .A2(new_n492), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(new_n328), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n304), .B1(new_n245), .B2(G900), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n731), .A2(new_n747), .A3(new_n703), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n745), .A2(new_n714), .A3(new_n716), .A4(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n755), .A2(new_n700), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n739), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  AOI211_X1 g728(.A(new_n908), .B(new_n909), .C1(new_n914), .C2(new_n304), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n909), .A2(G900), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n661), .A2(new_n912), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n745), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n645), .A2(new_n572), .A3(new_n709), .A4(new_n766), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT126), .Z(new_n922));
  NAND3_X1  g736(.A1(new_n922), .A2(new_n304), .A3(new_n739), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n916), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n915), .B1(new_n924), .B2(new_n908), .ZN(G72));
  NAND2_X1  g739(.A1(new_n914), .A2(new_n782), .ZN(new_n926));
  NAND2_X1  g740(.A1(G472), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT63), .Z(new_n928));
  AOI211_X1 g742(.A(new_n497), .B(new_n540), .C1(new_n926), .C2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n922), .A2(new_n739), .A3(new_n782), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n920), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n931), .A2(new_n497), .A3(new_n540), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n856), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n794), .B(new_n928), .C1(new_n543), .C2(new_n651), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT127), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  AOI211_X1 g751(.A(new_n929), .B(new_n933), .C1(new_n936), .C2(new_n937), .ZN(G57));
endmodule


