

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X2 U550 ( .A(n662), .Z(n679) );
  AND2_X2 U551 ( .A1(n677), .A2(n519), .ZN(n688) );
  NOR2_X2 U552 ( .A1(n694), .A2(KEYINPUT33), .ZN(n695) );
  BUF_X1 U553 ( .A(n707), .Z(n708) );
  XNOR2_X2 U554 ( .A(n689), .B(KEYINPUT101), .ZN(n703) );
  NOR2_X2 U555 ( .A1(n688), .A2(n687), .ZN(n689) );
  INV_X1 U556 ( .A(G2105), .ZN(n530) );
  NAND2_X1 U557 ( .A1(G8), .A2(n662), .ZN(n753) );
  INV_X1 U558 ( .A(KEYINPUT87), .ZN(n526) );
  NOR2_X1 U559 ( .A1(n627), .A2(G1384), .ZN(n748) );
  XNOR2_X1 U560 ( .A(n700), .B(n699), .ZN(n702) );
  INV_X1 U561 ( .A(KEYINPUT104), .ZN(n699) );
  INV_X1 U562 ( .A(n933), .ZN(n701) );
  XNOR2_X1 U563 ( .A(n525), .B(n524), .ZN(n707) );
  NOR2_X1 U564 ( .A1(G2105), .A2(G2104), .ZN(n525) );
  XNOR2_X1 U565 ( .A(n538), .B(n537), .ZN(n540) );
  INV_X1 U566 ( .A(KEYINPUT23), .ZN(n537) );
  BUF_X1 U567 ( .A(n627), .Z(G164) );
  BUF_X1 U568 ( .A(n626), .Z(G160) );
  XNOR2_X1 U569 ( .A(KEYINPUT105), .B(KEYINPUT40), .ZN(n518) );
  XOR2_X1 U570 ( .A(KEYINPUT95), .B(n676), .Z(n519) );
  OR2_X1 U571 ( .A1(n754), .A2(n753), .ZN(n520) );
  AND2_X1 U572 ( .A1(n755), .A2(n520), .ZN(n521) );
  OR2_X1 U573 ( .A1(n753), .A2(n697), .ZN(n522) );
  INV_X1 U574 ( .A(KEYINPUT28), .ZN(n650) );
  INV_X1 U575 ( .A(KEYINPUT29), .ZN(n654) );
  NOR2_X1 U576 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U577 ( .A1(G1966), .A2(n753), .ZN(n672) );
  INV_X1 U578 ( .A(KEYINPUT17), .ZN(n524) );
  NAND2_X1 U579 ( .A1(n813), .A2(G56), .ZN(n621) );
  INV_X1 U580 ( .A(KEYINPUT1), .ZN(n547) );
  INV_X1 U581 ( .A(KEYINPUT66), .ZN(n531) );
  NOR2_X1 U582 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U583 ( .A1(n994), .A2(G114), .ZN(n533) );
  XOR2_X1 U584 ( .A(G543), .B(KEYINPUT0), .Z(n588) );
  INV_X1 U585 ( .A(KEYINPUT7), .ZN(n575) );
  XNOR2_X1 U586 ( .A(n576), .B(n575), .ZN(n577) );
  NOR2_X1 U587 ( .A1(n536), .A2(n535), .ZN(n627) );
  NOR2_X1 U588 ( .A1(n565), .A2(n564), .ZN(G171) );
  NOR2_X2 U589 ( .A1(n530), .A2(G2104), .ZN(n993) );
  NAND2_X1 U590 ( .A1(G126), .A2(n993), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n523), .B(KEYINPUT86), .ZN(n529) );
  NAND2_X1 U592 ( .A1(G138), .A2(n707), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(n528) );
  NAND2_X1 U594 ( .A1(n529), .A2(n528), .ZN(n536) );
  AND2_X4 U595 ( .A1(n530), .A2(G2104), .ZN(n997) );
  NAND2_X1 U596 ( .A1(G102), .A2(n997), .ZN(n534) );
  NAND2_X1 U597 ( .A1(G2104), .A2(G2105), .ZN(n532) );
  XNOR2_X2 U598 ( .A(n532), .B(n531), .ZN(n994) );
  NAND2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n535) );
  INV_X1 U600 ( .A(KEYINPUT65), .ZN(n542) );
  NAND2_X1 U601 ( .A1(n997), .A2(G101), .ZN(n538) );
  NAND2_X1 U602 ( .A1(n993), .A2(G125), .ZN(n539) );
  NAND2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U604 ( .A(n542), .B(n541), .ZN(n546) );
  NAND2_X1 U605 ( .A1(G137), .A2(n707), .ZN(n544) );
  NAND2_X1 U606 ( .A1(G113), .A2(n994), .ZN(n543) );
  NAND2_X1 U607 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X2 U608 ( .A1(n546), .A2(n545), .ZN(n626) );
  INV_X1 U609 ( .A(G651), .ZN(n553) );
  NOR2_X1 U610 ( .A1(G543), .A2(n553), .ZN(n548) );
  XNOR2_X2 U611 ( .A(n548), .B(n547), .ZN(n813) );
  NAND2_X1 U612 ( .A1(n813), .A2(G65), .ZN(n551) );
  NOR2_X1 U613 ( .A1(G651), .A2(n588), .ZN(n549) );
  XNOR2_X2 U614 ( .A(KEYINPUT64), .B(n549), .ZN(n809) );
  NAND2_X1 U615 ( .A1(G53), .A2(n809), .ZN(n550) );
  NAND2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(KEYINPUT69), .B(n552), .ZN(n557) );
  NOR2_X2 U618 ( .A1(G543), .A2(G651), .ZN(n805) );
  NAND2_X1 U619 ( .A1(G91), .A2(n805), .ZN(n555) );
  NOR2_X2 U620 ( .A1(n588), .A2(n553), .ZN(n806) );
  NAND2_X1 U621 ( .A1(G78), .A2(n806), .ZN(n554) );
  AND2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(G299) );
  NAND2_X1 U624 ( .A1(G90), .A2(n805), .ZN(n559) );
  NAND2_X1 U625 ( .A1(G77), .A2(n806), .ZN(n558) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(KEYINPUT9), .ZN(n562) );
  NAND2_X1 U628 ( .A1(G52), .A2(n809), .ZN(n561) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n813), .A2(G64), .ZN(n563) );
  XOR2_X1 U631 ( .A(KEYINPUT68), .B(n563), .Z(n564) );
  NAND2_X1 U632 ( .A1(G51), .A2(n809), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n813), .A2(G63), .ZN(n566) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(KEYINPUT6), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n805), .A2(G89), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n569), .B(KEYINPUT4), .ZN(n571) );
  NAND2_X1 U638 ( .A1(G76), .A2(n806), .ZN(n570) );
  NAND2_X1 U639 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U640 ( .A(n572), .B(KEYINPUT5), .Z(n573) );
  NOR2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n576) );
  XNOR2_X1 U642 ( .A(KEYINPUT74), .B(n577), .ZN(G168) );
  XOR2_X1 U643 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U644 ( .A1(G88), .A2(n805), .ZN(n579) );
  NAND2_X1 U645 ( .A1(G75), .A2(n806), .ZN(n578) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U647 ( .A1(n813), .A2(G62), .ZN(n581) );
  NAND2_X1 U648 ( .A1(G50), .A2(n809), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U650 ( .A1(n583), .A2(n582), .ZN(G166) );
  INV_X1 U651 ( .A(G166), .ZN(G303) );
  NAND2_X1 U652 ( .A1(G651), .A2(G74), .ZN(n585) );
  NAND2_X1 U653 ( .A1(G49), .A2(n809), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U655 ( .A1(n813), .A2(n586), .ZN(n587) );
  XOR2_X1 U656 ( .A(KEYINPUT81), .B(n587), .Z(n590) );
  NAND2_X1 U657 ( .A1(n588), .A2(G87), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n590), .A2(n589), .ZN(G288) );
  NAND2_X1 U659 ( .A1(G73), .A2(n806), .ZN(n591) );
  XNOR2_X1 U660 ( .A(n591), .B(KEYINPUT2), .ZN(n598) );
  NAND2_X1 U661 ( .A1(n813), .A2(G61), .ZN(n593) );
  NAND2_X1 U662 ( .A1(G48), .A2(n809), .ZN(n592) );
  NAND2_X1 U663 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U664 ( .A1(n805), .A2(G86), .ZN(n594) );
  XOR2_X1 U665 ( .A(KEYINPUT82), .B(n594), .Z(n595) );
  NOR2_X1 U666 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U667 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U668 ( .A(KEYINPUT83), .B(n599), .Z(G305) );
  NAND2_X1 U669 ( .A1(n813), .A2(G60), .ZN(n601) );
  NAND2_X1 U670 ( .A1(G47), .A2(n809), .ZN(n600) );
  NAND2_X1 U671 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U672 ( .A1(G85), .A2(n805), .ZN(n603) );
  NAND2_X1 U673 ( .A1(G72), .A2(n806), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U675 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U676 ( .A(n606), .B(KEYINPUT67), .ZN(G290) );
  NAND2_X1 U677 ( .A1(G66), .A2(n813), .ZN(n613) );
  NAND2_X1 U678 ( .A1(G92), .A2(n805), .ZN(n608) );
  NAND2_X1 U679 ( .A1(G54), .A2(n809), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U681 ( .A1(G79), .A2(n806), .ZN(n609) );
  XNOR2_X1 U682 ( .A(KEYINPUT73), .B(n609), .ZN(n610) );
  NOR2_X1 U683 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U684 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X2 U685 ( .A(n614), .B(KEYINPUT15), .ZN(n1018) );
  INV_X1 U686 ( .A(n1018), .ZN(n625) );
  NAND2_X1 U687 ( .A1(n805), .A2(G81), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n615), .B(KEYINPUT12), .ZN(n617) );
  NAND2_X1 U689 ( .A1(G68), .A2(n806), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U691 ( .A(n618), .B(KEYINPUT13), .ZN(n620) );
  NAND2_X1 U692 ( .A1(G43), .A2(n809), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n623) );
  XOR2_X1 U694 ( .A(KEYINPUT14), .B(n621), .Z(n622) );
  XOR2_X1 U695 ( .A(KEYINPUT70), .B(n624), .Z(n778) );
  NOR2_X1 U696 ( .A1(n625), .A2(n778), .ZN(n633) );
  NAND2_X1 U697 ( .A1(n626), .A2(G40), .ZN(n747) );
  INV_X1 U698 ( .A(n747), .ZN(n628) );
  NAND2_X2 U699 ( .A1(n628), .A2(n748), .ZN(n662) );
  INV_X2 U700 ( .A(n662), .ZN(n656) );
  NAND2_X1 U701 ( .A1(n656), .A2(G1996), .ZN(n629) );
  XNOR2_X1 U702 ( .A(n629), .B(KEYINPUT26), .ZN(n631) );
  NAND2_X1 U703 ( .A1(n679), .A2(G1341), .ZN(n630) );
  NAND2_X1 U704 ( .A1(n631), .A2(n630), .ZN(n639) );
  INV_X1 U705 ( .A(n639), .ZN(n632) );
  NAND2_X1 U706 ( .A1(n633), .A2(n632), .ZN(n638) );
  AND2_X1 U707 ( .A1(n656), .A2(G2067), .ZN(n634) );
  XOR2_X1 U708 ( .A(n634), .B(KEYINPUT98), .Z(n636) );
  NAND2_X1 U709 ( .A1(n679), .A2(G1348), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U711 ( .A1(n638), .A2(n637), .ZN(n642) );
  NOR2_X1 U712 ( .A1(n639), .A2(n778), .ZN(n640) );
  OR2_X2 U713 ( .A1(n640), .A2(n1018), .ZN(n641) );
  NAND2_X1 U714 ( .A1(n642), .A2(n641), .ZN(n648) );
  INV_X1 U715 ( .A(G299), .ZN(n819) );
  NAND2_X1 U716 ( .A1(n656), .A2(G2072), .ZN(n643) );
  XNOR2_X1 U717 ( .A(n643), .B(KEYINPUT27), .ZN(n646) );
  NAND2_X1 U718 ( .A1(G1956), .A2(n662), .ZN(n644) );
  XNOR2_X1 U719 ( .A(n644), .B(KEYINPUT97), .ZN(n645) );
  NOR2_X1 U720 ( .A1(n646), .A2(n645), .ZN(n649) );
  NAND2_X1 U721 ( .A1(n819), .A2(n649), .ZN(n647) );
  NAND2_X1 U722 ( .A1(n648), .A2(n647), .ZN(n653) );
  NOR2_X1 U723 ( .A1(n649), .A2(n819), .ZN(n651) );
  XNOR2_X1 U724 ( .A(n651), .B(n650), .ZN(n652) );
  NAND2_X1 U725 ( .A1(n653), .A2(n652), .ZN(n655) );
  XNOR2_X1 U726 ( .A(n655), .B(n654), .ZN(n661) );
  XOR2_X1 U727 ( .A(G2078), .B(KEYINPUT25), .Z(n857) );
  NAND2_X1 U728 ( .A1(n656), .A2(n857), .ZN(n658) );
  NAND2_X1 U729 ( .A1(G1961), .A2(n679), .ZN(n657) );
  NAND2_X1 U730 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U731 ( .A(KEYINPUT96), .B(n659), .Z(n666) );
  NAND2_X1 U732 ( .A1(n666), .A2(G171), .ZN(n660) );
  NAND2_X1 U733 ( .A1(n661), .A2(n660), .ZN(n671) );
  NOR2_X1 U734 ( .A1(G2084), .A2(n679), .ZN(n675) );
  NOR2_X1 U735 ( .A1(n675), .A2(n672), .ZN(n663) );
  NAND2_X1 U736 ( .A1(G8), .A2(n663), .ZN(n664) );
  XNOR2_X1 U737 ( .A(n664), .B(KEYINPUT30), .ZN(n665) );
  NOR2_X1 U738 ( .A1(n665), .A2(G168), .ZN(n668) );
  NOR2_X1 U739 ( .A1(G171), .A2(n666), .ZN(n667) );
  XOR2_X1 U740 ( .A(KEYINPUT31), .B(n669), .Z(n670) );
  NAND2_X1 U741 ( .A1(n671), .A2(n670), .ZN(n678) );
  XNOR2_X1 U742 ( .A(n678), .B(KEYINPUT99), .ZN(n673) );
  NOR2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U744 ( .A(n674), .B(KEYINPUT100), .ZN(n677) );
  NAND2_X1 U745 ( .A1(G8), .A2(n675), .ZN(n676) );
  NAND2_X1 U746 ( .A1(G286), .A2(n678), .ZN(n684) );
  NOR2_X1 U747 ( .A1(G1971), .A2(n753), .ZN(n681) );
  NOR2_X1 U748 ( .A1(G2090), .A2(n679), .ZN(n680) );
  NOR2_X1 U749 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U750 ( .A1(n682), .A2(G303), .ZN(n683) );
  NAND2_X1 U751 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U752 ( .A1(n685), .A2(G8), .ZN(n686) );
  XOR2_X1 U753 ( .A(KEYINPUT32), .B(n686), .Z(n687) );
  NOR2_X1 U754 ( .A1(G1976), .A2(G288), .ZN(n696) );
  NOR2_X1 U755 ( .A1(G1971), .A2(G303), .ZN(n690) );
  NOR2_X1 U756 ( .A1(n696), .A2(n690), .ZN(n918) );
  NAND2_X1 U757 ( .A1(n703), .A2(n918), .ZN(n691) );
  NAND2_X1 U758 ( .A1(G1976), .A2(G288), .ZN(n917) );
  NAND2_X1 U759 ( .A1(n691), .A2(n917), .ZN(n692) );
  XNOR2_X1 U760 ( .A(n692), .B(KEYINPUT102), .ZN(n693) );
  NOR2_X1 U761 ( .A1(n693), .A2(n753), .ZN(n694) );
  XNOR2_X1 U762 ( .A(n695), .B(KEYINPUT103), .ZN(n698) );
  NAND2_X1 U763 ( .A1(n696), .A2(KEYINPUT33), .ZN(n697) );
  NAND2_X1 U764 ( .A1(n698), .A2(n522), .ZN(n700) );
  XNOR2_X1 U765 ( .A(G1981), .B(G305), .ZN(n933) );
  NAND2_X1 U766 ( .A1(n702), .A2(n701), .ZN(n756) );
  NOR2_X1 U767 ( .A1(G2090), .A2(G303), .ZN(n704) );
  NAND2_X1 U768 ( .A1(G8), .A2(n704), .ZN(n705) );
  NAND2_X1 U769 ( .A1(n703), .A2(n705), .ZN(n706) );
  NAND2_X1 U770 ( .A1(n753), .A2(n706), .ZN(n750) );
  NAND2_X1 U771 ( .A1(n994), .A2(G117), .ZN(n715) );
  NAND2_X1 U772 ( .A1(G129), .A2(n993), .ZN(n710) );
  NAND2_X1 U773 ( .A1(G141), .A2(n708), .ZN(n709) );
  NAND2_X1 U774 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U775 ( .A1(n997), .A2(G105), .ZN(n711) );
  XOR2_X1 U776 ( .A(KEYINPUT38), .B(n711), .Z(n712) );
  NOR2_X1 U777 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U778 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U779 ( .A(n716), .B(KEYINPUT92), .ZN(n992) );
  NOR2_X1 U780 ( .A1(G1996), .A2(n992), .ZN(n895) );
  NAND2_X1 U781 ( .A1(G1996), .A2(n992), .ZN(n717) );
  XOR2_X1 U782 ( .A(KEYINPUT93), .B(n717), .Z(n727) );
  NAND2_X1 U783 ( .A1(G119), .A2(n993), .ZN(n718) );
  XNOR2_X1 U784 ( .A(n718), .B(KEYINPUT90), .ZN(n725) );
  NAND2_X1 U785 ( .A1(G95), .A2(n997), .ZN(n720) );
  NAND2_X1 U786 ( .A1(G131), .A2(n708), .ZN(n719) );
  NAND2_X1 U787 ( .A1(n720), .A2(n719), .ZN(n723) );
  NAND2_X1 U788 ( .A1(G107), .A2(n994), .ZN(n721) );
  XNOR2_X1 U789 ( .A(KEYINPUT91), .B(n721), .ZN(n722) );
  NOR2_X1 U790 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U791 ( .A1(n725), .A2(n724), .ZN(n1006) );
  NAND2_X1 U792 ( .A1(G1991), .A2(n1006), .ZN(n726) );
  NAND2_X1 U793 ( .A1(n727), .A2(n726), .ZN(n758) );
  NOR2_X1 U794 ( .A1(G1986), .A2(G290), .ZN(n728) );
  NOR2_X1 U795 ( .A1(G1991), .A2(n1006), .ZN(n900) );
  NOR2_X1 U796 ( .A1(n728), .A2(n900), .ZN(n729) );
  NOR2_X1 U797 ( .A1(n758), .A2(n729), .ZN(n730) );
  NOR2_X1 U798 ( .A1(n895), .A2(n730), .ZN(n731) );
  XNOR2_X1 U799 ( .A(n731), .B(KEYINPUT39), .ZN(n744) );
  XNOR2_X1 U800 ( .A(G2067), .B(KEYINPUT37), .ZN(n732) );
  XNOR2_X1 U801 ( .A(n732), .B(KEYINPUT88), .ZN(n745) );
  NAND2_X1 U802 ( .A1(n997), .A2(G104), .ZN(n733) );
  XOR2_X1 U803 ( .A(KEYINPUT89), .B(n733), .Z(n735) );
  NAND2_X1 U804 ( .A1(n708), .A2(G140), .ZN(n734) );
  NAND2_X1 U805 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U806 ( .A(KEYINPUT34), .B(n736), .ZN(n741) );
  NAND2_X1 U807 ( .A1(G128), .A2(n993), .ZN(n738) );
  NAND2_X1 U808 ( .A1(G116), .A2(n994), .ZN(n737) );
  NAND2_X1 U809 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U810 ( .A(KEYINPUT35), .B(n739), .Z(n740) );
  NOR2_X1 U811 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U812 ( .A(KEYINPUT36), .B(n742), .ZN(n1015) );
  NOR2_X1 U813 ( .A1(n745), .A2(n1015), .ZN(n759) );
  INV_X1 U814 ( .A(n759), .ZN(n743) );
  NAND2_X1 U815 ( .A1(n744), .A2(n743), .ZN(n746) );
  NAND2_X1 U816 ( .A1(n745), .A2(n1015), .ZN(n901) );
  NAND2_X1 U817 ( .A1(n746), .A2(n901), .ZN(n749) );
  NOR2_X1 U818 ( .A1(n748), .A2(n747), .ZN(n760) );
  NAND2_X1 U819 ( .A1(n749), .A2(n760), .ZN(n757) );
  AND2_X1 U820 ( .A1(n750), .A2(n757), .ZN(n755) );
  NOR2_X1 U821 ( .A1(G1981), .A2(G305), .ZN(n751) );
  XOR2_X1 U822 ( .A(n751), .B(KEYINPUT94), .Z(n752) );
  XNOR2_X1 U823 ( .A(KEYINPUT24), .B(n752), .ZN(n754) );
  NAND2_X1 U824 ( .A1(n756), .A2(n521), .ZN(n765) );
  INV_X1 U825 ( .A(n757), .ZN(n763) );
  XOR2_X1 U826 ( .A(G1986), .B(G290), .Z(n914) );
  NOR2_X1 U827 ( .A1(n759), .A2(n758), .ZN(n892) );
  NAND2_X1 U828 ( .A1(n914), .A2(n892), .ZN(n761) );
  NAND2_X1 U829 ( .A1(n761), .A2(n760), .ZN(n762) );
  OR2_X1 U830 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U831 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U832 ( .A(n766), .B(n518), .ZN(G329) );
  XOR2_X1 U833 ( .A(G2443), .B(G2454), .Z(n768) );
  XNOR2_X1 U834 ( .A(G1341), .B(G1348), .ZN(n767) );
  XNOR2_X1 U835 ( .A(n768), .B(n767), .ZN(n774) );
  XOR2_X1 U836 ( .A(G2427), .B(G2446), .Z(n770) );
  XNOR2_X1 U837 ( .A(G2430), .B(G2451), .ZN(n769) );
  XNOR2_X1 U838 ( .A(n770), .B(n769), .ZN(n772) );
  XOR2_X1 U839 ( .A(G2435), .B(G2438), .Z(n771) );
  XNOR2_X1 U840 ( .A(n772), .B(n771), .ZN(n773) );
  XOR2_X1 U841 ( .A(n774), .B(n773), .Z(n775) );
  AND2_X1 U842 ( .A1(G14), .A2(n775), .ZN(G401) );
  AND2_X1 U843 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U844 ( .A(G57), .ZN(G237) );
  NAND2_X1 U845 ( .A1(G7), .A2(G661), .ZN(n776) );
  XNOR2_X1 U846 ( .A(n776), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U847 ( .A(G223), .ZN(n844) );
  NAND2_X1 U848 ( .A1(n844), .A2(G567), .ZN(n777) );
  XOR2_X1 U849 ( .A(KEYINPUT11), .B(n777), .Z(G234) );
  INV_X1 U850 ( .A(G860), .ZN(n785) );
  BUF_X1 U851 ( .A(n778), .Z(n925) );
  OR2_X1 U852 ( .A1(n785), .A2(n925), .ZN(G153) );
  XNOR2_X1 U853 ( .A(G171), .B(KEYINPUT71), .ZN(G301) );
  NAND2_X1 U854 ( .A1(G868), .A2(G301), .ZN(n779) );
  XNOR2_X1 U855 ( .A(n779), .B(KEYINPUT72), .ZN(n781) );
  INV_X1 U856 ( .A(G868), .ZN(n827) );
  NAND2_X1 U857 ( .A1(n827), .A2(n625), .ZN(n780) );
  NAND2_X1 U858 ( .A1(n781), .A2(n780), .ZN(G284) );
  NOR2_X1 U859 ( .A1(G286), .A2(n827), .ZN(n782) );
  XOR2_X1 U860 ( .A(KEYINPUT75), .B(n782), .Z(n784) );
  NOR2_X1 U861 ( .A1(G868), .A2(G299), .ZN(n783) );
  NOR2_X1 U862 ( .A1(n784), .A2(n783), .ZN(G297) );
  NAND2_X1 U863 ( .A1(n785), .A2(G559), .ZN(n786) );
  NAND2_X1 U864 ( .A1(n786), .A2(n1018), .ZN(n787) );
  XNOR2_X1 U865 ( .A(n787), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U866 ( .A1(n925), .A2(G868), .ZN(n790) );
  NAND2_X1 U867 ( .A1(G868), .A2(n1018), .ZN(n788) );
  NOR2_X1 U868 ( .A1(G559), .A2(n788), .ZN(n789) );
  NOR2_X1 U869 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U870 ( .A(KEYINPUT76), .B(n791), .ZN(G282) );
  NAND2_X1 U871 ( .A1(G123), .A2(n993), .ZN(n792) );
  XOR2_X1 U872 ( .A(KEYINPUT18), .B(n792), .Z(n793) );
  XNOR2_X1 U873 ( .A(n793), .B(KEYINPUT77), .ZN(n795) );
  NAND2_X1 U874 ( .A1(G135), .A2(n708), .ZN(n794) );
  NAND2_X1 U875 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U876 ( .A(KEYINPUT78), .B(n796), .Z(n798) );
  NAND2_X1 U877 ( .A1(n997), .A2(G99), .ZN(n797) );
  NAND2_X1 U878 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U879 ( .A1(G111), .A2(n994), .ZN(n799) );
  XNOR2_X1 U880 ( .A(KEYINPUT79), .B(n799), .ZN(n800) );
  NOR2_X1 U881 ( .A1(n801), .A2(n800), .ZN(n990) );
  XNOR2_X1 U882 ( .A(n990), .B(G2096), .ZN(n803) );
  INV_X1 U883 ( .A(G2100), .ZN(n802) );
  NAND2_X1 U884 ( .A1(n803), .A2(n802), .ZN(G156) );
  NAND2_X1 U885 ( .A1(n1018), .A2(G559), .ZN(n825) );
  XNOR2_X1 U886 ( .A(n925), .B(n825), .ZN(n804) );
  NOR2_X1 U887 ( .A1(G860), .A2(n804), .ZN(n816) );
  NAND2_X1 U888 ( .A1(G93), .A2(n805), .ZN(n808) );
  NAND2_X1 U889 ( .A1(G80), .A2(n806), .ZN(n807) );
  NAND2_X1 U890 ( .A1(n808), .A2(n807), .ZN(n812) );
  NAND2_X1 U891 ( .A1(n809), .A2(G55), .ZN(n810) );
  XOR2_X1 U892 ( .A(KEYINPUT80), .B(n810), .Z(n811) );
  NOR2_X1 U893 ( .A1(n812), .A2(n811), .ZN(n815) );
  NAND2_X1 U894 ( .A1(n813), .A2(G67), .ZN(n814) );
  NAND2_X1 U895 ( .A1(n815), .A2(n814), .ZN(n828) );
  XOR2_X1 U896 ( .A(n816), .B(n828), .Z(G145) );
  XOR2_X1 U897 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n817) );
  XNOR2_X1 U898 ( .A(G305), .B(n817), .ZN(n818) );
  XNOR2_X1 U899 ( .A(G288), .B(n818), .ZN(n821) );
  XNOR2_X1 U900 ( .A(G166), .B(n819), .ZN(n820) );
  XNOR2_X1 U901 ( .A(n821), .B(n820), .ZN(n822) );
  XNOR2_X1 U902 ( .A(n822), .B(G290), .ZN(n823) );
  XNOR2_X1 U903 ( .A(n823), .B(n828), .ZN(n824) );
  XNOR2_X1 U904 ( .A(n925), .B(n824), .ZN(n1021) );
  XNOR2_X1 U905 ( .A(n825), .B(n1021), .ZN(n826) );
  NAND2_X1 U906 ( .A1(n826), .A2(G868), .ZN(n830) );
  NAND2_X1 U907 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U908 ( .A1(n830), .A2(n829), .ZN(G295) );
  NAND2_X1 U909 ( .A1(G2084), .A2(G2078), .ZN(n831) );
  XOR2_X1 U910 ( .A(KEYINPUT20), .B(n831), .Z(n832) );
  NAND2_X1 U911 ( .A1(G2090), .A2(n832), .ZN(n833) );
  XNOR2_X1 U912 ( .A(KEYINPUT21), .B(n833), .ZN(n834) );
  NAND2_X1 U913 ( .A1(n834), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U914 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U915 ( .A(KEYINPUT85), .B(KEYINPUT22), .Z(n836) );
  NAND2_X1 U916 ( .A1(G132), .A2(G82), .ZN(n835) );
  XNOR2_X1 U917 ( .A(n836), .B(n835), .ZN(n837) );
  NOR2_X1 U918 ( .A1(n837), .A2(G218), .ZN(n838) );
  NAND2_X1 U919 ( .A1(G96), .A2(n838), .ZN(n967) );
  NAND2_X1 U920 ( .A1(n967), .A2(G2106), .ZN(n842) );
  NAND2_X1 U921 ( .A1(G69), .A2(G120), .ZN(n839) );
  NOR2_X1 U922 ( .A1(G237), .A2(n839), .ZN(n840) );
  NAND2_X1 U923 ( .A1(G108), .A2(n840), .ZN(n968) );
  NAND2_X1 U924 ( .A1(n968), .A2(G567), .ZN(n841) );
  NAND2_X1 U925 ( .A1(n842), .A2(n841), .ZN(n969) );
  NAND2_X1 U926 ( .A1(G483), .A2(G661), .ZN(n843) );
  NOR2_X1 U927 ( .A1(n969), .A2(n843), .ZN(n847) );
  NAND2_X1 U928 ( .A1(n847), .A2(G36), .ZN(G176) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n844), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n845) );
  NAND2_X1 U931 ( .A1(G661), .A2(n845), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n846) );
  NAND2_X1 U933 ( .A1(n847), .A2(n846), .ZN(G188) );
  NAND2_X1 U935 ( .A1(n994), .A2(G112), .ZN(n854) );
  NAND2_X1 U936 ( .A1(G100), .A2(n997), .ZN(n849) );
  NAND2_X1 U937 ( .A1(G136), .A2(n708), .ZN(n848) );
  NAND2_X1 U938 ( .A1(n849), .A2(n848), .ZN(n852) );
  NAND2_X1 U939 ( .A1(n993), .A2(G124), .ZN(n850) );
  XOR2_X1 U940 ( .A(KEYINPUT44), .B(n850), .Z(n851) );
  NOR2_X1 U941 ( .A1(n852), .A2(n851), .ZN(n853) );
  NAND2_X1 U942 ( .A1(n854), .A2(n853), .ZN(n855) );
  XNOR2_X1 U943 ( .A(n855), .B(KEYINPUT109), .ZN(G162) );
  XOR2_X1 U944 ( .A(G1991), .B(G25), .Z(n856) );
  NAND2_X1 U945 ( .A1(n856), .A2(G28), .ZN(n862) );
  XNOR2_X1 U946 ( .A(n857), .B(G27), .ZN(n859) );
  XNOR2_X1 U947 ( .A(G32), .B(G1996), .ZN(n858) );
  NOR2_X1 U948 ( .A1(n859), .A2(n858), .ZN(n860) );
  XOR2_X1 U949 ( .A(KEYINPUT122), .B(n860), .Z(n861) );
  NOR2_X1 U950 ( .A1(n862), .A2(n861), .ZN(n866) );
  XNOR2_X1 U951 ( .A(G2067), .B(G26), .ZN(n864) );
  XNOR2_X1 U952 ( .A(G33), .B(G2072), .ZN(n863) );
  NOR2_X1 U953 ( .A1(n864), .A2(n863), .ZN(n865) );
  NAND2_X1 U954 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U955 ( .A(n867), .B(KEYINPUT53), .ZN(n870) );
  XOR2_X1 U956 ( .A(G2084), .B(G34), .Z(n868) );
  XNOR2_X1 U957 ( .A(KEYINPUT54), .B(n868), .ZN(n869) );
  NAND2_X1 U958 ( .A1(n870), .A2(n869), .ZN(n873) );
  XOR2_X1 U959 ( .A(G35), .B(G2090), .Z(n871) );
  XNOR2_X1 U960 ( .A(KEYINPUT121), .B(n871), .ZN(n872) );
  NOR2_X1 U961 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U962 ( .A(KEYINPUT55), .B(n874), .ZN(n876) );
  INV_X1 U963 ( .A(G29), .ZN(n875) );
  NAND2_X1 U964 ( .A1(n876), .A2(n875), .ZN(n877) );
  NAND2_X1 U965 ( .A1(n877), .A2(G11), .ZN(n913) );
  NAND2_X1 U966 ( .A1(G103), .A2(n997), .ZN(n879) );
  NAND2_X1 U967 ( .A1(G139), .A2(n708), .ZN(n878) );
  NAND2_X1 U968 ( .A1(n879), .A2(n878), .ZN(n886) );
  XNOR2_X1 U969 ( .A(KEYINPUT47), .B(KEYINPUT112), .ZN(n884) );
  NAND2_X1 U970 ( .A1(G115), .A2(n994), .ZN(n882) );
  NAND2_X1 U971 ( .A1(n993), .A2(G127), .ZN(n880) );
  XOR2_X1 U972 ( .A(KEYINPUT111), .B(n880), .Z(n881) );
  NAND2_X1 U973 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U974 ( .A(n884), .B(n883), .Z(n885) );
  NOR2_X1 U975 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U976 ( .A(KEYINPUT113), .B(n887), .Z(n991) );
  XOR2_X1 U977 ( .A(G2072), .B(n991), .Z(n889) );
  XOR2_X1 U978 ( .A(G164), .B(G2078), .Z(n888) );
  NOR2_X1 U979 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U980 ( .A(n890), .B(KEYINPUT118), .ZN(n891) );
  XNOR2_X1 U981 ( .A(n891), .B(KEYINPUT50), .ZN(n893) );
  NAND2_X1 U982 ( .A1(n893), .A2(n892), .ZN(n898) );
  XOR2_X1 U983 ( .A(G2090), .B(G162), .Z(n894) );
  NOR2_X1 U984 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U985 ( .A(n896), .B(KEYINPUT51), .ZN(n897) );
  NOR2_X1 U986 ( .A1(n898), .A2(n897), .ZN(n905) );
  XOR2_X1 U987 ( .A(G160), .B(G2084), .Z(n899) );
  NOR2_X1 U988 ( .A1(n900), .A2(n899), .ZN(n902) );
  NAND2_X1 U989 ( .A1(n902), .A2(n901), .ZN(n903) );
  NOR2_X1 U990 ( .A1(n903), .A2(n990), .ZN(n904) );
  NAND2_X1 U991 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U992 ( .A(KEYINPUT119), .B(n906), .ZN(n907) );
  XNOR2_X1 U993 ( .A(KEYINPUT52), .B(n907), .ZN(n909) );
  INV_X1 U994 ( .A(KEYINPUT55), .ZN(n908) );
  NAND2_X1 U995 ( .A1(n909), .A2(n908), .ZN(n910) );
  NAND2_X1 U996 ( .A1(n910), .A2(G29), .ZN(n911) );
  XOR2_X1 U997 ( .A(KEYINPUT120), .B(n911), .Z(n912) );
  NOR2_X1 U998 ( .A1(n913), .A2(n912), .ZN(n940) );
  XNOR2_X1 U999 ( .A(G16), .B(KEYINPUT56), .ZN(n938) );
  XNOR2_X1 U1000 ( .A(G171), .B(G1961), .ZN(n915) );
  NAND2_X1 U1001 ( .A1(n915), .A2(n914), .ZN(n931) );
  XNOR2_X1 U1002 ( .A(G299), .B(G1956), .ZN(n923) );
  INV_X1 U1003 ( .A(G1971), .ZN(n916) );
  NOR2_X1 U1004 ( .A1(G166), .A2(n916), .ZN(n920) );
  NAND2_X1 U1005 ( .A1(n918), .A2(n917), .ZN(n919) );
  NOR2_X1 U1006 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1007 ( .A(KEYINPUT123), .B(n921), .ZN(n922) );
  NOR2_X1 U1008 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1009 ( .A(KEYINPUT124), .B(n924), .ZN(n929) );
  XNOR2_X1 U1010 ( .A(n625), .B(G1348), .ZN(n927) );
  XNOR2_X1 U1011 ( .A(G1341), .B(n925), .ZN(n926) );
  NOR2_X1 U1012 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1013 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1014 ( .A1(n931), .A2(n930), .ZN(n936) );
  XOR2_X1 U1015 ( .A(G168), .B(G1966), .Z(n932) );
  NOR2_X1 U1016 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1017 ( .A(KEYINPUT57), .B(n934), .Z(n935) );
  NAND2_X1 U1018 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1019 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1020 ( .A1(n940), .A2(n939), .ZN(n965) );
  XOR2_X1 U1021 ( .A(G1976), .B(G23), .Z(n942) );
  XOR2_X1 U1022 ( .A(G1971), .B(G22), .Z(n941) );
  NAND2_X1 U1023 ( .A1(n942), .A2(n941), .ZN(n944) );
  XNOR2_X1 U1024 ( .A(G24), .B(G1986), .ZN(n943) );
  NOR2_X1 U1025 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1026 ( .A(KEYINPUT58), .B(n945), .Z(n961) );
  XOR2_X1 U1027 ( .A(G1961), .B(G5), .Z(n956) );
  XOR2_X1 U1028 ( .A(G1348), .B(KEYINPUT59), .Z(n946) );
  XNOR2_X1 U1029 ( .A(G4), .B(n946), .ZN(n948) );
  XNOR2_X1 U1030 ( .A(G6), .B(G1981), .ZN(n947) );
  NOR2_X1 U1031 ( .A1(n948), .A2(n947), .ZN(n952) );
  XNOR2_X1 U1032 ( .A(G1341), .B(G19), .ZN(n950) );
  XNOR2_X1 U1033 ( .A(G1956), .B(G20), .ZN(n949) );
  NOR2_X1 U1034 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1035 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1036 ( .A(n953), .B(KEYINPUT125), .ZN(n954) );
  XNOR2_X1 U1037 ( .A(n954), .B(KEYINPUT60), .ZN(n955) );
  NAND2_X1 U1038 ( .A1(n956), .A2(n955), .ZN(n958) );
  XNOR2_X1 U1039 ( .A(G21), .B(G1966), .ZN(n957) );
  NOR2_X1 U1040 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1041 ( .A(KEYINPUT126), .B(n959), .Z(n960) );
  NOR2_X1 U1042 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1043 ( .A(KEYINPUT61), .B(n962), .Z(n963) );
  NOR2_X1 U1044 ( .A1(G16), .A2(n963), .ZN(n964) );
  NOR2_X1 U1045 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1046 ( .A(n966), .B(KEYINPUT62), .ZN(G311) );
  XNOR2_X1 U1047 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1048 ( .A(G132), .ZN(G219) );
  INV_X1 U1049 ( .A(G120), .ZN(G236) );
  INV_X1 U1050 ( .A(G96), .ZN(G221) );
  INV_X1 U1051 ( .A(G82), .ZN(G220) );
  INV_X1 U1052 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1053 ( .A1(n968), .A2(n967), .ZN(G325) );
  INV_X1 U1054 ( .A(G325), .ZN(G261) );
  INV_X1 U1055 ( .A(n969), .ZN(G319) );
  XOR2_X1 U1056 ( .A(G2678), .B(KEYINPUT42), .Z(n971) );
  XNOR2_X1 U1057 ( .A(G2096), .B(G2100), .ZN(n970) );
  XNOR2_X1 U1058 ( .A(n971), .B(n970), .ZN(n975) );
  XOR2_X1 U1059 ( .A(KEYINPUT43), .B(G2072), .Z(n973) );
  XNOR2_X1 U1060 ( .A(G2090), .B(G2067), .ZN(n972) );
  XNOR2_X1 U1061 ( .A(n973), .B(n972), .ZN(n974) );
  XOR2_X1 U1062 ( .A(n975), .B(n974), .Z(n977) );
  XNOR2_X1 U1063 ( .A(G2084), .B(G2078), .ZN(n976) );
  XNOR2_X1 U1064 ( .A(n977), .B(n976), .ZN(G227) );
  XOR2_X1 U1065 ( .A(G2474), .B(KEYINPUT106), .Z(n979) );
  XNOR2_X1 U1066 ( .A(G1966), .B(G1961), .ZN(n978) );
  XNOR2_X1 U1067 ( .A(n979), .B(n978), .ZN(n989) );
  XOR2_X1 U1068 ( .A(KEYINPUT107), .B(KEYINPUT41), .Z(n981) );
  XNOR2_X1 U1069 ( .A(G1986), .B(G1991), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(n981), .B(n980), .ZN(n985) );
  XOR2_X1 U1071 ( .A(G1976), .B(G1981), .Z(n983) );
  XNOR2_X1 U1072 ( .A(G1956), .B(G1971), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(n983), .B(n982), .ZN(n984) );
  XOR2_X1 U1074 ( .A(n985), .B(n984), .Z(n987) );
  XNOR2_X1 U1075 ( .A(G1996), .B(KEYINPUT108), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(n987), .B(n986), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(n989), .B(n988), .ZN(G229) );
  XNOR2_X1 U1078 ( .A(G160), .B(n990), .ZN(n1014) );
  XNOR2_X1 U1079 ( .A(n992), .B(n991), .ZN(n1005) );
  NAND2_X1 U1080 ( .A1(G130), .A2(n993), .ZN(n996) );
  NAND2_X1 U1081 ( .A1(G118), .A2(n994), .ZN(n995) );
  NAND2_X1 U1082 ( .A1(n996), .A2(n995), .ZN(n1003) );
  NAND2_X1 U1083 ( .A1(G106), .A2(n997), .ZN(n999) );
  NAND2_X1 U1084 ( .A1(G142), .A2(n708), .ZN(n998) );
  NAND2_X1 U1085 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1086 ( .A(KEYINPUT45), .B(n1000), .Z(n1001) );
  XNOR2_X1 U1087 ( .A(KEYINPUT110), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1088 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1089 ( .A(n1005), .B(n1004), .ZN(n1010) );
  XNOR2_X1 U1090 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n1008) );
  XNOR2_X1 U1091 ( .A(n1006), .B(KEYINPUT114), .ZN(n1007) );
  XNOR2_X1 U1092 ( .A(n1008), .B(n1007), .ZN(n1009) );
  XOR2_X1 U1093 ( .A(n1010), .B(n1009), .Z(n1012) );
  XNOR2_X1 U1094 ( .A(G164), .B(G162), .ZN(n1011) );
  XNOR2_X1 U1095 ( .A(n1012), .B(n1011), .ZN(n1013) );
  XNOR2_X1 U1096 ( .A(n1014), .B(n1013), .ZN(n1016) );
  XOR2_X1 U1097 ( .A(n1016), .B(n1015), .Z(n1017) );
  NOR2_X1 U1098 ( .A1(G37), .A2(n1017), .ZN(G395) );
  XNOR2_X1 U1099 ( .A(G286), .B(KEYINPUT115), .ZN(n1020) );
  XNOR2_X1 U1100 ( .A(G171), .B(n1018), .ZN(n1019) );
  XNOR2_X1 U1101 ( .A(n1020), .B(n1019), .ZN(n1022) );
  XNOR2_X1 U1102 ( .A(n1022), .B(n1021), .ZN(n1023) );
  NOR2_X1 U1103 ( .A1(G37), .A2(n1023), .ZN(n1024) );
  XNOR2_X1 U1104 ( .A(KEYINPUT116), .B(n1024), .ZN(G397) );
  NOR2_X1 U1105 ( .A1(G227), .A2(G229), .ZN(n1025) );
  XNOR2_X1 U1106 ( .A(n1025), .B(KEYINPUT49), .ZN(n1026) );
  NOR2_X1 U1107 ( .A1(G401), .A2(n1026), .ZN(n1027) );
  NAND2_X1 U1108 ( .A1(G319), .A2(n1027), .ZN(n1028) );
  XNOR2_X1 U1109 ( .A(KEYINPUT117), .B(n1028), .ZN(n1030) );
  NOR2_X1 U1110 ( .A1(G395), .A2(G397), .ZN(n1029) );
  NAND2_X1 U1111 ( .A1(n1030), .A2(n1029), .ZN(G225) );
  INV_X1 U1112 ( .A(G225), .ZN(G308) );
  INV_X1 U1113 ( .A(G108), .ZN(G238) );
endmodule

