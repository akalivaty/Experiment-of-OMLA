

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718;

  INV_X1 U363 ( .A(G953), .ZN(n707) );
  AND2_X2 U364 ( .A1(n589), .A2(n468), .ZN(n375) );
  OR2_X2 U365 ( .A1(n636), .A2(n504), .ZN(n505) );
  OR2_X2 U366 ( .A1(n610), .A2(G902), .ZN(n368) );
  XNOR2_X2 U367 ( .A(n435), .B(n434), .ZN(n555) );
  OR2_X1 U368 ( .A1(n549), .A2(n548), .ZN(n552) );
  NOR2_X1 U369 ( .A1(n662), .A2(n660), .ZN(n481) );
  NOR2_X1 U370 ( .A1(n705), .A2(KEYINPUT83), .ZN(n582) );
  NAND2_X1 U371 ( .A1(n488), .A2(n532), .ZN(n634) );
  NAND2_X1 U372 ( .A1(n364), .A2(n361), .ZN(n532) );
  XNOR2_X1 U373 ( .A(n345), .B(n395), .ZN(n461) );
  XNOR2_X1 U374 ( .A(G143), .B(KEYINPUT65), .ZN(n345) );
  XNOR2_X1 U375 ( .A(G101), .B(KEYINPUT90), .ZN(n411) );
  OR2_X2 U376 ( .A1(n644), .A2(n555), .ZN(n436) );
  BUF_X2 U377 ( .A(n647), .Z(n339) );
  XNOR2_X1 U378 ( .A(n448), .B(n371), .ZN(n647) );
  INV_X1 U379 ( .A(KEYINPUT46), .ZN(n483) );
  XNOR2_X1 U380 ( .A(n373), .B(n372), .ZN(n347) );
  INV_X1 U381 ( .A(KEYINPUT77), .ZN(n372) );
  NOR2_X1 U382 ( .A1(n498), .A2(n497), .ZN(n373) );
  XNOR2_X1 U383 ( .A(n438), .B(n437), .ZN(n699) );
  XOR2_X1 U384 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n379) );
  INV_X1 U385 ( .A(KEYINPUT78), .ZN(n522) );
  NAND2_X1 U386 ( .A1(n521), .A2(n642), .ZN(n354) );
  XNOR2_X1 U387 ( .A(n461), .B(G134), .ZN(n408) );
  XNOR2_X1 U388 ( .A(n408), .B(G131), .ZN(n438) );
  XNOR2_X1 U389 ( .A(n460), .B(n356), .ZN(n437) );
  INV_X1 U390 ( .A(G137), .ZN(n356) );
  XNOR2_X1 U391 ( .A(n360), .B(n410), .ZN(n458) );
  XNOR2_X1 U392 ( .A(G107), .B(G104), .ZN(n410) );
  XNOR2_X1 U393 ( .A(n411), .B(n409), .ZN(n360) );
  INV_X1 U394 ( .A(G110), .ZN(n409) );
  XNOR2_X1 U395 ( .A(n476), .B(n475), .ZN(n516) );
  AND2_X1 U396 ( .A1(n369), .A2(n479), .ZN(n480) );
  AND2_X1 U397 ( .A1(n503), .A2(n647), .ZN(n370) );
  XNOR2_X1 U398 ( .A(n406), .B(G478), .ZN(n493) );
  NAND2_X1 U399 ( .A1(n532), .A2(n531), .ZN(n533) );
  INV_X1 U400 ( .A(G237), .ZN(n449) );
  INV_X1 U401 ( .A(G902), .ZN(n450) );
  NOR2_X1 U402 ( .A1(G953), .A2(G237), .ZN(n439) );
  NAND2_X1 U403 ( .A1(G234), .A2(G237), .ZN(n452) );
  XNOR2_X1 U404 ( .A(n346), .B(n342), .ZN(n587) );
  NOR2_X1 U405 ( .A1(n499), .A2(n374), .ZN(n348) );
  INV_X1 U406 ( .A(n477), .ZN(n352) );
  NAND2_X1 U407 ( .A1(n486), .A2(n487), .ZN(n365) );
  XNOR2_X1 U408 ( .A(G128), .B(G137), .ZN(n421) );
  XOR2_X1 U409 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n397) );
  XNOR2_X1 U410 ( .A(G116), .B(G107), .ZN(n399) );
  INV_X1 U411 ( .A(G146), .ZN(n380) );
  INV_X1 U412 ( .A(G128), .ZN(n395) );
  INV_X1 U413 ( .A(KEYINPUT1), .ZN(n367) );
  AND2_X1 U414 ( .A1(n351), .A2(n349), .ZN(n495) );
  XNOR2_X1 U415 ( .A(n350), .B(n451), .ZN(n349) );
  NOR2_X1 U416 ( .A1(n543), .A2(n352), .ZN(n351) );
  INV_X1 U417 ( .A(KEYINPUT30), .ZN(n451) );
  NAND2_X1 U418 ( .A1(n363), .A2(n362), .ZN(n361) );
  AND2_X1 U419 ( .A1(n366), .A2(n365), .ZN(n364) );
  NOR2_X1 U420 ( .A1(n486), .A2(n487), .ZN(n362) );
  NOR2_X1 U421 ( .A1(n591), .A2(G902), .ZN(n448) );
  XNOR2_X1 U422 ( .A(n359), .B(n459), .ZN(n694) );
  XNOR2_X1 U423 ( .A(n458), .B(n457), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n438), .B(n355), .ZN(n610) );
  XNOR2_X1 U425 ( .A(n357), .B(n437), .ZN(n355) );
  XNOR2_X1 U426 ( .A(n458), .B(n413), .ZN(n357) );
  XNOR2_X1 U427 ( .A(n353), .B(n341), .ZN(n718) );
  XNOR2_X1 U428 ( .A(KEYINPUT74), .B(KEYINPUT34), .ZN(n534) );
  INV_X1 U429 ( .A(n521), .ZN(n520) );
  XOR2_X1 U430 ( .A(n416), .B(n415), .Z(n340) );
  XOR2_X1 U431 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n341) );
  XOR2_X1 U432 ( .A(KEYINPUT87), .B(KEYINPUT48), .Z(n342) );
  XNOR2_X1 U433 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n343) );
  XOR2_X1 U434 ( .A(n591), .B(KEYINPUT62), .Z(n344) );
  XNOR2_X1 U435 ( .A(KEYINPUT15), .B(G902), .ZN(n590) );
  OR2_X2 U436 ( .A1(n553), .A2(n505), .ZN(n510) );
  INV_X1 U437 ( .A(n587), .ZN(n519) );
  NAND2_X1 U438 ( .A1(n348), .A2(n347), .ZN(n346) );
  NAND2_X1 U439 ( .A1(n339), .A2(n657), .ZN(n350) );
  NOR2_X1 U440 ( .A1(n718), .A2(n717), .ZN(n484) );
  NAND2_X1 U441 ( .A1(n516), .A2(n490), .ZN(n353) );
  XNOR2_X1 U442 ( .A(n540), .B(KEYINPUT104), .ZN(n524) );
  XNOR2_X2 U443 ( .A(n354), .B(n522), .ZN(n540) );
  XNOR2_X2 U444 ( .A(n500), .B(n367), .ZN(n521) );
  INV_X1 U445 ( .A(n358), .ZN(n686) );
  NAND2_X1 U446 ( .A1(n358), .A2(n588), .ZN(n589) );
  XNOR2_X2 U447 ( .A(n581), .B(n343), .ZN(n358) );
  NAND2_X1 U448 ( .A1(n358), .A2(n582), .ZN(n377) );
  INV_X1 U449 ( .A(n513), .ZN(n363) );
  NAND2_X1 U450 ( .A1(n513), .A2(n487), .ZN(n366) );
  XNOR2_X2 U451 ( .A(n473), .B(n472), .ZN(n513) );
  NAND2_X1 U452 ( .A1(n561), .A2(n573), .ZN(n571) );
  NAND2_X1 U453 ( .A1(n598), .A2(n570), .ZN(n573) );
  XNOR2_X2 U454 ( .A(n368), .B(n340), .ZN(n500) );
  XNOR2_X1 U455 ( .A(n370), .B(KEYINPUT28), .ZN(n369) );
  INV_X1 U456 ( .A(G472), .ZN(n371) );
  INV_X1 U457 ( .A(n712), .ZN(n374) );
  NAND2_X1 U458 ( .A1(n376), .A2(n589), .ZN(n676) );
  AND2_X4 U459 ( .A1(n376), .A2(n375), .ZN(n679) );
  NAND2_X2 U460 ( .A1(n377), .A2(n583), .ZN(n376) );
  XNOR2_X1 U461 ( .A(n484), .B(n483), .ZN(n499) );
  INV_X1 U462 ( .A(n553), .ZN(n523) );
  XNOR2_X1 U463 ( .A(n424), .B(n423), .ZN(n425) );
  INV_X1 U464 ( .A(KEYINPUT33), .ZN(n525) );
  XNOR2_X1 U465 ( .A(n699), .B(n447), .ZN(n591) );
  XNOR2_X1 U466 ( .A(n426), .B(n425), .ZN(n427) );
  INV_X1 U467 ( .A(n500), .ZN(n479) );
  INV_X1 U468 ( .A(KEYINPUT73), .ZN(n474) );
  XNOR2_X1 U469 ( .A(n474), .B(KEYINPUT39), .ZN(n475) );
  INV_X1 U470 ( .A(n683), .ZN(n594) );
  XNOR2_X1 U471 ( .A(G125), .B(G140), .ZN(n378) );
  XNOR2_X1 U472 ( .A(n379), .B(n378), .ZN(n698) );
  XNOR2_X1 U473 ( .A(n698), .B(n380), .ZN(n428) );
  XOR2_X1 U474 ( .A(G104), .B(G113), .Z(n382) );
  XNOR2_X1 U475 ( .A(G143), .B(G131), .ZN(n381) );
  XNOR2_X1 U476 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U477 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n384) );
  XNOR2_X1 U478 ( .A(G122), .B(KEYINPUT96), .ZN(n383) );
  XNOR2_X1 U479 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U480 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U481 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n388) );
  NAND2_X1 U482 ( .A1(G214), .A2(n439), .ZN(n387) );
  XNOR2_X1 U483 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U484 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U485 ( .A(n428), .B(n391), .ZN(n604) );
  NOR2_X1 U486 ( .A1(G902), .A2(n604), .ZN(n393) );
  XNOR2_X1 U487 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n392) );
  XNOR2_X1 U488 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U489 ( .A(n394), .B(G475), .ZN(n494) );
  INV_X1 U490 ( .A(n494), .ZN(n407) );
  XNOR2_X1 U491 ( .A(G122), .B(KEYINPUT100), .ZN(n396) );
  XNOR2_X1 U492 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U493 ( .A(n398), .B(KEYINPUT101), .Z(n400) );
  XNOR2_X1 U494 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U495 ( .A(n408), .B(n401), .Z(n405) );
  XOR2_X1 U496 ( .A(KEYINPUT86), .B(KEYINPUT8), .Z(n403) );
  NAND2_X1 U497 ( .A1(G234), .A2(n707), .ZN(n402) );
  XNOR2_X1 U498 ( .A(n403), .B(n402), .ZN(n420) );
  NAND2_X1 U499 ( .A1(G217), .A2(n420), .ZN(n404) );
  XNOR2_X1 U500 ( .A(n405), .B(n404), .ZN(n680) );
  NOR2_X1 U501 ( .A1(n680), .A2(G902), .ZN(n406) );
  NAND2_X1 U502 ( .A1(n407), .A2(n493), .ZN(n636) );
  INV_X1 U503 ( .A(n636), .ZN(n490) );
  NAND2_X1 U504 ( .A1(G227), .A2(n707), .ZN(n412) );
  XOR2_X1 U505 ( .A(G140), .B(n412), .Z(n413) );
  XNOR2_X1 U506 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n414) );
  XNOR2_X1 U507 ( .A(n414), .B(G146), .ZN(n460) );
  XNOR2_X1 U508 ( .A(KEYINPUT71), .B(KEYINPUT70), .ZN(n416) );
  INV_X1 U509 ( .A(G469), .ZN(n415) );
  NAND2_X1 U510 ( .A1(G234), .A2(n590), .ZN(n417) );
  XNOR2_X1 U511 ( .A(KEYINPUT20), .B(n417), .ZN(n429) );
  AND2_X1 U512 ( .A1(n429), .A2(G221), .ZN(n419) );
  INV_X1 U513 ( .A(KEYINPUT21), .ZN(n418) );
  XNOR2_X1 U514 ( .A(n419), .B(n418), .ZN(n644) );
  NAND2_X1 U515 ( .A1(G221), .A2(n420), .ZN(n426) );
  XOR2_X1 U516 ( .A(G110), .B(G119), .Z(n422) );
  XNOR2_X1 U517 ( .A(n422), .B(n421), .ZN(n424) );
  XOR2_X1 U518 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n423) );
  XNOR2_X1 U519 ( .A(n428), .B(n427), .ZN(n599) );
  NAND2_X1 U520 ( .A1(n599), .A2(n450), .ZN(n435) );
  AND2_X1 U521 ( .A1(n429), .A2(G217), .ZN(n431) );
  XNOR2_X1 U522 ( .A(KEYINPUT95), .B(KEYINPUT25), .ZN(n430) );
  XNOR2_X1 U523 ( .A(n431), .B(n430), .ZN(n433) );
  XOR2_X1 U524 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n432) );
  XNOR2_X1 U525 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X2 U526 ( .A(n436), .B(KEYINPUT67), .ZN(n642) );
  NAND2_X1 U527 ( .A1(n479), .A2(n642), .ZN(n543) );
  XOR2_X1 U528 ( .A(KEYINPUT79), .B(KEYINPUT5), .Z(n442) );
  NAND2_X1 U529 ( .A1(n439), .A2(G210), .ZN(n440) );
  XNOR2_X1 U530 ( .A(n440), .B(G101), .ZN(n441) );
  XOR2_X1 U531 ( .A(n442), .B(n441), .Z(n446) );
  XNOR2_X1 U532 ( .A(G119), .B(G116), .ZN(n443) );
  XNOR2_X1 U533 ( .A(n443), .B(KEYINPUT3), .ZN(n445) );
  XNOR2_X1 U534 ( .A(G113), .B(KEYINPUT72), .ZN(n444) );
  XNOR2_X1 U535 ( .A(n445), .B(n444), .ZN(n459) );
  XNOR2_X1 U536 ( .A(n446), .B(n459), .ZN(n447) );
  NAND2_X1 U537 ( .A1(n450), .A2(n449), .ZN(n469) );
  NAND2_X1 U538 ( .A1(n469), .A2(G214), .ZN(n657) );
  XNOR2_X1 U539 ( .A(n452), .B(KEYINPUT14), .ZN(n454) );
  NAND2_X1 U540 ( .A1(G952), .A2(n454), .ZN(n453) );
  XOR2_X1 U541 ( .A(KEYINPUT92), .B(n453), .Z(n669) );
  NAND2_X1 U542 ( .A1(n707), .A2(n669), .ZN(n529) );
  NAND2_X1 U543 ( .A1(G902), .A2(n454), .ZN(n527) );
  NOR2_X1 U544 ( .A1(G900), .A2(n527), .ZN(n455) );
  NAND2_X1 U545 ( .A1(G953), .A2(n455), .ZN(n456) );
  NAND2_X1 U546 ( .A1(n529), .A2(n456), .ZN(n477) );
  XNOR2_X1 U547 ( .A(KEYINPUT16), .B(G122), .ZN(n457) );
  XNOR2_X1 U548 ( .A(n461), .B(n460), .ZN(n466) );
  XOR2_X1 U549 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n464) );
  NAND2_X1 U550 ( .A1(G224), .A2(n707), .ZN(n462) );
  XNOR2_X1 U551 ( .A(n462), .B(G125), .ZN(n463) );
  XNOR2_X1 U552 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U553 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U554 ( .A(n694), .B(n467), .ZN(n617) );
  INV_X1 U555 ( .A(n590), .ZN(n468) );
  OR2_X1 U556 ( .A1(n617), .A2(n468), .ZN(n473) );
  NAND2_X1 U557 ( .A1(n469), .A2(G210), .ZN(n471) );
  INV_X1 U558 ( .A(KEYINPUT91), .ZN(n470) );
  XNOR2_X1 U559 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U560 ( .A(n513), .B(KEYINPUT38), .ZN(n658) );
  NAND2_X1 U561 ( .A1(n495), .A2(n658), .ZN(n476) );
  NAND2_X1 U562 ( .A1(n555), .A2(n477), .ZN(n478) );
  NOR2_X1 U563 ( .A1(n644), .A2(n478), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n480), .B(KEYINPUT107), .ZN(n485) );
  NAND2_X1 U565 ( .A1(n658), .A2(n657), .ZN(n662) );
  NAND2_X1 U566 ( .A1(n493), .A2(n494), .ZN(n660) );
  XNOR2_X1 U567 ( .A(n481), .B(KEYINPUT41), .ZN(n672) );
  NOR2_X1 U568 ( .A1(n485), .A2(n672), .ZN(n482) );
  XNOR2_X1 U569 ( .A(KEYINPUT42), .B(n482), .ZN(n717) );
  INV_X1 U570 ( .A(n485), .ZN(n488) );
  INV_X1 U571 ( .A(n657), .ZN(n486) );
  XNOR2_X1 U572 ( .A(KEYINPUT80), .B(KEYINPUT19), .ZN(n487) );
  INV_X1 U573 ( .A(n493), .ZN(n489) );
  AND2_X1 U574 ( .A1(n489), .A2(n494), .ZN(n626) );
  NOR2_X1 U575 ( .A1(n626), .A2(n490), .ZN(n491) );
  XNOR2_X1 U576 ( .A(n491), .B(KEYINPUT102), .ZN(n661) );
  NOR2_X1 U577 ( .A1(n634), .A2(n661), .ZN(n492) );
  XOR2_X1 U578 ( .A(KEYINPUT47), .B(n492), .Z(n498) );
  NOR2_X1 U579 ( .A1(n494), .A2(n493), .ZN(n536) );
  NAND2_X1 U580 ( .A1(n495), .A2(n536), .ZN(n496) );
  NOR2_X1 U581 ( .A1(n496), .A2(n513), .ZN(n597) );
  XOR2_X1 U582 ( .A(KEYINPUT85), .B(n597), .Z(n497) );
  INV_X1 U583 ( .A(KEYINPUT103), .ZN(n501) );
  XNOR2_X1 U584 ( .A(n501), .B(KEYINPUT6), .ZN(n502) );
  XNOR2_X1 U585 ( .A(n339), .B(n502), .ZN(n553) );
  NAND2_X1 U586 ( .A1(n503), .A2(n657), .ZN(n504) );
  NOR2_X1 U587 ( .A1(n510), .A2(n513), .ZN(n507) );
  XNOR2_X1 U588 ( .A(KEYINPUT36), .B(KEYINPUT89), .ZN(n506) );
  XNOR2_X1 U589 ( .A(n507), .B(n506), .ZN(n508) );
  NOR2_X1 U590 ( .A1(n520), .A2(n508), .ZN(n509) );
  XNOR2_X1 U591 ( .A(n509), .B(KEYINPUT109), .ZN(n712) );
  XOR2_X1 U592 ( .A(n510), .B(KEYINPUT105), .Z(n511) );
  NOR2_X1 U593 ( .A1(n521), .A2(n511), .ZN(n512) );
  XNOR2_X1 U594 ( .A(n512), .B(KEYINPUT43), .ZN(n514) );
  NOR2_X1 U595 ( .A1(n514), .A2(n363), .ZN(n515) );
  XNOR2_X1 U596 ( .A(n515), .B(KEYINPUT106), .ZN(n715) );
  NAND2_X1 U597 ( .A1(n626), .A2(n516), .ZN(n641) );
  INV_X1 U598 ( .A(n641), .ZN(n517) );
  NOR2_X1 U599 ( .A1(n715), .A2(n517), .ZN(n518) );
  NAND2_X1 U600 ( .A1(n519), .A2(n518), .ZN(n705) );
  NAND2_X1 U601 ( .A1(n524), .A2(n523), .ZN(n526) );
  XNOR2_X2 U602 ( .A(n526), .B(n525), .ZN(n671) );
  XNOR2_X1 U603 ( .A(G898), .B(KEYINPUT93), .ZN(n690) );
  NAND2_X1 U604 ( .A1(G953), .A2(n690), .ZN(n693) );
  OR2_X1 U605 ( .A1(n527), .A2(n693), .ZN(n528) );
  NAND2_X1 U606 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U607 ( .A(n530), .B(KEYINPUT94), .ZN(n531) );
  XNOR2_X2 U608 ( .A(n533), .B(KEYINPUT0), .ZN(n549) );
  NOR2_X2 U609 ( .A1(n671), .A2(n549), .ZN(n535) );
  XNOR2_X1 U610 ( .A(n535), .B(n534), .ZN(n537) );
  NAND2_X1 U611 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X2 U612 ( .A(n538), .B(KEYINPUT35), .ZN(n713) );
  INV_X1 U613 ( .A(n713), .ZN(n539) );
  NAND2_X1 U614 ( .A1(n539), .A2(n576), .ZN(n560) );
  NAND2_X1 U615 ( .A1(n339), .A2(n540), .ZN(n652) );
  OR2_X1 U616 ( .A1(n652), .A2(n549), .ZN(n542) );
  INV_X1 U617 ( .A(KEYINPUT31), .ZN(n541) );
  XNOR2_X1 U618 ( .A(n542), .B(n541), .ZN(n638) );
  NOR2_X1 U619 ( .A1(n543), .A2(n339), .ZN(n545) );
  INV_X1 U620 ( .A(n549), .ZN(n544) );
  NAND2_X1 U621 ( .A1(n545), .A2(n544), .ZN(n627) );
  NAND2_X1 U622 ( .A1(n638), .A2(n627), .ZN(n547) );
  INV_X1 U623 ( .A(n661), .ZN(n546) );
  NAND2_X1 U624 ( .A1(n547), .A2(n546), .ZN(n558) );
  OR2_X1 U625 ( .A1(n660), .A2(n644), .ZN(n548) );
  XNOR2_X1 U626 ( .A(KEYINPUT76), .B(KEYINPUT22), .ZN(n550) );
  XNOR2_X1 U627 ( .A(n550), .B(KEYINPUT75), .ZN(n551) );
  XNOR2_X1 U628 ( .A(n552), .B(n551), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n568), .A2(n553), .ZN(n562) );
  INV_X1 U630 ( .A(KEYINPUT88), .ZN(n554) );
  XNOR2_X1 U631 ( .A(n562), .B(n554), .ZN(n557) );
  INV_X1 U632 ( .A(n555), .ZN(n566) );
  AND2_X1 U633 ( .A1(n520), .A2(n566), .ZN(n556) );
  NAND2_X1 U634 ( .A1(n557), .A2(n556), .ZN(n622) );
  AND2_X1 U635 ( .A1(n558), .A2(n622), .ZN(n561) );
  AND2_X1 U636 ( .A1(KEYINPUT66), .A2(n561), .ZN(n559) );
  NAND2_X1 U637 ( .A1(n560), .A2(n559), .ZN(n572) );
  INV_X1 U638 ( .A(n562), .ZN(n564) );
  NOR2_X1 U639 ( .A1(n520), .A2(n566), .ZN(n563) );
  NAND2_X1 U640 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U641 ( .A(n565), .B(KEYINPUT32), .ZN(n598) );
  NOR2_X1 U642 ( .A1(n339), .A2(n566), .ZN(n567) );
  AND2_X1 U643 ( .A1(n520), .A2(n567), .ZN(n569) );
  AND2_X1 U644 ( .A1(n569), .A2(n568), .ZN(n630) );
  INV_X1 U645 ( .A(n630), .ZN(n570) );
  NAND2_X1 U646 ( .A1(n572), .A2(n571), .ZN(n580) );
  NAND2_X1 U647 ( .A1(n573), .A2(KEYINPUT66), .ZN(n575) );
  INV_X1 U648 ( .A(KEYINPUT44), .ZN(n576) );
  NOR2_X1 U649 ( .A1(n713), .A2(n576), .ZN(n574) );
  NAND2_X1 U650 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U651 ( .A1(n576), .A2(KEYINPUT66), .ZN(n577) );
  NAND2_X1 U652 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U653 ( .A1(n580), .A2(n579), .ZN(n581) );
  INV_X1 U654 ( .A(KEYINPUT2), .ZN(n583) );
  XOR2_X1 U655 ( .A(n641), .B(KEYINPUT83), .Z(n584) );
  NAND2_X1 U656 ( .A1(KEYINPUT2), .A2(n584), .ZN(n585) );
  OR2_X1 U657 ( .A1(n715), .A2(n585), .ZN(n586) );
  NOR2_X1 U658 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n679), .A2(G472), .ZN(n592) );
  XNOR2_X1 U660 ( .A(n592), .B(n344), .ZN(n595) );
  INV_X1 U661 ( .A(G952), .ZN(n593) );
  AND2_X1 U662 ( .A1(n593), .A2(G953), .ZN(n683) );
  NAND2_X1 U663 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U664 ( .A(n596), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U665 ( .A(G143), .B(n597), .Z(G45) );
  XNOR2_X1 U666 ( .A(n598), .B(G119), .ZN(G21) );
  NAND2_X1 U667 ( .A1(n679), .A2(G217), .ZN(n601) );
  XNOR2_X1 U668 ( .A(n599), .B(KEYINPUT119), .ZN(n600) );
  XNOR2_X1 U669 ( .A(n601), .B(n600), .ZN(n602) );
  NOR2_X2 U670 ( .A1(n602), .A2(n683), .ZN(n603) );
  XNOR2_X1 U671 ( .A(n603), .B(KEYINPUT120), .ZN(G66) );
  NAND2_X1 U672 ( .A1(n679), .A2(G475), .ZN(n606) );
  XOR2_X1 U673 ( .A(n604), .B(KEYINPUT59), .Z(n605) );
  XNOR2_X1 U674 ( .A(n606), .B(n605), .ZN(n607) );
  NOR2_X2 U675 ( .A1(n607), .A2(n683), .ZN(n608) );
  XNOR2_X1 U676 ( .A(n608), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U677 ( .A1(n679), .A2(G469), .ZN(n612) );
  XOR2_X1 U678 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n609) );
  XNOR2_X1 U679 ( .A(n610), .B(n609), .ZN(n611) );
  XNOR2_X1 U680 ( .A(n612), .B(n611), .ZN(n613) );
  NOR2_X2 U681 ( .A1(n613), .A2(n683), .ZN(n614) );
  XNOR2_X1 U682 ( .A(n614), .B(KEYINPUT116), .ZN(G54) );
  NAND2_X1 U683 ( .A1(n679), .A2(G210), .ZN(n619) );
  XNOR2_X1 U684 ( .A(KEYINPUT84), .B(KEYINPUT54), .ZN(n615) );
  XOR2_X1 U685 ( .A(n615), .B(KEYINPUT55), .Z(n616) );
  XNOR2_X1 U686 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U687 ( .A(n619), .B(n618), .ZN(n620) );
  NOR2_X2 U688 ( .A1(n620), .A2(n683), .ZN(n621) );
  XNOR2_X1 U689 ( .A(n621), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U690 ( .A(G101), .B(n622), .ZN(G3) );
  NOR2_X1 U691 ( .A1(n636), .A2(n627), .ZN(n623) );
  XOR2_X1 U692 ( .A(G104), .B(n623), .Z(G6) );
  XOR2_X1 U693 ( .A(KEYINPUT110), .B(KEYINPUT26), .Z(n625) );
  XNOR2_X1 U694 ( .A(G107), .B(KEYINPUT27), .ZN(n624) );
  XNOR2_X1 U695 ( .A(n625), .B(n624), .ZN(n629) );
  INV_X1 U696 ( .A(n626), .ZN(n639) );
  NOR2_X1 U697 ( .A1(n639), .A2(n627), .ZN(n628) );
  XOR2_X1 U698 ( .A(n629), .B(n628), .Z(G9) );
  XNOR2_X1 U699 ( .A(G110), .B(n630), .ZN(n631) );
  XNOR2_X1 U700 ( .A(n631), .B(KEYINPUT111), .ZN(G12) );
  NOR2_X1 U701 ( .A1(n634), .A2(n639), .ZN(n633) );
  XNOR2_X1 U702 ( .A(G128), .B(KEYINPUT29), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n633), .B(n632), .ZN(G30) );
  NOR2_X1 U704 ( .A1(n634), .A2(n636), .ZN(n635) );
  XOR2_X1 U705 ( .A(G146), .B(n635), .Z(G48) );
  NOR2_X1 U706 ( .A1(n636), .A2(n638), .ZN(n637) );
  XOR2_X1 U707 ( .A(G113), .B(n637), .Z(G15) );
  NOR2_X1 U708 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U709 ( .A(G116), .B(n640), .Z(G18) );
  XNOR2_X1 U710 ( .A(G134), .B(n641), .ZN(G36) );
  XNOR2_X1 U711 ( .A(KEYINPUT51), .B(KEYINPUT114), .ZN(n654) );
  NOR2_X1 U712 ( .A1(n521), .A2(n642), .ZN(n643) );
  XOR2_X1 U713 ( .A(KEYINPUT50), .B(n643), .Z(n650) );
  XOR2_X1 U714 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n646) );
  NAND2_X1 U715 ( .A1(n644), .A2(n555), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n646), .B(n645), .ZN(n648) );
  NOR2_X1 U717 ( .A1(n648), .A2(n339), .ZN(n649) );
  NAND2_X1 U718 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U719 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U720 ( .A(n654), .B(n653), .ZN(n655) );
  NOR2_X1 U721 ( .A1(n672), .A2(n655), .ZN(n656) );
  XOR2_X1 U722 ( .A(KEYINPUT115), .B(n656), .Z(n667) );
  NOR2_X1 U723 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U724 ( .A1(n660), .A2(n659), .ZN(n664) );
  NOR2_X1 U725 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U726 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U727 ( .A1(n665), .A2(n671), .ZN(n666) );
  NOR2_X1 U728 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U729 ( .A(KEYINPUT52), .B(n668), .Z(n670) );
  AND2_X1 U730 ( .A1(n670), .A2(n669), .ZN(n674) );
  NOR2_X1 U731 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U732 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U733 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U734 ( .A1(n707), .A2(n677), .ZN(n678) );
  XOR2_X1 U735 ( .A(KEYINPUT53), .B(n678), .Z(G75) );
  NAND2_X1 U736 ( .A1(n679), .A2(G478), .ZN(n682) );
  XOR2_X1 U737 ( .A(n680), .B(KEYINPUT117), .Z(n681) );
  XNOR2_X1 U738 ( .A(n682), .B(n681), .ZN(n684) );
  NOR2_X2 U739 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U740 ( .A(n685), .B(KEYINPUT118), .ZN(G63) );
  NOR2_X1 U741 ( .A1(n686), .A2(G953), .ZN(n692) );
  NAND2_X1 U742 ( .A1(G224), .A2(G953), .ZN(n687) );
  XNOR2_X1 U743 ( .A(n687), .B(KEYINPUT61), .ZN(n688) );
  XNOR2_X1 U744 ( .A(n688), .B(KEYINPUT121), .ZN(n689) );
  NOR2_X1 U745 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U746 ( .A1(n692), .A2(n691), .ZN(n697) );
  NAND2_X1 U747 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U748 ( .A(n695), .B(KEYINPUT122), .ZN(n696) );
  XNOR2_X1 U749 ( .A(n697), .B(n696), .ZN(G69) );
  XOR2_X1 U750 ( .A(n699), .B(n698), .Z(n704) );
  XOR2_X1 U751 ( .A(G227), .B(n704), .Z(n700) );
  NAND2_X1 U752 ( .A1(n700), .A2(G900), .ZN(n701) );
  XOR2_X1 U753 ( .A(KEYINPUT124), .B(n701), .Z(n702) );
  NOR2_X1 U754 ( .A1(n707), .A2(n702), .ZN(n703) );
  XNOR2_X1 U755 ( .A(n703), .B(KEYINPUT125), .ZN(n710) );
  XNOR2_X1 U756 ( .A(n704), .B(KEYINPUT123), .ZN(n706) );
  XNOR2_X1 U757 ( .A(n706), .B(n705), .ZN(n708) );
  NAND2_X1 U758 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U759 ( .A1(n710), .A2(n709), .ZN(G72) );
  XOR2_X1 U760 ( .A(G125), .B(KEYINPUT37), .Z(n711) );
  XNOR2_X1 U761 ( .A(n712), .B(n711), .ZN(G27) );
  XOR2_X1 U762 ( .A(G122), .B(n713), .Z(G24) );
  XOR2_X1 U763 ( .A(G140), .B(KEYINPUT112), .Z(n714) );
  XNOR2_X1 U764 ( .A(n715), .B(n714), .ZN(G42) );
  XOR2_X1 U765 ( .A(G137), .B(KEYINPUT126), .Z(n716) );
  XNOR2_X1 U766 ( .A(n717), .B(n716), .ZN(G39) );
  XOR2_X1 U767 ( .A(n718), .B(G131), .Z(G33) );
endmodule

