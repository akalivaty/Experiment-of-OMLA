//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979, new_n980;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT67), .B1(new_n203), .B2(G190gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT28), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207));
  OAI211_X1 g006(.A(KEYINPUT67), .B(KEYINPUT28), .C1(new_n203), .C2(G190gat), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  INV_X1    g008(.A(G176gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT26), .ZN(new_n212));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n214), .B1(new_n212), .B2(new_n213), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n206), .A2(new_n207), .A3(new_n208), .A4(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(KEYINPUT23), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n218), .B1(G169gat), .B2(G176gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n217), .B1(new_n219), .B2(new_n213), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT24), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(KEYINPUT24), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(new_n207), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(KEYINPUT64), .ZN(new_n226));
  AND2_X1   g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n220), .B1(new_n230), .B2(KEYINPUT65), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n224), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT25), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n220), .ZN(new_n235));
  INV_X1    g034(.A(G183gat), .ZN(new_n236));
  INV_X1    g035(.A(G190gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n238), .B(new_n207), .C1(KEYINPUT66), .C2(KEYINPUT24), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT25), .ZN(new_n240));
  NOR2_X1   g039(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n240), .B1(new_n227), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n235), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n216), .B1(new_n234), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G113gat), .A2(G120gat), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(G113gat), .A2(G120gat), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT69), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G113gat), .ZN(new_n250));
  INV_X1    g049(.A(G120gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(new_n253), .A3(new_n246), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT1), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n249), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(G127gat), .A2(G134gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT68), .B(G127gat), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n257), .B1(new_n258), .B2(G134gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  NOR3_X1   g059(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT1), .ZN(new_n261));
  INV_X1    g060(.A(G127gat), .ZN(new_n262));
  INV_X1    g061(.A(G134gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n261), .B1(new_n257), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n245), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n225), .A2(KEYINPUT64), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n226), .B1(new_n227), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n222), .B1(new_n238), .B2(new_n207), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT65), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(new_n233), .A3(new_n235), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n240), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(new_n243), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(new_n266), .A3(new_n216), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n268), .A2(new_n276), .A3(G227gat), .A4(G233gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT32), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n281));
  XNOR2_X1  g080(.A(G15gat), .B(G43gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(G71gat), .B(G99gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT33), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n284), .B1(new_n277), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n280), .A2(new_n281), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n268), .A2(new_n276), .ZN(new_n288));
  NAND2_X1  g087(.A1(G227gat), .A2(G233gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT34), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n277), .B(KEYINPUT32), .C1(new_n285), .C2(new_n284), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n287), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n292), .B1(new_n287), .B2(new_n293), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(G141gat), .A2(G148gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT2), .ZN(new_n301));
  XNOR2_X1  g100(.A(G155gat), .B(G162gat), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n299), .B(new_n301), .C1(new_n302), .C2(KEYINPUT74), .ZN(new_n303));
  OR2_X1    g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(G141gat), .A2(G148gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n301), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(KEYINPUT74), .A3(new_n305), .ZN(new_n307));
  INV_X1    g106(.A(new_n300), .ZN(new_n308));
  NOR2_X1   g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n306), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n260), .A2(new_n303), .A3(new_n311), .A4(new_n265), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n303), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT3), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT3), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n311), .A2(new_n303), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n266), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT4), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n312), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G225gat), .A2(G233gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n324), .A2(KEYINPUT5), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n315), .A2(new_n320), .A3(new_n322), .A4(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n323), .B1(new_n312), .B2(new_n321), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n320), .A2(new_n314), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n327), .B1(new_n328), .B2(new_n312), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n260), .A2(new_n265), .B1(new_n303), .B2(new_n311), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n324), .B1(new_n313), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT5), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n326), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G1gat), .B(G29gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(KEYINPUT0), .ZN(new_n335));
  XNOR2_X1  g134(.A(G57gat), .B(G85gat), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n335), .B(new_n336), .Z(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT6), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n337), .B(new_n326), .C1(new_n329), .C2(new_n332), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n339), .A2(KEYINPUT76), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n333), .A2(KEYINPUT6), .A3(new_n338), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT6), .B1(new_n333), .B2(new_n338), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT76), .B1(new_n345), .B2(new_n341), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G8gat), .B(G36gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(G64gat), .B(G92gat), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n348), .B(new_n349), .Z(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G211gat), .A2(G218gat), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT22), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(G197gat), .A2(G204gat), .ZN(new_n355));
  AND2_X1   g154(.A1(G197gat), .A2(G204gat), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(G211gat), .B(G218gat), .Z(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G211gat), .B(G218gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(G197gat), .B(G204gat), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(new_n361), .A3(new_n354), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(G226gat), .ZN(new_n365));
  INV_X1    g164(.A(G233gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n367), .B1(new_n245), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n367), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n370), .B1(new_n275), .B2(new_n216), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n364), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n245), .A2(new_n367), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT29), .B1(new_n275), .B2(new_n216), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n363), .B(new_n373), .C1(new_n374), .C2(new_n367), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n372), .A2(new_n375), .A3(KEYINPUT72), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT72), .B1(new_n372), .B2(new_n375), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n351), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n372), .A2(new_n375), .A3(new_n350), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT73), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT30), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT30), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n379), .A2(KEYINPUT73), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n378), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n347), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n386));
  AND2_X1   g185(.A1(G228gat), .A2(G233gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n357), .A2(new_n358), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n360), .B1(new_n354), .B2(new_n361), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n368), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n390), .A2(new_n318), .B1(new_n303), .B2(new_n311), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n363), .B1(new_n319), .B2(new_n368), .ZN(new_n392));
  OAI211_X1 g191(.A(KEYINPUT77), .B(new_n387), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n319), .A2(new_n368), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n364), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT29), .B1(new_n359), .B2(new_n362), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n316), .B1(new_n396), .B2(KEYINPUT3), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n387), .A2(KEYINPUT77), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n387), .A2(KEYINPUT77), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n395), .A2(new_n397), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n393), .A2(G22gat), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT78), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT78), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n393), .A2(new_n400), .A3(new_n403), .A4(G22gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n393), .A2(new_n400), .ZN(new_n406));
  INV_X1    g205(.A(G22gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT79), .ZN(new_n409));
  XNOR2_X1  g208(.A(G78gat), .B(G106gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT31), .B(G50gat), .ZN(new_n411));
  XOR2_X1   g210(.A(new_n410), .B(new_n411), .Z(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT79), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n406), .A2(new_n414), .A3(new_n407), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n405), .A2(new_n409), .A3(new_n413), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT80), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n412), .B1(new_n408), .B2(KEYINPUT79), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT80), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n418), .A2(new_n405), .A3(new_n419), .A4(new_n415), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n413), .B1(new_n408), .B2(new_n401), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n386), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  AOI211_X1 g223(.A(KEYINPUT81), .B(new_n422), .C1(new_n417), .C2(new_n420), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n296), .B(new_n385), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n426), .A2(KEYINPUT83), .A3(KEYINPUT35), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT83), .B1(new_n426), .B2(KEYINPUT35), .ZN(new_n428));
  INV_X1    g227(.A(new_n384), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n429), .B(new_n296), .C1(new_n424), .C2(new_n425), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n345), .A2(KEYINPUT82), .A3(new_n341), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n343), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT82), .B1(new_n345), .B2(new_n341), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OR2_X1    g233(.A1(new_n434), .A2(KEYINPUT35), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n427), .A2(new_n428), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n296), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT36), .B1(new_n438), .B2(KEYINPUT71), .ZN(new_n439));
  OAI211_X1 g238(.A(KEYINPUT71), .B(KEYINPUT36), .C1(new_n294), .C2(new_n295), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n424), .ZN(new_n443));
  INV_X1    g242(.A(new_n425), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n315), .A2(new_n320), .A3(new_n322), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n324), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n447), .A2(KEYINPUT39), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT39), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n313), .A2(new_n330), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n449), .B1(new_n450), .B2(new_n323), .ZN(new_n451));
  AOI211_X1 g250(.A(new_n338), .B(new_n448), .C1(new_n447), .C2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n339), .B1(new_n452), .B2(KEYINPUT40), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n453), .B1(KEYINPUT40), .B2(new_n452), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n384), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n376), .A2(new_n377), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT37), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n372), .A2(new_n375), .A3(new_n457), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n459), .A2(KEYINPUT38), .A3(new_n351), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n351), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n372), .A2(new_n375), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n461), .B1(KEYINPUT37), .B2(new_n462), .ZN(new_n463));
  OAI22_X1  g262(.A1(new_n458), .A2(new_n460), .B1(new_n463), .B2(KEYINPUT38), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n464), .A2(new_n379), .A3(new_n434), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n445), .A2(new_n455), .A3(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n443), .B(new_n444), .C1(new_n347), .C2(new_n384), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n442), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT84), .B1(new_n437), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n426), .A2(KEYINPUT35), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n430), .A2(new_n435), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n426), .A2(KEYINPUT83), .A3(KEYINPUT35), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT84), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n442), .A2(new_n466), .A3(new_n467), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n469), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(G113gat), .B(G141gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(G169gat), .B(G197gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n480), .B(new_n481), .ZN(new_n482));
  XOR2_X1   g281(.A(KEYINPUT85), .B(KEYINPUT11), .Z(new_n483));
  XNOR2_X1  g282(.A(new_n482), .B(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(KEYINPUT12), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT92), .ZN(new_n487));
  XNOR2_X1  g286(.A(G15gat), .B(G22gat), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT89), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT90), .ZN(new_n491));
  OAI21_X1  g290(.A(G8gat), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n488), .B(KEYINPUT89), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT16), .ZN(new_n494));
  AOI21_X1  g293(.A(G1gat), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(G8gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(KEYINPUT90), .A3(new_n496), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n492), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n493), .A2(new_n494), .ZN(new_n499));
  INV_X1    g298(.A(G1gat), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n492), .A2(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n487), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT15), .ZN(new_n503));
  XNOR2_X1  g302(.A(KEYINPUT87), .B(G50gat), .ZN(new_n504));
  INV_X1    g303(.A(G43gat), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(G50gat), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n503), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n509));
  NOR3_X1   g308(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n510), .A2(KEYINPUT88), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(KEYINPUT88), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n505), .A2(G50gat), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n514), .A2(new_n507), .A3(new_n503), .ZN(new_n515));
  AND2_X1   g314(.A1(G29gat), .A2(G36gat), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n508), .A2(new_n513), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n509), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(new_n510), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n515), .B1(new_n520), .B2(new_n516), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n499), .A2(new_n500), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n490), .A2(new_n491), .A3(G8gat), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n496), .B1(new_n493), .B2(KEYINPUT90), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n492), .A2(new_n495), .A3(new_n497), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(KEYINPUT92), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n502), .A2(new_n522), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT91), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(new_n498), .B2(new_n501), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n522), .A2(KEYINPUT17), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n533), .A3(new_n521), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n526), .A2(KEYINPUT91), .A3(new_n527), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n531), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G229gat), .A2(G233gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n529), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT18), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(new_n538), .B(KEYINPUT13), .Z(new_n542));
  INV_X1    g341(.A(new_n529), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n522), .B1(new_n502), .B2(new_n528), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n529), .A2(new_n537), .A3(KEYINPUT18), .A4(new_n538), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT93), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n547), .A2(KEYINPUT93), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n546), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT86), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n486), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n547), .B(KEYINPUT93), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n541), .A2(new_n545), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n555), .A2(KEYINPUT86), .A3(new_n485), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n559));
  INV_X1    g358(.A(G155gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G183gat), .B(G211gat), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n561), .B(new_n562), .Z(new_n563));
  NAND2_X1  g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564));
  OR2_X1    g363(.A1(G71gat), .A2(G78gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(G57gat), .B(G64gat), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT9), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n564), .B(new_n565), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT94), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n565), .A2(new_n564), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n571), .B(KEYINPUT94), .C1(new_n567), .C2(new_n566), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT95), .ZN(new_n574));
  INV_X1    g373(.A(G64gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n574), .B1(new_n575), .B2(G57gat), .ZN(new_n576));
  INV_X1    g375(.A(G57gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n577), .A2(KEYINPUT95), .A3(G64gat), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n576), .B(new_n578), .C1(new_n577), .C2(G64gat), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n564), .B1(new_n565), .B2(new_n567), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT96), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(KEYINPUT96), .A3(new_n580), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n573), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT21), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(new_n262), .ZN(new_n589));
  NOR3_X1   g388(.A1(new_n498), .A2(new_n501), .A3(new_n487), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT92), .B1(new_n526), .B2(new_n527), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n584), .A2(new_n585), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n588), .B(G127gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n594), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n563), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n595), .A2(new_n598), .A3(new_n563), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(KEYINPUT97), .B(G85gat), .ZN(new_n603));
  INV_X1    g402(.A(G92gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G85gat), .A2(G92gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT7), .ZN(new_n607));
  INV_X1    g406(.A(G99gat), .ZN(new_n608));
  INV_X1    g407(.A(G106gat), .ZN(new_n609));
  OAI21_X1  g408(.A(KEYINPUT8), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n605), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G99gat), .B(G106gat), .Z(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n612), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n614), .A2(new_n605), .A3(new_n607), .A4(new_n610), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n535), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n616), .ZN(new_n618));
  AND2_X1   g417(.A1(G232gat), .A2(G233gat), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n522), .A2(new_n618), .B1(KEYINPUT41), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G190gat), .B(G218gat), .Z(new_n622));
  AND2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n619), .A2(KEYINPUT41), .ZN(new_n625));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  OR3_X1    g427(.A1(new_n623), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n628), .B1(new_n623), .B2(new_n624), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT98), .B1(new_n602), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n601), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n631), .B(KEYINPUT98), .C1(new_n633), .C2(new_n599), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G230gat), .A2(G233gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n584), .A2(new_n616), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n579), .A2(KEYINPUT96), .A3(new_n580), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n640), .A2(new_n581), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n641), .A2(new_n573), .A3(new_n615), .A4(new_n613), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n638), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G120gat), .B(G148gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(G176gat), .B(G204gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n644), .B(new_n645), .Z(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n638), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT10), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n639), .A2(new_n649), .A3(new_n642), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT99), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n639), .A2(KEYINPUT99), .A3(new_n642), .A4(new_n649), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n642), .A2(new_n649), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n648), .B1(new_n655), .B2(KEYINPUT100), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n652), .A2(new_n657), .A3(new_n653), .A4(new_n654), .ZN(new_n658));
  AOI211_X1 g457(.A(new_n643), .B(new_n647), .C1(new_n656), .C2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n646), .B(KEYINPUT101), .Z(new_n661));
  AND2_X1   g460(.A1(new_n655), .A2(new_n638), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n661), .B1(new_n662), .B2(new_n643), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n637), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n479), .A2(new_n558), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n557), .B1(new_n469), .B2(new_n478), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n669), .A2(KEYINPUT102), .A3(new_n665), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n347), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g472(.A(KEYINPUT16), .B(G8gat), .Z(new_n674));
  AND3_X1   g473(.A1(new_n671), .A2(new_n384), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT103), .B1(new_n675), .B2(KEYINPUT42), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n496), .B1(new_n671), .B2(new_n384), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n677), .B1(new_n675), .B2(KEYINPUT42), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n671), .A2(new_n384), .A3(new_n674), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n676), .A2(new_n678), .A3(new_n682), .ZN(G1325gat));
  INV_X1    g482(.A(G15gat), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n671), .A2(new_n684), .A3(new_n296), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n442), .B1(new_n668), .B2(new_n670), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n685), .B1(new_n686), .B2(new_n684), .ZN(G1326gat));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n688));
  INV_X1    g487(.A(new_n445), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n671), .B2(new_n689), .ZN(new_n690));
  AOI211_X1 g489(.A(KEYINPUT104), .B(new_n445), .C1(new_n668), .C2(new_n670), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT43), .B(G22gat), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n690), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n670), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT102), .B1(new_n669), .B2(new_n665), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n689), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT104), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n671), .A2(new_n688), .A3(new_n689), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n692), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n694), .A2(new_n700), .ZN(G1327gat));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702));
  INV_X1    g501(.A(new_n631), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n702), .B1(new_n479), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n475), .A2(new_n477), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(KEYINPUT106), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n707), .B1(new_n475), .B2(new_n477), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n703), .A2(new_n702), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n706), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n704), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n602), .B(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(new_n557), .A3(new_n664), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n347), .ZN(new_n717));
  OAI21_X1  g516(.A(G29gat), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n602), .A2(new_n664), .A3(new_n631), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n669), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n717), .A2(G29gat), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n719), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n669), .A2(KEYINPUT45), .A3(new_n720), .A4(new_n722), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n718), .A2(new_n724), .A3(new_n725), .ZN(G1328gat));
  OAI21_X1  g525(.A(G36gat), .B1(new_n716), .B2(new_n429), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n429), .A2(G36gat), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT46), .B1(new_n721), .B2(new_n729), .ZN(new_n730));
  OR3_X1    g529(.A1(new_n721), .A2(KEYINPUT46), .A3(new_n729), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n727), .A2(new_n730), .A3(new_n731), .ZN(G1329gat));
  NAND2_X1  g531(.A1(new_n296), .A2(new_n505), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n721), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n442), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n735), .B(new_n715), .C1(new_n704), .C2(new_n710), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n734), .B1(new_n736), .B2(G43gat), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT47), .ZN(G1330gat));
  OR2_X1    g537(.A1(new_n445), .A2(new_n504), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n721), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n689), .B(new_n715), .C1(new_n704), .C2(new_n710), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(new_n504), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g542(.A1(new_n706), .A2(new_n708), .ZN(new_n744));
  INV_X1    g543(.A(new_n664), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n637), .A2(new_n558), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(new_n717), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(new_n577), .ZN(G1332gat));
  NOR2_X1   g548(.A1(new_n747), .A2(new_n429), .ZN(new_n750));
  NOR2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  AND2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n750), .B2(new_n751), .ZN(G1333gat));
  OAI21_X1  g553(.A(G71gat), .B1(new_n747), .B2(new_n442), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n438), .A2(G71gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n747), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g557(.A1(new_n747), .A2(new_n445), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n759), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g559(.A1(new_n558), .A2(new_n602), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n703), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n762), .B1(new_n475), .B2(new_n477), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n763), .A2(KEYINPUT51), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(KEYINPUT51), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT107), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n767), .A2(new_n347), .A3(new_n603), .A4(new_n664), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n761), .A2(new_n664), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n711), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n717), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n768), .B1(new_n772), .B2(new_n603), .ZN(G1336gat));
  OAI211_X1 g572(.A(new_n384), .B(new_n770), .C1(new_n704), .C2(new_n710), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G92gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n766), .A2(new_n664), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n384), .A2(new_n604), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT52), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n775), .B(new_n780), .C1(new_n776), .C2(new_n777), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(G1337gat));
  OAI21_X1  g581(.A(G99gat), .B1(new_n771), .B2(new_n442), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n767), .A2(new_n608), .A3(new_n296), .A4(new_n664), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1338gat));
  INV_X1    g584(.A(KEYINPUT108), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n689), .B(new_n770), .C1(new_n704), .C2(new_n710), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n786), .B1(new_n787), .B2(G106gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n689), .A2(new_n609), .ZN(new_n789));
  AOI211_X1 g588(.A(new_n745), .B(new_n789), .C1(new_n764), .C2(new_n765), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n787), .B2(G106gat), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n788), .A2(new_n791), .A3(KEYINPUT53), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793));
  AOI221_X4 g592(.A(new_n790), .B1(new_n786), .B2(new_n793), .C1(new_n787), .C2(G106gat), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n792), .A2(new_n794), .ZN(G1339gat));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n655), .A2(new_n796), .A3(new_n638), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n647), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n656), .A2(new_n658), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT54), .B1(new_n655), .B2(new_n638), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n798), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n659), .B1(new_n802), .B2(KEYINPUT55), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n800), .B1(new_n658), .B2(new_n656), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(new_n798), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n552), .A2(new_n556), .A3(new_n803), .A4(new_n806), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n543), .A2(new_n544), .A3(new_n542), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n538), .B1(new_n529), .B2(new_n537), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n484), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n553), .A2(new_n554), .A3(new_n485), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n664), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n703), .B1(new_n807), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n811), .A2(new_n810), .ZN(new_n814));
  AND4_X1   g613(.A1(new_n703), .A2(new_n814), .A3(new_n806), .A4(new_n803), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n713), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n636), .A2(new_n557), .A3(new_n745), .ZN(new_n817));
  AOI211_X1 g616(.A(new_n717), .B(new_n430), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(G113gat), .B1(new_n818), .B2(new_n558), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n689), .B1(new_n816), .B2(new_n817), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n717), .A2(new_n384), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(new_n438), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n557), .A2(new_n250), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n819), .B1(new_n823), .B2(new_n824), .ZN(G1340gat));
  AOI21_X1  g624(.A(G120gat), .B1(new_n818), .B2(new_n664), .ZN(new_n826));
  INV_X1    g625(.A(new_n822), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n745), .A2(new_n438), .A3(new_n251), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(G1341gat));
  NAND2_X1  g628(.A1(new_n823), .A2(new_n714), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n258), .ZN(new_n831));
  INV_X1    g630(.A(new_n602), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(new_n258), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT109), .ZN(G1342gat));
  NAND3_X1  g635(.A1(new_n818), .A2(new_n263), .A3(new_n703), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT56), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n263), .B1(new_n823), .B2(new_n703), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT110), .ZN(G1343gat));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n816), .A2(new_n817), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n442), .A2(new_n689), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n384), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n843), .A2(new_n347), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(G141gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n847), .A3(new_n558), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT113), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n842), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n850), .B1(new_n848), .B2(new_n849), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT112), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n802), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT112), .B1(new_n805), .B2(new_n798), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(new_n855), .A3(new_n804), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n856), .A2(new_n552), .A3(new_n556), .A4(new_n803), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n703), .B1(new_n857), .B2(new_n812), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n832), .B1(new_n858), .B2(new_n815), .ZN(new_n859));
  AOI211_X1 g658(.A(new_n852), .B(new_n445), .C1(new_n859), .C2(new_n817), .ZN(new_n860));
  XNOR2_X1  g659(.A(KEYINPUT111), .B(KEYINPUT57), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n862), .B1(new_n843), .B2(new_n689), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n442), .A2(new_n821), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n558), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(G141gat), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n851), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n851), .B2(new_n868), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n868), .A2(new_n848), .ZN(new_n872));
  OAI22_X1  g671(.A1(new_n870), .A2(new_n871), .B1(new_n872), .B2(new_n842), .ZN(G1344gat));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n874));
  INV_X1    g673(.A(G148gat), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n843), .A2(new_n689), .A3(new_n862), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n445), .B1(new_n859), .B2(new_n817), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(KEYINPUT57), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT116), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n664), .B1(new_n865), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n880), .B1(new_n879), .B2(new_n865), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n875), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n874), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n859), .A2(new_n817), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT57), .B1(new_n885), .B2(new_n689), .ZN(new_n886));
  AOI211_X1 g685(.A(new_n445), .B(new_n861), .C1(new_n816), .C2(new_n817), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n881), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(G148gat), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(KEYINPUT117), .A3(KEYINPUT59), .ZN(new_n890));
  INV_X1    g689(.A(new_n865), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n664), .B(new_n891), .C1(new_n860), .C2(new_n863), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n875), .A2(KEYINPUT59), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT115), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n892), .A2(KEYINPUT115), .A3(new_n893), .ZN(new_n897));
  AOI22_X1  g696(.A1(new_n884), .A2(new_n890), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n846), .A2(new_n875), .A3(new_n664), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT118), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT117), .B1(new_n889), .B2(KEYINPUT59), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n882), .A2(new_n874), .A3(new_n883), .ZN(new_n903));
  INV_X1    g702(.A(new_n897), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT115), .B1(new_n892), .B2(new_n893), .ZN(new_n905));
  OAI22_X1  g704(.A1(new_n902), .A2(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n907), .A3(new_n899), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n901), .A2(new_n908), .ZN(G1345gat));
  AOI21_X1  g708(.A(KEYINPUT119), .B1(new_n846), .B2(new_n602), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(G155gat), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n846), .A2(KEYINPUT119), .A3(new_n602), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n713), .A2(new_n560), .ZN(new_n913));
  AOI22_X1  g712(.A1(new_n911), .A2(new_n912), .B1(new_n866), .B2(new_n913), .ZN(G1346gat));
  AOI21_X1  g713(.A(G162gat), .B1(new_n846), .B2(new_n703), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n703), .A2(G162gat), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n866), .B2(new_n916), .ZN(G1347gat));
  AOI21_X1  g716(.A(new_n347), .B1(new_n816), .B2(new_n817), .ZN(new_n918));
  AND4_X1   g717(.A1(new_n445), .A2(new_n918), .A3(new_n384), .A4(new_n296), .ZN(new_n919));
  AOI21_X1  g718(.A(G169gat), .B1(new_n919), .B2(new_n558), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n429), .A2(new_n347), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n820), .A2(new_n296), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n557), .A2(new_n209), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(G1348gat));
  AOI21_X1  g723(.A(G176gat), .B1(new_n919), .B2(new_n664), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT120), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n745), .A2(new_n210), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n926), .B1(new_n922), .B2(new_n927), .ZN(G1349gat));
  NAND2_X1  g727(.A1(new_n922), .A2(new_n714), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n236), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n931), .B1(new_n930), .B2(new_n929), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n919), .A2(new_n202), .A3(new_n602), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g734(.A(new_n237), .B1(new_n922), .B2(new_n703), .ZN(new_n936));
  XOR2_X1   g735(.A(new_n936), .B(KEYINPUT61), .Z(new_n937));
  NAND3_X1  g736(.A1(new_n919), .A2(new_n237), .A3(new_n703), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1351gat));
  NOR2_X1   g738(.A1(new_n844), .A2(new_n429), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n918), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(G197gat), .B1(new_n942), .B2(new_n558), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n878), .B(KEYINPUT122), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n442), .A2(new_n921), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n946), .A2(G197gat), .A3(new_n558), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n943), .B1(new_n944), .B2(new_n947), .ZN(G1352gat));
  INV_X1    g747(.A(KEYINPUT124), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n745), .A2(G204gat), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(KEYINPUT123), .B1(new_n941), .B2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n941), .A2(KEYINPUT123), .A3(new_n951), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(new_n954), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT62), .B1(new_n957), .B2(new_n952), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(G204gat), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n945), .A2(new_n745), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n960), .B1(new_n944), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n949), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n956), .A2(new_n958), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n944), .A2(new_n961), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n964), .B(KEYINPUT124), .C1(new_n965), .C2(new_n960), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n963), .A2(new_n966), .ZN(G1353gat));
  NAND3_X1  g766(.A1(new_n878), .A2(new_n602), .A3(new_n946), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n968), .B(G211gat), .C1(new_n969), .C2(KEYINPUT63), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n969), .A2(KEYINPUT63), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OR3_X1    g771(.A1(new_n941), .A2(G211gat), .A3(new_n832), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n970), .A2(new_n971), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(G1354gat));
  AOI21_X1  g774(.A(G218gat), .B1(new_n942), .B2(new_n703), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n703), .A2(G218gat), .ZN(new_n977));
  XOR2_X1   g776(.A(new_n977), .B(KEYINPUT126), .Z(new_n978));
  NOR2_X1   g777(.A1(new_n945), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n976), .B1(new_n944), .B2(new_n979), .ZN(new_n980));
  XOR2_X1   g779(.A(new_n980), .B(KEYINPUT127), .Z(G1355gat));
endmodule


