//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997;
  XOR2_X1   g000(.A(KEYINPUT73), .B(KEYINPUT0), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT74), .ZN(new_n203));
  XNOR2_X1  g002(.A(G1gat), .B(G29gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G57gat), .B(G85gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(G141gat), .B(G148gat), .Z(new_n208));
  INV_X1    g007(.A(G155gat), .ZN(new_n209));
  INV_X1    g008(.A(G162gat), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT2), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G155gat), .B(G162gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(G113gat), .B(G120gat), .Z(new_n216));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G127gat), .B(G134gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n208), .A2(new_n213), .A3(new_n211), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n216), .A2(new_n217), .A3(new_n219), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n215), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(KEYINPUT4), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n215), .A2(new_n222), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT3), .ZN(new_n227));
  XOR2_X1   g026(.A(KEYINPUT71), .B(KEYINPUT3), .Z(new_n228));
  NAND3_X1  g027(.A1(new_n215), .A2(new_n222), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n221), .A2(new_n223), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n225), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G225gat), .A2(G233gat), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n207), .B1(new_n235), .B2(KEYINPUT39), .ZN(new_n236));
  INV_X1    g035(.A(new_n224), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n215), .A2(new_n222), .B1(new_n221), .B2(new_n223), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT39), .B1(new_n239), .B2(new_n234), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n240), .B1(new_n234), .B2(new_n232), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT78), .B1(new_n236), .B2(new_n241), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n242), .A2(KEYINPUT40), .ZN(new_n243));
  INV_X1    g042(.A(new_n207), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n234), .B1(new_n237), .B2(new_n238), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT5), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n233), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT4), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n237), .A2(KEYINPUT72), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT72), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n251), .B1(new_n224), .B2(KEYINPUT4), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n224), .A2(KEYINPUT4), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n246), .B1(new_n248), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT5), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n224), .A2(KEYINPUT4), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n224), .A2(KEYINPUT4), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n259), .A2(new_n247), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n244), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n242), .A2(KEYINPUT40), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n243), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G169gat), .ZN(new_n264));
  INV_X1    g063(.A(G176gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(G169gat), .A2(G176gat), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n266), .B1(KEYINPUT23), .B2(new_n267), .ZN(new_n268));
  OR3_X1    g067(.A1(new_n267), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT64), .B1(new_n267), .B2(KEYINPUT23), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n268), .A2(KEYINPUT25), .A3(new_n269), .A4(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT24), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n273), .A2(KEYINPUT65), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(KEYINPUT65), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n272), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT66), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(G183gat), .B2(G190gat), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n280), .B1(new_n276), .B2(new_n277), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n271), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n272), .A2(new_n273), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n283), .B(new_n279), .C1(G183gat), .C2(G190gat), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n268), .A2(new_n284), .A3(new_n269), .A4(new_n270), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT25), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT27), .B(G183gat), .ZN(new_n289));
  INV_X1    g088(.A(G190gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT28), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n267), .A2(KEYINPUT26), .ZN(new_n293));
  INV_X1    g092(.A(new_n267), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT26), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n272), .B(new_n293), .C1(new_n296), .C2(new_n266), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G226gat), .A2(G233gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  OAI22_X1  g099(.A1(new_n288), .A2(new_n298), .B1(KEYINPUT29), .B2(new_n300), .ZN(new_n301));
  OR2_X1    g100(.A1(new_n292), .A2(new_n297), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n302), .B(new_n299), .C1(new_n287), .C2(new_n282), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT68), .B(G211gat), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT22), .B1(new_n304), .B2(G218gat), .ZN(new_n305));
  XOR2_X1   g104(.A(G197gat), .B(G204gat), .Z(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G211gat), .B(G218gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT69), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n307), .B(new_n310), .ZN(new_n311));
  AND3_X1   g110(.A1(new_n301), .A2(new_n303), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(KEYINPUT70), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n305), .A2(new_n306), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(new_n310), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n307), .B1(new_n309), .B2(new_n308), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT70), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n301), .A2(new_n303), .B1(new_n313), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G8gat), .B(G36gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(G64gat), .B(G92gat), .ZN(new_n322));
  XOR2_X1   g121(.A(new_n321), .B(new_n322), .Z(new_n323));
  OR3_X1    g122(.A1(new_n312), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n323), .B1(new_n312), .B2(new_n320), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(KEYINPUT30), .A3(new_n325), .ZN(new_n326));
  OR2_X1    g125(.A1(new_n312), .A2(new_n320), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT30), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(new_n328), .A3(new_n323), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n263), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT38), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT37), .ZN(new_n333));
  OR2_X1    g132(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT79), .B(KEYINPUT37), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(new_n312), .B2(new_n320), .ZN(new_n336));
  INV_X1    g135(.A(new_n323), .ZN(new_n337));
  AND2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n332), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT6), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n248), .A2(new_n256), .A3(new_n225), .ZN(new_n341));
  NOR3_X1   g140(.A1(new_n224), .A2(new_n251), .A3(KEYINPUT4), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n342), .A2(new_n257), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n247), .B1(new_n343), .B2(new_n252), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n341), .B(new_n207), .C1(new_n344), .C2(new_n246), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n261), .A2(new_n340), .A3(new_n345), .ZN(new_n346));
  OAI211_X1 g145(.A(KEYINPUT6), .B(new_n244), .C1(new_n255), .C2(new_n260), .ZN(new_n347));
  AND2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n301), .A2(new_n303), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n333), .B1(new_n349), .B2(new_n317), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n301), .A2(new_n303), .A3(new_n313), .A4(new_n319), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT38), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n352), .A2(KEYINPUT80), .A3(new_n337), .A4(new_n336), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n300), .A2(KEYINPUT29), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n282), .A2(new_n287), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n354), .B1(new_n355), .B2(new_n302), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n288), .A2(new_n298), .A3(new_n300), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n317), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n358), .A2(KEYINPUT37), .A3(new_n351), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n336), .A2(new_n359), .A3(new_n332), .A4(new_n337), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT80), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n348), .A2(new_n325), .A3(new_n353), .A4(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT81), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n339), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n346), .A2(new_n347), .A3(new_n325), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n366), .A2(KEYINPUT81), .A3(new_n353), .A4(new_n362), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n331), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n230), .B1(new_n288), .B2(new_n298), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n221), .A2(new_n223), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n302), .B(new_n370), .C1(new_n287), .C2(new_n282), .ZN(new_n371));
  INV_X1    g170(.A(G227gat), .ZN(new_n372));
  INV_X1    g171(.A(G233gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n369), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT34), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(G15gat), .B(G43gat), .Z(new_n379));
  XNOR2_X1  g178(.A(G71gat), .B(G99gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n375), .B1(new_n369), .B2(new_n371), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n381), .B1(new_n382), .B2(KEYINPUT33), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT32), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n387));
  AOI221_X4 g186(.A(new_n384), .B1(KEYINPUT33), .B2(new_n381), .C1(new_n387), .C2(new_n374), .ZN(new_n388));
  OAI211_X1 g187(.A(KEYINPUT67), .B(new_n378), .C1(new_n386), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n374), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT32), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT33), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(new_n393), .A3(new_n381), .ZN(new_n394));
  INV_X1    g193(.A(new_n388), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n376), .B(KEYINPUT34), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n378), .A2(KEYINPUT67), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n389), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT36), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n378), .B1(new_n386), .B2(new_n388), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT36), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n397), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT76), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT29), .ZN(new_n406));
  INV_X1    g205(.A(new_n308), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n406), .B1(new_n307), .B2(new_n407), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n305), .A2(new_n308), .A3(new_n306), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n228), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n229), .A2(new_n406), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n410), .A2(new_n226), .B1(new_n311), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G228gat), .A2(G233gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT77), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT77), .ZN(new_n416));
  INV_X1    g215(.A(new_n226), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n314), .A2(new_n308), .ZN(new_n418));
  INV_X1    g217(.A(new_n409), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n418), .A2(new_n406), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n417), .B1(new_n420), .B2(new_n228), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n411), .A2(new_n316), .A3(new_n315), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n416), .B(new_n413), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n415), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(G22gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n311), .A2(KEYINPUT29), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n226), .B1(new_n426), .B2(KEYINPUT3), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n313), .A2(new_n319), .A3(new_n411), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n428), .A3(new_n414), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n424), .A2(new_n425), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n425), .B1(new_n424), .B2(new_n429), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n405), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G78gat), .B(G106gat), .ZN(new_n433));
  INV_X1    g232(.A(G50gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n424), .A2(new_n429), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(G22gat), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n424), .A2(new_n425), .A3(new_n429), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n435), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n405), .A3(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT75), .B(KEYINPUT31), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n436), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n443), .B1(new_n436), .B2(new_n442), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n404), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n326), .A2(new_n329), .B1(new_n346), .B2(new_n347), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n397), .A2(new_n401), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n443), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n441), .B1(new_n440), .B2(new_n405), .ZN(new_n451));
  AOI211_X1 g250(.A(KEYINPUT76), .B(new_n435), .C1(new_n438), .C2(new_n439), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n442), .A3(new_n443), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n449), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI22_X1  g254(.A1(new_n368), .A2(new_n446), .B1(KEYINPUT35), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n447), .ZN(new_n457));
  OAI211_X1 g256(.A(KEYINPUT35), .B(new_n399), .C1(new_n444), .C2(new_n445), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n404), .A2(new_n454), .A3(new_n453), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT87), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n425), .A2(G15gat), .ZN(new_n463));
  INV_X1    g262(.A(G15gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G22gat), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT16), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(G1gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(G15gat), .B(G22gat), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n467), .A2(new_n468), .B1(new_n469), .B2(KEYINPUT84), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n469), .A2(KEYINPUT84), .A3(KEYINPUT16), .A4(new_n468), .ZN(new_n472));
  XOR2_X1   g271(.A(KEYINPUT85), .B(G8gat), .Z(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n472), .ZN(new_n475));
  INV_X1    g274(.A(G8gat), .ZN(new_n476));
  OAI22_X1  g275(.A1(new_n475), .A2(new_n470), .B1(KEYINPUT85), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT83), .B1(G29gat), .B2(G36gat), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT14), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n481), .A2(new_n482), .B1(G29gat), .B2(G36gat), .ZN(new_n483));
  OR3_X1    g282(.A1(KEYINPUT83), .A2(G29gat), .A3(G36gat), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(KEYINPUT14), .A3(new_n480), .ZN(new_n485));
  INV_X1    g284(.A(G43gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n434), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT15), .ZN(new_n488));
  NAND2_X1  g287(.A1(G43gat), .A2(G50gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n483), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G43gat), .B(G50gat), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n488), .B1(new_n492), .B2(KEYINPUT82), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT82), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n487), .A2(new_n494), .A3(new_n489), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n493), .A2(new_n483), .A3(new_n495), .A4(new_n485), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(KEYINPUT17), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT17), .B1(new_n497), .B2(new_n498), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n479), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G229gat), .A2(G233gat), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n497), .A2(new_n498), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n478), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n507));
  AOI21_X1  g306(.A(new_n462), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G113gat), .B(G141gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(G197gat), .ZN(new_n510));
  XOR2_X1   g309(.A(KEYINPUT11), .B(G169gat), .Z(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT12), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n498), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n515), .A2(new_n474), .A3(new_n477), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n505), .A2(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(new_n503), .B(KEYINPUT13), .Z(new_n518));
  AOI22_X1  g317(.A1(new_n506), .A2(new_n507), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n502), .A2(KEYINPUT18), .A3(new_n503), .A4(new_n505), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n519), .B(new_n520), .C1(new_n508), .C2(new_n513), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n461), .A2(new_n525), .ZN(new_n526));
  XOR2_X1   g325(.A(G127gat), .B(G155gat), .Z(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(KEYINPUT20), .ZN(new_n528));
  NAND2_X1  g327(.A1(G231gat), .A2(G233gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT91), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n528), .B(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G183gat), .B(G211gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT89), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n535), .A2(KEYINPUT88), .A3(G57gat), .ZN(new_n536));
  OR2_X1    g335(.A1(KEYINPUT88), .A2(G57gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(G64gat), .ZN(new_n539));
  INV_X1    g338(.A(G71gat), .ZN(new_n540));
  INV_X1    g339(.A(G78gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n541), .A3(KEYINPUT9), .ZN(new_n542));
  NAND2_X1  g341(.A1(G71gat), .A2(G78gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n535), .A2(G57gat), .ZN(new_n544));
  INV_X1    g343(.A(G64gat), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n542), .A2(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G57gat), .A2(G64gat), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n540), .A2(new_n541), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n551), .A2(new_n543), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n539), .A2(new_n546), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT93), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n543), .B(new_n551), .C1(new_n548), .C2(new_n549), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n542), .A2(new_n543), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n544), .A2(new_n545), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n545), .B1(new_n536), .B2(new_n537), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n555), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT93), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n554), .A2(new_n562), .A3(KEYINPUT21), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n479), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT94), .ZN(new_n565));
  XOR2_X1   g364(.A(KEYINPUT90), .B(KEYINPUT21), .Z(new_n566));
  NAND2_X1  g365(.A1(new_n560), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n565), .A2(new_n569), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n534), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n572), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(new_n570), .A3(new_n533), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n578), .A2(KEYINPUT41), .ZN(new_n579));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(KEYINPUT96), .A2(G85gat), .A3(G92gat), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT95), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(KEYINPUT95), .A2(G85gat), .A3(G92gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n585), .A2(KEYINPUT7), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G99gat), .B(G106gat), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT7), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n583), .A2(new_n584), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G99gat), .A2(G106gat), .ZN(new_n591));
  INV_X1    g390(.A(G85gat), .ZN(new_n592));
  INV_X1    g391(.A(G92gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(KEYINPUT8), .A2(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n587), .A2(new_n588), .A3(new_n590), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT97), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n594), .A2(new_n590), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT97), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n597), .A2(new_n598), .A3(new_n588), .A4(new_n587), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT98), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n583), .A2(new_n584), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n586), .A2(KEYINPUT7), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n590), .B(new_n594), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n588), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n601), .A3(new_n605), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n600), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n609), .B1(new_n500), .B2(new_n501), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n604), .A2(new_n605), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT98), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n612), .A2(new_n607), .B1(new_n596), .B2(new_n599), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n504), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n578), .A2(KEYINPUT41), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n610), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G190gat), .B(G218gat), .Z(new_n617));
  AND2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n582), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n616), .A2(new_n617), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n616), .A2(new_n617), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n621), .A2(new_n622), .A3(new_n581), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n577), .A2(KEYINPUT99), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT99), .ZN(new_n626));
  INV_X1    g425(.A(new_n624), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n576), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G230gat), .A2(G233gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n609), .A2(new_n560), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n611), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n603), .B1(new_n584), .B2(new_n583), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n594), .A2(new_n590), .ZN(new_n635));
  OAI211_X1 g434(.A(KEYINPUT100), .B(new_n605), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n600), .A2(new_n553), .A3(new_n633), .A4(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n630), .B1(new_n631), .B2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT101), .B(KEYINPUT10), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n637), .B(new_n639), .C1(new_n613), .C2(new_n553), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n554), .A2(new_n562), .A3(KEYINPUT10), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n613), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n638), .B1(new_n644), .B2(new_n630), .ZN(new_n645));
  XNOR2_X1  g444(.A(G120gat), .B(G148gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(G176gat), .B(G204gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n646), .B(new_n647), .Z(new_n648));
  NOR2_X1   g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n638), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n609), .A2(new_n641), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n553), .ZN(new_n652));
  AOI21_X1  g451(.A(KEYINPUT100), .B1(new_n604), .B2(new_n605), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n609), .A2(new_n560), .B1(new_n654), .B2(new_n600), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n651), .B1(new_n655), .B2(new_n639), .ZN(new_n656));
  INV_X1    g455(.A(new_n630), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n650), .B(new_n648), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n645), .A2(KEYINPUT102), .A3(new_n648), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n649), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n629), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n526), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n348), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(new_n468), .ZN(G1324gat));
  INV_X1    g466(.A(new_n330), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT103), .B(KEYINPUT16), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(new_n476), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n526), .A2(new_n668), .A3(new_n663), .A4(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(G8gat), .B1(new_n664), .B2(new_n330), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n671), .ZN(new_n673));
  MUX2_X1   g472(.A(new_n671), .B(new_n673), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g473(.A(G15gat), .B1(new_n664), .B2(new_n404), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n448), .A2(new_n464), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n675), .B1(new_n664), .B2(new_n676), .ZN(G1326gat));
  NOR2_X1   g476(.A1(new_n444), .A2(new_n445), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n526), .A2(new_n678), .A3(new_n663), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  NAND2_X1  g480(.A1(new_n363), .A2(new_n364), .ZN(new_n682));
  INV_X1    g481(.A(new_n339), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n682), .A2(new_n367), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n331), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n453), .A2(new_n454), .B1(new_n400), .B2(new_n403), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n447), .B(new_n448), .C1(new_n444), .C2(new_n445), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT35), .ZN(new_n689));
  AOI22_X1  g488(.A1(new_n686), .A2(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n458), .A2(new_n459), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n447), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n576), .A2(new_n662), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n694), .A2(new_n525), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(new_n627), .A3(new_n695), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n696), .A2(G29gat), .A3(new_n665), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n627), .B1(new_n456), .B2(new_n460), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI211_X1 g501(.A(KEYINPUT44), .B(new_n627), .C1(new_n456), .C2(new_n460), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(new_n695), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(G29gat), .B1(new_n704), .B2(new_n665), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n699), .A2(new_n705), .ZN(G1328gat));
  OR2_X1    g505(.A1(new_n330), .A2(G36gat), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT46), .B1(new_n696), .B2(new_n707), .ZN(new_n708));
  OR3_X1    g507(.A1(new_n696), .A2(KEYINPUT46), .A3(new_n707), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n702), .A2(new_n668), .A3(new_n695), .A4(new_n703), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G36gat), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n710), .A2(new_n711), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n708), .B(new_n709), .C1(new_n713), .C2(new_n714), .ZN(G1329gat));
  INV_X1    g514(.A(new_n448), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n486), .B1(new_n696), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n404), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G43gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n717), .B1(new_n704), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g520(.A1(new_n702), .A2(new_n678), .A3(new_n695), .A4(new_n703), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(G50gat), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n694), .A2(G50gat), .A3(new_n624), .ZN(new_n724));
  AND4_X1   g523(.A1(new_n524), .A2(new_n693), .A3(new_n678), .A4(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT48), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n725), .B1(new_n722), .B2(G50gat), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n730), .A2(KEYINPUT106), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n729), .A2(new_n732), .ZN(G1331gat));
  AOI21_X1  g532(.A(KEYINPUT102), .B1(new_n645), .B2(new_n648), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n657), .B1(new_n640), .B2(new_n643), .ZN(new_n735));
  INV_X1    g534(.A(new_n648), .ZN(new_n736));
  NOR4_X1   g535(.A1(new_n735), .A2(new_n638), .A3(new_n659), .A4(new_n736), .ZN(new_n737));
  OAI22_X1  g536(.A1(new_n734), .A2(new_n737), .B1(new_n645), .B2(new_n648), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n629), .A2(new_n525), .A3(new_n738), .ZN(new_n739));
  OR2_X1    g538(.A1(new_n461), .A2(new_n739), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n740), .A2(new_n665), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT88), .B(G57gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1332gat));
  NOR2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  OR3_X1    g546(.A1(new_n461), .A2(new_n746), .A3(new_n739), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n330), .B(KEYINPUT108), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n751), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n745), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n752), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n749), .A2(new_n744), .A3(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n753), .A2(new_n755), .ZN(G1333gat));
  NAND4_X1  g555(.A1(new_n747), .A2(G71gat), .A3(new_n718), .A4(new_n748), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n540), .B1(new_n740), .B2(new_n716), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n757), .A2(KEYINPUT50), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT50), .B1(new_n757), .B2(new_n758), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(G1334gat));
  XNOR2_X1  g560(.A(KEYINPUT109), .B(G78gat), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n750), .A2(new_n678), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n762), .ZN(new_n764));
  INV_X1    g563(.A(new_n678), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n749), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n766), .ZN(G1335gat));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT51), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n577), .A2(new_n524), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n768), .B2(KEYINPUT51), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n770), .B1(new_n700), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n772), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n693), .A2(new_n627), .A3(new_n774), .A4(new_n769), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n773), .A2(new_n738), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n776), .A2(new_n592), .A3(new_n348), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n577), .A2(new_n524), .A3(new_n662), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n702), .A2(new_n348), .A3(new_n703), .A4(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G85gat), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n779), .A2(new_n780), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n777), .B1(new_n782), .B2(new_n783), .ZN(G1336gat));
  NOR2_X1   g583(.A1(new_n751), .A2(G92gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n776), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n702), .A2(new_n703), .A3(new_n778), .ZN(new_n788));
  OAI21_X1  g587(.A(G92gat), .B1(new_n788), .B2(new_n751), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n702), .A2(new_n668), .A3(new_n703), .A4(new_n778), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n776), .A2(new_n785), .B1(G92gat), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n790), .B1(new_n792), .B2(new_n787), .ZN(G1337gat));
  NAND2_X1  g592(.A1(new_n718), .A2(G99gat), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n788), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n773), .A2(new_n775), .A3(new_n448), .A4(new_n738), .ZN(new_n796));
  INV_X1    g595(.A(G99gat), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT112), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT112), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n795), .A2(new_n798), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(G1338gat));
  NAND4_X1  g602(.A1(new_n702), .A2(new_n678), .A3(new_n703), .A4(new_n778), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n804), .A2(G106gat), .B1(KEYINPUT113), .B2(KEYINPUT53), .ZN(new_n805));
  OR2_X1    g604(.A1(KEYINPUT113), .A2(KEYINPUT53), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n765), .A2(G106gat), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n773), .A2(new_n775), .A3(new_n738), .A4(new_n807), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n805), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n806), .B1(new_n805), .B2(new_n808), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(G1339gat));
  NAND2_X1  g610(.A1(new_n660), .A2(new_n661), .ZN(new_n812));
  INV_X1    g611(.A(new_n735), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n630), .B1(new_n642), .B2(new_n613), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n640), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n640), .A2(new_n814), .A3(KEYINPUT114), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n813), .A2(new_n817), .A3(KEYINPUT54), .A4(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n648), .B1(new_n735), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n819), .A2(KEYINPUT55), .A3(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n812), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n644), .A2(new_n820), .A3(new_n630), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n736), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n735), .A2(new_n820), .ZN(new_n827));
  INV_X1    g626(.A(new_n818), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT114), .B1(new_n640), .B2(new_n814), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n826), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n824), .B1(new_n831), .B2(KEYINPUT55), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n819), .A2(new_n821), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n833), .A2(KEYINPUT115), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n503), .B1(new_n502), .B2(new_n505), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n517), .A2(new_n518), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n512), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT116), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n506), .A2(new_n507), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n517), .A2(new_n518), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n840), .A2(new_n513), .A3(new_n520), .A4(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n843), .B(new_n512), .C1(new_n836), .C2(new_n837), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n839), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n624), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n823), .A2(new_n832), .A3(new_n835), .A4(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT115), .B1(new_n833), .B2(new_n834), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n812), .A2(new_n822), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n852), .A2(KEYINPUT117), .A3(new_n835), .A4(new_n846), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n662), .A2(new_n855), .A3(new_n845), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n839), .A2(new_n842), .A3(new_n844), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT118), .B1(new_n738), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n823), .A2(new_n832), .A3(new_n524), .A4(new_n835), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n627), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n576), .B1(new_n854), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n625), .A2(new_n525), .A3(new_n628), .A4(new_n662), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AND4_X1   g663(.A1(new_n348), .A2(new_n864), .A3(new_n399), .A4(new_n765), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n865), .A2(new_n751), .ZN(new_n866));
  AOI21_X1  g665(.A(G113gat), .B1(new_n866), .B2(new_n524), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n678), .B1(new_n862), .B2(new_n863), .ZN(new_n868));
  INV_X1    g667(.A(new_n751), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n869), .A2(new_n665), .A3(new_n716), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n524), .A2(G113gat), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n867), .B1(new_n871), .B2(new_n872), .ZN(G1340gat));
  AOI21_X1  g672(.A(G120gat), .B1(new_n866), .B2(new_n738), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n738), .A2(G120gat), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n871), .B2(new_n875), .ZN(G1341gat));
  NAND3_X1  g675(.A1(new_n871), .A2(G127gat), .A3(new_n577), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT119), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n865), .A2(new_n577), .A3(new_n751), .ZN(new_n879));
  AOI21_X1  g678(.A(G127gat), .B1(new_n879), .B2(KEYINPUT120), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n879), .A2(KEYINPUT120), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(G1342gat));
  AND2_X1   g681(.A1(new_n871), .A2(new_n627), .ZN(new_n883));
  INV_X1    g682(.A(G134gat), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n668), .A2(new_n624), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n865), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n885), .B1(KEYINPUT56), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(KEYINPUT56), .B2(new_n887), .ZN(G1343gat));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n718), .A2(new_n869), .A3(new_n665), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT57), .B1(new_n864), .B2(new_n678), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n678), .A2(KEYINPUT57), .ZN(new_n893));
  XOR2_X1   g692(.A(KEYINPUT121), .B(KEYINPUT55), .Z(new_n894));
  NAND2_X1  g693(.A1(new_n833), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n895), .A2(new_n524), .A3(new_n812), .A4(new_n822), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n738), .A2(new_n857), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n627), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n576), .B1(new_n854), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n893), .B1(new_n899), .B2(new_n863), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n524), .B(new_n891), .C1(new_n892), .C2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n890), .B1(new_n901), .B2(G141gat), .ZN(new_n902));
  INV_X1    g701(.A(new_n459), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n665), .B1(new_n862), .B2(new_n863), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n525), .A2(G141gat), .ZN(new_n905));
  AND4_X1   g704(.A1(new_n903), .A2(new_n904), .A3(new_n751), .A4(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n906), .B1(new_n901), .B2(G141gat), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n902), .A2(new_n907), .A3(KEYINPUT58), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT58), .ZN(new_n909));
  AOI221_X4 g708(.A(new_n906), .B1(new_n890), .B2(new_n909), .C1(new_n901), .C2(G141gat), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n908), .A2(new_n910), .ZN(G1344gat));
  NAND2_X1  g710(.A1(new_n904), .A2(new_n903), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n912), .A2(new_n869), .ZN(new_n913));
  INV_X1    g712(.A(G148gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n913), .A2(new_n914), .A3(new_n738), .ZN(new_n915));
  XNOR2_X1  g714(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n893), .B1(new_n862), .B2(new_n863), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n896), .A2(new_n897), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n624), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n577), .B1(new_n919), .B2(new_n847), .ZN(new_n920));
  INV_X1    g719(.A(new_n863), .ZN(new_n921));
  OAI21_X1  g720(.A(KEYINPUT124), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n847), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n576), .B1(new_n923), .B2(new_n898), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(new_n925), .A3(new_n863), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n922), .A2(new_n926), .A3(new_n678), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT57), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n917), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n891), .A2(new_n738), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n914), .B1(new_n931), .B2(KEYINPUT125), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n933), .B1(new_n929), .B2(new_n930), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n916), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n891), .B1(new_n892), .B2(new_n900), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n936), .A2(new_n662), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n937), .A2(KEYINPUT59), .A3(new_n914), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n915), .B1(new_n935), .B2(new_n938), .ZN(G1345gat));
  OAI21_X1  g738(.A(G155gat), .B1(new_n936), .B2(new_n576), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n913), .A2(new_n209), .A3(new_n577), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1346gat));
  OAI21_X1  g741(.A(G162gat), .B1(new_n936), .B2(new_n624), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n886), .A2(new_n210), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n912), .B2(new_n944), .ZN(G1347gat));
  NOR2_X1   g744(.A1(new_n330), .A2(new_n348), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n947), .A2(new_n716), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n868), .A2(new_n948), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n949), .A2(new_n264), .A3(new_n525), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n348), .B1(new_n862), .B2(new_n863), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n765), .A2(new_n399), .A3(new_n869), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n953), .A2(KEYINPUT126), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(KEYINPUT126), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n954), .A2(new_n524), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n950), .B1(new_n956), .B2(new_n264), .ZN(G1348gat));
  OAI21_X1  g756(.A(G176gat), .B1(new_n949), .B2(new_n662), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n954), .A2(new_n955), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n738), .A2(new_n265), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(G1349gat));
  OAI21_X1  g760(.A(G183gat), .B1(new_n949), .B2(new_n576), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n577), .A2(new_n289), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n953), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g764(.A(G190gat), .B1(new_n949), .B2(new_n624), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n966), .A2(KEYINPUT61), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n966), .A2(KEYINPUT61), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n627), .A2(new_n290), .ZN(new_n969));
  OAI22_X1  g768(.A1(new_n967), .A2(new_n968), .B1(new_n959), .B2(new_n969), .ZN(G1351gat));
  NOR2_X1   g769(.A1(new_n459), .A2(new_n751), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n951), .A2(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(G197gat), .B1(new_n973), .B2(new_n524), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n718), .A2(new_n947), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n929), .A2(new_n976), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n524), .A2(G197gat), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(G1352gat));
  NOR3_X1   g778(.A1(new_n972), .A2(G204gat), .A3(new_n662), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT62), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n977), .A2(new_n738), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(G204gat), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n981), .A2(new_n983), .ZN(G1353gat));
  OR3_X1    g783(.A1(new_n972), .A2(new_n304), .A3(new_n576), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n977), .A2(new_n577), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n986), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT63), .B1(new_n986), .B2(G211gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(G1354gat));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n990));
  NOR3_X1   g789(.A1(new_n929), .A2(new_n624), .A3(new_n976), .ZN(new_n991));
  INV_X1    g790(.A(G218gat), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n627), .A2(new_n992), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n972), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n990), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  OAI221_X1 g795(.A(KEYINPUT127), .B1(new_n972), .B2(new_n994), .C1(new_n991), .C2(new_n992), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n996), .A2(new_n997), .ZN(G1355gat));
endmodule


