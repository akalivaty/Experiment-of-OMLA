//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n211), .A2(new_n212), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n202), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n218), .B1(new_n212), .B2(new_n211), .C1(new_n227), .C2(KEYINPUT1), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT64), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XOR2_X1   g0039(.A(G50), .B(G58), .Z(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT65), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  AND2_X1   g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  OAI21_X1  g0047(.A(KEYINPUT66), .B1(new_n247), .B2(new_n213), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT66), .ZN(new_n252));
  NAND4_X1  g0052(.A1(new_n251), .A2(new_n252), .A3(G1), .A4(G13), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n248), .A2(new_n250), .A3(G274), .A4(new_n253), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n248), .A2(G232), .A3(new_n253), .A4(new_n249), .ZN(new_n255));
  AOI21_X1  g0055(.A(KEYINPUT74), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(new_n255), .A3(KEYINPUT74), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n247), .A2(new_n213), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT68), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT68), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G1698), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(new_n266), .A3(G223), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G226), .A2(G1698), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n262), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G87), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n259), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n257), .A2(new_n258), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G169), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n276), .B1(G179), .B2(new_n274), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n213), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n280), .B1(G1), .B2(new_n207), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G13), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(G1), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G20), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n282), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT73), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT73), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n284), .A2(new_n291), .A3(new_n288), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G58), .ZN(new_n294));
  INV_X1    g0094(.A(G68), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(G20), .B1(new_n296), .B2(new_n201), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G159), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT3), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n270), .ZN(new_n303));
  NAND2_X1  g0103(.A1(KEYINPUT3), .A2(G33), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n303), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT67), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n260), .A2(new_n261), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT67), .B1(new_n303), .B2(new_n304), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n207), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT7), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n306), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n301), .B1(new_n312), .B2(new_n295), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT16), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n303), .A2(new_n207), .A3(new_n304), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n311), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n305), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n300), .B1(new_n318), .B2(G68), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n280), .B1(new_n319), .B2(KEYINPUT16), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n293), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n277), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT18), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n322), .B(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G200), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n273), .A2(new_n258), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(new_n256), .ZN(new_n327));
  INV_X1    g0127(.A(G190), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n257), .A2(new_n328), .A3(new_n258), .A4(new_n273), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n307), .B1(new_n260), .B2(new_n261), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n303), .A2(KEYINPUT67), .A3(new_n304), .ZN(new_n332));
  AOI21_X1  g0132(.A(G20), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n305), .B1(new_n333), .B2(KEYINPUT7), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n300), .B1(new_n334), .B2(G68), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n320), .B1(new_n335), .B2(KEYINPUT16), .ZN(new_n336));
  INV_X1    g0136(.A(new_n293), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT17), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n330), .A2(new_n336), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT75), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT75), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n321), .A2(new_n341), .A3(new_n338), .A4(new_n330), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n330), .A2(new_n336), .A3(new_n337), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT17), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT76), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n343), .A2(KEYINPUT76), .A3(new_n345), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n324), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n281), .A2(G50), .ZN(new_n351));
  INV_X1    g0151(.A(new_n287), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n351), .B1(G50), .B2(new_n352), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n298), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n207), .A2(G33), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n354), .B1(new_n282), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n279), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n259), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n331), .A2(new_n332), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n264), .A2(new_n266), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(G222), .B1(G77), .B2(new_n361), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT69), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n361), .B2(new_n263), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n331), .A2(new_n332), .A3(KEYINPUT69), .A4(G1698), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(G223), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n360), .B1(new_n364), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n254), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n248), .A2(new_n253), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(new_n250), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n370), .B1(G226), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G169), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n369), .A2(new_n374), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G179), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n359), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n358), .B(KEYINPUT9), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n377), .B2(new_n325), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n369), .A2(new_n328), .A3(new_n374), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT10), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n375), .A2(G200), .ZN(new_n384));
  INV_X1    g0184(.A(new_n382), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT10), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .A4(new_n380), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n379), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n352), .A2(G77), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n389), .B1(new_n281), .B2(G77), .ZN(new_n390));
  XOR2_X1   g0190(.A(new_n282), .B(KEYINPUT70), .Z(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n298), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT15), .B(G87), .ZN(new_n393));
  OAI221_X1 g0193(.A(new_n392), .B1(new_n207), .B2(new_n221), .C1(new_n355), .C2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n390), .B1(new_n394), .B2(new_n279), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n366), .A2(G238), .A3(new_n367), .ZN(new_n396));
  AND3_X1   g0196(.A1(new_n331), .A2(new_n332), .A3(G232), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT68), .B(G1698), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n397), .A2(new_n398), .B1(G107), .B2(new_n361), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n360), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n370), .B1(G244), .B2(new_n372), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n325), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n400), .A2(G190), .A3(new_n402), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n395), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(G179), .ZN(new_n408));
  OR3_X1    g0208(.A1(new_n400), .A2(new_n408), .A3(new_n402), .ZN(new_n409));
  OAI21_X1  g0209(.A(G169), .B1(new_n400), .B2(new_n402), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n395), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n388), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n248), .A2(G238), .A3(new_n253), .A4(new_n249), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n254), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n331), .A2(new_n332), .A3(G226), .A4(new_n398), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n331), .A2(new_n332), .A3(G232), .A4(G1698), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G97), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n415), .B1(new_n419), .B2(new_n259), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT13), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI211_X1 g0222(.A(KEYINPUT13), .B(new_n415), .C1(new_n419), .C2(new_n259), .ZN(new_n423));
  OAI21_X1  g0223(.A(G169), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT14), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT14), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n426), .B(G169), .C1(new_n422), .C2(new_n423), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n422), .A2(KEYINPUT71), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n420), .A2(new_n421), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT71), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n420), .B2(new_n421), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n428), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n425), .B(new_n427), .C1(new_n432), .C2(new_n408), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT12), .ZN(new_n434));
  INV_X1    g0234(.A(new_n286), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n295), .A2(G20), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n286), .A2(KEYINPUT12), .A3(G20), .A4(new_n295), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n437), .B(new_n438), .C1(new_n281), .C2(new_n295), .ZN(new_n439));
  XOR2_X1   g0239(.A(new_n439), .B(KEYINPUT72), .Z(new_n440));
  NAND2_X1  g0240(.A1(new_n298), .A2(G50), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(new_n436), .C1(new_n221), .C2(new_n355), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n279), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n443), .B(KEYINPUT11), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n433), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n445), .ZN(new_n447));
  OAI21_X1  g0247(.A(G200), .B1(new_n422), .B2(new_n423), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n447), .B(new_n448), .C1(new_n432), .C2(new_n328), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n350), .A2(new_n413), .A3(KEYINPUT77), .A4(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT77), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n322), .B(KEYINPUT18), .ZN(new_n454));
  AOI221_X4 g0254(.A(new_n347), .B1(KEYINPUT17), .B2(new_n344), .C1(new_n340), .C2(new_n342), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT76), .B1(new_n343), .B2(new_n345), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n388), .A2(new_n446), .A3(new_n449), .A4(new_n412), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n453), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G107), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G20), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n435), .A2(new_n462), .ZN(new_n463));
  XOR2_X1   g0263(.A(new_n463), .B(KEYINPUT25), .Z(new_n464));
  OAI211_X1 g0264(.A(new_n280), .B(new_n287), .C1(G1), .C2(new_n270), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(new_n461), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n462), .B(KEYINPUT23), .ZN(new_n468));
  INV_X1    g0268(.A(G116), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n270), .A2(new_n469), .A3(G20), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n303), .A2(new_n304), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(new_n207), .A3(G87), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(KEYINPUT87), .A3(KEYINPUT22), .ZN(new_n474));
  OR3_X1    g0274(.A1(new_n271), .A2(KEYINPUT22), .A3(G20), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n474), .B1(new_n361), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT87), .B1(new_n473), .B2(KEYINPUT22), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n471), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT24), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n279), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n477), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n481), .B(new_n474), .C1(new_n361), .C2(new_n475), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT24), .B1(new_n482), .B2(new_n471), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n467), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n371), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT88), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT5), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G41), .ZN(new_n488));
  INV_X1    g0288(.A(G41), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT5), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n488), .A2(new_n490), .A3(new_n206), .A4(G45), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n485), .A2(new_n486), .A3(G264), .A4(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n264), .A2(new_n266), .A3(G250), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G257), .A2(G1698), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n262), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(G294), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n270), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n259), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(G274), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n206), .A2(G45), .ZN(new_n500));
  AOI211_X1 g0300(.A(new_n499), .B(new_n500), .C1(new_n487), .C2(G41), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT79), .ZN(new_n502));
  XNOR2_X1  g0302(.A(new_n490), .B(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n485), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n491), .A2(new_n248), .A3(G264), .A4(new_n253), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT88), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n492), .A2(new_n498), .A3(new_n504), .A4(new_n506), .ZN(new_n507));
  OR2_X1    g0307(.A1(new_n507), .A2(G190), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n492), .A2(new_n498), .A3(new_n506), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT89), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT89), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n492), .A2(new_n498), .A3(new_n511), .A4(new_n506), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n504), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n325), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n484), .B1(new_n508), .B2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n510), .A2(G179), .A3(new_n504), .A4(new_n512), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n507), .A2(G169), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n484), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT90), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n484), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n514), .A2(new_n508), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT90), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n484), .A2(new_n518), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  MUX2_X1   g0327(.A(new_n287), .B(new_n465), .S(G97), .Z(new_n528));
  INV_X1    g0328(.A(KEYINPUT6), .ZN(new_n529));
  INV_X1    g0329(.A(G97), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(new_n461), .ZN(new_n531));
  NOR2_X1   g0331(.A1(G97), .A2(G107), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n461), .A2(KEYINPUT6), .A3(G97), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G20), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n298), .A2(G77), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(G107), .B2(new_n334), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n528), .B1(new_n539), .B2(new_n280), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT78), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n264), .A2(new_n266), .A3(G244), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n541), .B1(new_n542), .B2(new_n262), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n472), .A2(new_n398), .A3(KEYINPUT78), .A4(G244), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT4), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n308), .A2(new_n309), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G250), .A2(G1698), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n542), .B2(new_n545), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G283), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n546), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n259), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n485), .A2(G257), .A3(new_n491), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n504), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n325), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n540), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n553), .A2(new_n556), .A3(KEYINPUT80), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT80), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n547), .A2(new_n549), .B1(G33), .B2(G283), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n360), .B1(new_n561), .B2(new_n546), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n560), .B1(new_n562), .B2(new_n555), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n559), .A2(new_n563), .A3(G190), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(G169), .B1(new_n559), .B2(new_n563), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n553), .A2(new_n556), .A3(new_n408), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n540), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n565), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n465), .A2(new_n271), .ZN(new_n570));
  INV_X1    g0370(.A(new_n393), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n571), .A2(new_n287), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT19), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n207), .B1(new_n418), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(G87), .A2(G97), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n461), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n575), .A2(new_n577), .B1(new_n574), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n472), .A2(new_n207), .A3(G68), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(KEYINPUT82), .B(new_n573), .C1(new_n581), .C2(new_n280), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT82), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n280), .B1(new_n579), .B2(new_n580), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n583), .B1(new_n584), .B2(new_n572), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n570), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n500), .A2(G250), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n499), .B2(new_n500), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n485), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G244), .A2(G1698), .ZN(new_n590));
  OAI22_X1  g0390(.A1(new_n262), .A2(new_n590), .B1(new_n270), .B2(new_n469), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT81), .ZN(new_n592));
  OAI21_X1  g0392(.A(G238), .B1(new_n260), .B2(new_n261), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n593), .B2(new_n362), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n472), .A2(new_n398), .A3(KEYINPUT81), .A4(G238), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n591), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n589), .B1(new_n596), .B2(new_n360), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G200), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n586), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT83), .ZN(new_n600));
  INV_X1    g0400(.A(new_n597), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(G190), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT83), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n586), .A2(new_n603), .A3(new_n598), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n600), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n582), .A2(new_n585), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n393), .B2(new_n465), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n597), .A2(new_n275), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n601), .A2(new_n408), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n270), .A2(G97), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(new_n207), .A3(new_n551), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT86), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT86), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n612), .A2(new_n615), .A3(new_n207), .A4(new_n551), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT85), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n279), .B(new_n618), .C1(new_n207), .C2(G116), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n207), .A2(G116), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT85), .B1(new_n280), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n617), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT20), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n617), .A2(new_n621), .A3(KEYINPUT20), .A4(new_n619), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  MUX2_X1   g0426(.A(new_n287), .B(new_n465), .S(G116), .Z(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(G303), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n331), .B2(new_n332), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n264), .A2(new_n266), .A3(G257), .ZN(new_n631));
  NAND2_X1  g0431(.A1(G264), .A2(G1698), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n262), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n259), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT84), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n485), .A2(new_n635), .A3(G270), .A4(new_n491), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n491), .A2(new_n248), .A3(G270), .A4(new_n253), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT84), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n634), .A2(new_n636), .A3(new_n504), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(G169), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT21), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n639), .A2(new_n408), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n628), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n628), .ZN(new_n645));
  INV_X1    g0445(.A(new_n639), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(G200), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n639), .A2(G190), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n641), .B1(new_n645), .B2(new_n640), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n644), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n569), .A2(new_n611), .A3(new_n651), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n460), .A2(new_n527), .A3(new_n652), .ZN(G372));
  NAND2_X1  g0453(.A1(new_n348), .A2(new_n349), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n445), .A2(new_n433), .B1(new_n449), .B2(new_n411), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n454), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n383), .A2(new_n387), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n379), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n460), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n525), .A2(new_n650), .A3(new_n644), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n559), .A2(new_n563), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n275), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n540), .A2(new_n567), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n663), .A2(new_n664), .B1(new_n558), .B2(new_n564), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n602), .A2(new_n598), .A3(new_n586), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n661), .A2(new_n665), .A3(new_n523), .A4(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n608), .A2(KEYINPUT91), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n608), .A2(KEYINPUT91), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n609), .B(new_n607), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n566), .A2(new_n568), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n672), .A2(new_n605), .A3(KEYINPUT26), .A4(new_n610), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT92), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n672), .A2(new_n666), .A3(new_n670), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n673), .A2(KEYINPUT92), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n671), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n659), .B1(new_n660), .B2(new_n678), .ZN(G369));
  OR3_X1    g0479(.A1(new_n435), .A2(KEYINPUT27), .A3(G20), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT27), .B1(new_n435), .B2(G20), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n680), .A2(G213), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G343), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT93), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n527), .B1(new_n521), .B2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n684), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n519), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n644), .A2(new_n650), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n684), .A2(new_n645), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n693), .B1(new_n651), .B2(new_n692), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(G330), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n689), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n690), .A2(new_n684), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n685), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n519), .A2(new_n684), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n699), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n210), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n576), .A2(new_n461), .A3(new_n469), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n707), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n216), .B2(new_n707), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n678), .B2(new_n686), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n675), .A2(KEYINPUT26), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n672), .A2(new_n605), .A3(new_n676), .A4(new_n610), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n667), .A2(new_n715), .A3(new_n670), .A4(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(KEYINPUT29), .A3(new_n684), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n646), .A2(new_n601), .A3(G179), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n553), .A2(new_n556), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(new_n513), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n643), .A2(new_n510), .A3(new_n512), .A4(new_n601), .ZN(new_n725));
  OAI21_X1  g0525(.A(KEYINPUT94), .B1(new_n725), .B2(new_n662), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI211_X1 g0528(.A(KEYINPUT94), .B(KEYINPUT30), .C1(new_n725), .C2(new_n662), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n724), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n720), .B1(new_n730), .B2(new_n684), .ZN(new_n731));
  INV_X1    g0531(.A(new_n729), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n510), .A2(new_n512), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n639), .A2(new_n597), .A3(new_n408), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n733), .A2(new_n563), .A3(new_n559), .A4(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(KEYINPUT30), .B1(new_n735), .B2(KEYINPUT94), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n723), .B1(new_n732), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(KEYINPUT31), .A3(new_n686), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n731), .A2(new_n738), .A3(KEYINPUT95), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n652), .A2(new_n520), .A3(new_n526), .A4(new_n684), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(KEYINPUT95), .B1(new_n731), .B2(new_n738), .ZN(new_n742));
  OAI21_X1  g0542(.A(G330), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n719), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n712), .B1(new_n744), .B2(G1), .ZN(G364));
  NOR2_X1   g0545(.A1(new_n285), .A2(G20), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G45), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n707), .A2(G1), .A3(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT96), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n695), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n213), .B1(G20), .B2(new_n275), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n705), .A2(new_n472), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n241), .A2(G45), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n217), .A2(G45), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n705), .A2(new_n361), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n762), .A2(G355), .B1(new_n469), .B2(new_n705), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n757), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n408), .A2(new_n325), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n207), .A2(G190), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(KEYINPUT33), .B(G317), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n207), .A2(new_n328), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n408), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n768), .A2(new_n769), .B1(new_n773), .B2(G322), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n325), .A2(G179), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G179), .A2(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n766), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G303), .A2(new_n777), .B1(new_n780), .B2(G329), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n774), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n207), .B1(new_n778), .B2(G190), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n547), .B(new_n782), .C1(G294), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n770), .A2(new_n765), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n766), .A2(new_n771), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G326), .A2(new_n787), .B1(new_n789), .B2(G311), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n775), .A2(new_n766), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n785), .B(new_n790), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G159), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n779), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT32), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n784), .A2(G97), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n786), .A2(new_n202), .B1(new_n772), .B2(new_n294), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n767), .A2(new_n295), .B1(new_n788), .B2(new_n221), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n776), .A2(new_n271), .B1(new_n792), .B2(new_n461), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n361), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n796), .A2(new_n797), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n793), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n764), .B1(new_n804), .B2(new_n755), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n748), .B1(new_n754), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n695), .A2(new_n696), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n698), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n806), .B1(new_n808), .B2(new_n748), .ZN(G396));
  NOR2_X1   g0609(.A1(new_n678), .A2(new_n686), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n411), .A2(new_n684), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n395), .A2(new_n684), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n407), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g0613(.A(KEYINPUT99), .B(new_n811), .C1(new_n813), .C2(new_n411), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT99), .ZN(new_n815));
  INV_X1    g0615(.A(new_n812), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n411), .B1(new_n816), .B2(new_n406), .ZN(new_n817));
  INV_X1    g0617(.A(new_n811), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n815), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n810), .B(new_n820), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n821), .A2(new_n743), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT100), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  INV_X1    g0625(.A(new_n748), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n821), .B2(new_n743), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n824), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n755), .ZN(new_n829));
  INV_X1    g0629(.A(G143), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n772), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G137), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n786), .A2(new_n832), .B1(new_n788), .B2(new_n794), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n831), .B(new_n833), .C1(G150), .C2(new_n768), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n834), .A2(KEYINPUT34), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(KEYINPUT34), .ZN(new_n836));
  INV_X1    g0636(.A(G132), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n472), .B1(new_n779), .B2(new_n837), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n776), .A2(new_n202), .B1(new_n792), .B2(new_n295), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n838), .B(new_n839), .C1(G58), .C2(new_n784), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n835), .A2(new_n836), .A3(new_n840), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G294), .A2(new_n773), .B1(new_n780), .B2(G311), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n271), .B2(new_n792), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT97), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n767), .A2(new_n791), .B1(new_n788), .B2(new_n469), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(G303), .A2(new_n787), .B1(new_n777), .B2(G107), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n847), .A2(new_n361), .A3(new_n797), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n846), .B(new_n848), .C1(new_n844), .C2(new_n845), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n829), .B1(new_n841), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n755), .A2(new_n749), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n748), .B(new_n850), .C1(new_n221), .C2(new_n851), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT98), .Z(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n750), .B2(new_n820), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n828), .A2(new_n854), .ZN(G384));
  NOR2_X1   g0655(.A1(new_n446), .A2(new_n686), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT39), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT38), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT103), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n320), .B1(KEYINPUT16), .B2(new_n319), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n337), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT102), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n861), .B(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n682), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n457), .A2(new_n859), .A3(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  INV_X1    g0667(.A(new_n682), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n277), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n863), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n867), .B1(new_n870), .B2(new_n344), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n336), .A2(new_n337), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n682), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n874), .B(KEYINPUT104), .Z(new_n875));
  INV_X1    g0675(.A(new_n344), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n322), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n872), .B1(new_n878), .B2(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n866), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n859), .B1(new_n457), .B2(new_n865), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n858), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT103), .B1(new_n350), .B2(new_n864), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n883), .A2(KEYINPUT38), .A3(new_n866), .A4(new_n879), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n857), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n878), .B(new_n867), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n875), .B1(new_n454), .B2(new_n346), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n858), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  XOR2_X1   g0688(.A(KEYINPUT105), .B(KEYINPUT39), .Z(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n888), .A2(new_n884), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n856), .B1(new_n885), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n447), .A2(new_n684), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n450), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n450), .A2(new_n893), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n810), .A2(new_n820), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n897), .B1(new_n898), .B2(new_n811), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n882), .A2(new_n884), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n899), .A2(new_n900), .B1(new_n324), .B2(new_n868), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n892), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT106), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT106), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n892), .A2(new_n904), .A3(new_n901), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n714), .A2(new_n460), .A3(new_n718), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n659), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n906), .B(new_n908), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n894), .A2(new_n895), .B1(new_n819), .B2(new_n814), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n740), .A2(new_n731), .A3(new_n738), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(KEYINPUT40), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n884), .B2(new_n888), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n910), .A2(new_n911), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n874), .B(KEYINPUT104), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n916), .A2(new_n322), .A3(new_n876), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n871), .B1(new_n917), .B2(new_n867), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n864), .B1(new_n654), .B2(new_n454), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n918), .B1(new_n919), .B2(new_n859), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n920), .B2(new_n883), .ZN(new_n921));
  INV_X1    g0721(.A(new_n884), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n915), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT40), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n913), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n460), .A2(new_n911), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT107), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(G330), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n926), .B2(new_n928), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n909), .A2(new_n931), .B1(new_n206), .B2(new_n746), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n931), .B2(new_n909), .ZN(new_n933));
  OR3_X1    g0733(.A1(new_n216), .A2(new_n221), .A3(new_n296), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n202), .A2(G68), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n206), .B(G13), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n535), .B(KEYINPUT101), .Z(new_n937));
  OR2_X1    g0737(.A1(new_n937), .A2(KEYINPUT35), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(KEYINPUT35), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n938), .A2(G116), .A3(new_n214), .A4(new_n939), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT36), .Z(new_n941));
  OR3_X1    g0741(.A1(new_n933), .A2(new_n936), .A3(new_n941), .ZN(G367));
  NAND2_X1  g0742(.A1(new_n686), .A2(new_n540), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n665), .A2(new_n943), .ZN(new_n944));
  OR3_X1    g0744(.A1(new_n701), .A2(KEYINPUT42), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(KEYINPUT42), .B1(new_n701), .B2(new_n944), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n944), .A2(new_n525), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n684), .B1(new_n947), .B2(new_n672), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n684), .A2(new_n586), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n670), .B2(new_n666), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n670), .B2(new_n950), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT108), .Z(new_n953));
  INV_X1    g0753(.A(KEYINPUT43), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n949), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n699), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n672), .A2(new_n686), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n944), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n949), .A2(new_n962), .A3(new_n955), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n956), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n961), .B1(new_n956), .B2(new_n963), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n706), .B(KEYINPUT41), .Z(new_n967));
  INV_X1    g0767(.A(KEYINPUT45), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n703), .B2(new_n960), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n701), .A2(KEYINPUT45), .A3(new_n702), .A4(new_n959), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n959), .B1(new_n701), .B2(new_n702), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT44), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n971), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n699), .A2(KEYINPUT109), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n700), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n701), .B1(new_n688), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(new_n697), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n744), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n972), .B(KEYINPUT44), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n985), .A2(new_n971), .A3(new_n977), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n979), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n967), .B1(new_n987), .B2(new_n744), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n747), .A2(G1), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n966), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n237), .A2(new_n705), .A3(new_n472), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n756), .B1(new_n210), .B2(new_n393), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n776), .A2(new_n469), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(KEYINPUT46), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT111), .Z(new_n995));
  OAI22_X1  g0795(.A1(new_n772), .A2(new_n629), .B1(new_n788), .B2(new_n791), .ZN(new_n996));
  XNOR2_X1  g0796(.A(KEYINPUT110), .B(G311), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n996), .B1(new_n787), .B2(new_n998), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n767), .A2(new_n496), .B1(new_n792), .B2(new_n530), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n472), .B(new_n1000), .C1(G317), .C2(new_n780), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n993), .A2(KEYINPUT46), .B1(G107), .B2(new_n784), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n995), .A2(new_n999), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT112), .Z(new_n1004));
  NOR2_X1   g0804(.A1(new_n792), .A2(new_n221), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n786), .A2(new_n830), .B1(new_n767), .B2(new_n794), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(G150), .C2(new_n773), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n776), .A2(new_n294), .B1(new_n788), .B2(new_n202), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(G137), .B2(new_n780), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n783), .A2(new_n295), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1007), .A2(new_n547), .A3(new_n1009), .A4(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT113), .Z(new_n1013));
  NAND3_X1  g0813(.A1(new_n1004), .A2(KEYINPUT47), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n755), .ZN(new_n1015));
  AOI21_X1  g0815(.A(KEYINPUT47), .B1(new_n1004), .B2(new_n1013), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n826), .B1(new_n991), .B2(new_n992), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT114), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n752), .B2(new_n952), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n990), .A2(new_n1019), .ZN(G387));
  AOI22_X1  g0820(.A1(new_n777), .A2(G294), .B1(new_n784), .B2(G283), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n787), .A2(G322), .B1(new_n768), .B2(new_n998), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT116), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G317), .A2(new_n773), .B1(new_n789), .B2(G303), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT48), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1021), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n1026), .B2(new_n1025), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1028), .A2(KEYINPUT49), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(KEYINPUT49), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n262), .B1(new_n792), .B2(new_n469), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G326), .B2(new_n780), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n786), .A2(new_n794), .B1(new_n776), .B2(new_n221), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n767), .A2(new_n282), .B1(new_n788), .B2(new_n295), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n784), .A2(new_n571), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n792), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n262), .B1(new_n1038), .B2(G97), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G50), .A2(new_n773), .B1(new_n780), .B2(G150), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1036), .A2(new_n1037), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n829), .B1(new_n1033), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n391), .A2(new_n202), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT50), .Z(new_n1044));
  AOI21_X1  g0844(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1044), .A2(new_n709), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(G45), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1046), .B(new_n758), .C1(new_n233), .C2(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n762), .A2(new_n708), .B1(new_n461), .B2(new_n705), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1048), .A2(KEYINPUT115), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n756), .ZN(new_n1051));
  AOI21_X1  g0851(.A(KEYINPUT115), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n826), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1042), .B(new_n1053), .C1(new_n689), .C2(new_n753), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n982), .B2(new_n989), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n983), .A2(new_n706), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n982), .A2(new_n744), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1055), .B1(new_n1056), .B2(new_n1057), .ZN(G393));
  AOI22_X1  g0858(.A1(G317), .A2(new_n787), .B1(new_n773), .B2(G311), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT52), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n776), .A2(new_n791), .B1(new_n788), .B2(new_n496), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G303), .B2(new_n768), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n784), .A2(G116), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G107), .A2(new_n1038), .B1(new_n780), .B2(G322), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1062), .A2(new_n361), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n783), .A2(new_n221), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n262), .B(new_n1066), .C1(G87), .C2(new_n1038), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n391), .A2(new_n789), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n776), .A2(new_n295), .B1(new_n779), .B2(new_n830), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G50), .B2(new_n768), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(G150), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n786), .A2(new_n1072), .B1(new_n772), .B2(new_n794), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT51), .Z(new_n1074));
  OAI22_X1  g0874(.A1(new_n1060), .A2(new_n1065), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n755), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n758), .A2(new_n245), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n756), .B1(new_n530), .B2(new_n210), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1076), .B(new_n826), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n960), .B2(new_n751), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n976), .A2(new_n957), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n985), .A2(new_n699), .A3(new_n971), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n989), .ZN(new_n1085));
  OAI211_X1 g0885(.A(KEYINPUT117), .B(new_n1081), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT117), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1085), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1087), .B1(new_n1088), .B2(new_n1080), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n987), .A2(new_n706), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1084), .A2(new_n983), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1086), .A2(new_n1089), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(G390));
  NOR2_X1   g0893(.A1(new_n885), .A2(new_n891), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n856), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n818), .B1(new_n810), .B2(new_n820), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1095), .B1(new_n1096), .B2(new_n897), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n888), .A2(new_n884), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n717), .A2(new_n684), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n818), .B1(new_n1101), .B2(new_n820), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1095), .B1(new_n1102), .B2(new_n897), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(G330), .B(new_n910), .C1(new_n741), .C2(new_n742), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1098), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1104), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n696), .B1(new_n814), .B2(new_n819), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n911), .A2(new_n896), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1107), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n911), .A2(new_n1109), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n897), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1106), .A2(new_n1114), .A3(new_n1102), .ZN(new_n1115));
  OAI211_X1 g0915(.A(G330), .B(new_n820), .C1(new_n741), .C2(new_n742), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1110), .B1(new_n1116), .B2(new_n897), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1117), .B2(new_n1096), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n460), .A2(G330), .A3(new_n911), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n907), .A2(new_n1119), .A3(new_n659), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1112), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1122), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1107), .B(new_n1124), .C1(new_n1108), .C2(new_n1111), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1123), .A2(new_n706), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n851), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT54), .B(G143), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n767), .A2(new_n832), .B1(new_n788), .B2(new_n1128), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n361), .B(new_n1129), .C1(G159), .C2(new_n784), .ZN(new_n1130));
  INV_X1    g0930(.A(G128), .ZN(new_n1131));
  INV_X1    g0931(.A(G125), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n786), .A2(new_n1131), .B1(new_n779), .B2(new_n1132), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n772), .A2(new_n837), .B1(new_n792), .B2(new_n202), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT53), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n776), .B2(new_n1072), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n777), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1133), .B(new_n1134), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n776), .A2(new_n271), .B1(new_n792), .B2(new_n295), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n767), .A2(new_n461), .B1(new_n779), .B2(new_n496), .ZN(new_n1140));
  NOR4_X1   g0940(.A1(new_n1139), .A2(new_n1140), .A3(new_n547), .A4(new_n1066), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n772), .A2(new_n469), .B1(new_n788), .B2(new_n530), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G283), .B2(new_n787), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1130), .A2(new_n1138), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n826), .B1(new_n283), .B2(new_n1127), .C1(new_n1144), .C2(new_n829), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(new_n1094), .B2(new_n749), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT118), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1146), .B(new_n1147), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1107), .B(new_n989), .C1(new_n1111), .C2(new_n1108), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1148), .A2(new_n1149), .A3(KEYINPUT119), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT119), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1126), .B1(new_n1150), .B2(new_n1151), .ZN(G378));
  NOR2_X1   g0952(.A1(new_n472), .A2(G41), .ZN(new_n1153));
  AOI211_X1 g0953(.A(G50), .B(new_n1153), .C1(new_n270), .C2(new_n489), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1153), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n788), .A2(new_n393), .B1(new_n779), .B2(new_n791), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1155), .B(new_n1156), .C1(G107), .C2(new_n773), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(G77), .A2(new_n777), .B1(new_n768), .B2(G97), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(G116), .A2(new_n787), .B1(new_n1038), .B2(G58), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1157), .A2(new_n1011), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1154), .B1(new_n1161), .B2(KEYINPUT58), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n786), .A2(new_n1132), .B1(new_n767), .B2(new_n837), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1128), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1164), .A2(new_n777), .B1(new_n773), .B2(G128), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n832), .B2(new_n788), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1163), .B(new_n1166), .C1(G150), .C2(new_n784), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n270), .B(new_n489), .C1(new_n792), .C2(new_n794), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(G124), .B2(new_n780), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT59), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1171), .B1(new_n1167), .B2(new_n1172), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1162), .B1(KEYINPUT58), .B2(new_n1161), .C1(new_n1169), .C2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n755), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n748), .B1(new_n202), .B2(new_n851), .ZN(new_n1176));
  OR2_X1    g0976(.A1(new_n388), .A2(KEYINPUT120), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n388), .A2(KEYINPUT120), .ZN(new_n1178));
  AND4_X1   g0978(.A1(new_n358), .A2(new_n1177), .A3(new_n682), .A4(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1177), .A2(new_n1178), .B1(new_n358), .B2(new_n682), .ZN(new_n1180));
  XOR2_X1   g0980(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1181));
  OR3_X1    g0981(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1181), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1175), .B(new_n1176), .C1(new_n1184), .C2(new_n750), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n925), .A2(KEYINPUT121), .A3(G330), .A4(new_n1184), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT121), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n912), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1099), .A2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n914), .B1(new_n882), .B2(new_n884), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1190), .B(G330), .C1(new_n1191), .C2(KEYINPUT40), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1184), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1188), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1187), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n892), .A2(new_n904), .A3(new_n901), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n904), .B1(new_n892), .B2(new_n901), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1198), .A2(new_n1199), .A3(KEYINPUT122), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1187), .A2(new_n1194), .B1(new_n1193), .B2(new_n1192), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT122), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n903), .A2(new_n1203), .A3(new_n905), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1201), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1186), .B1(new_n1206), .B2(new_n989), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT57), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n1125), .B2(new_n1121), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1202), .A2(new_n906), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1202), .A2(new_n906), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1209), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n706), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1125), .A2(new_n1121), .ZN(new_n1214));
  AOI21_X1  g1014(.A(KEYINPUT57), .B1(new_n1206), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1207), .B1(new_n1213), .B2(new_n1215), .ZN(G375));
  INV_X1    g1016(.A(new_n967), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1120), .B(new_n1115), .C1(new_n1117), .C2(new_n1096), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1122), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n897), .A2(new_n749), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n826), .B1(G68), .B2(new_n1127), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT123), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n786), .A2(new_n837), .B1(new_n772), .B2(new_n832), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n262), .B(new_n1223), .C1(G58), .C2(new_n1038), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G159), .A2(new_n777), .B1(new_n768), .B2(new_n1164), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(G150), .A2(new_n789), .B1(new_n780), .B2(G128), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n784), .A2(G50), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n776), .A2(new_n530), .B1(new_n788), .B2(new_n461), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1005), .B(new_n1229), .C1(G294), .C2(new_n787), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n469), .A2(new_n767), .B1(new_n772), .B2(new_n791), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G303), .B2(new_n780), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1230), .A2(new_n361), .A3(new_n1037), .A4(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n829), .B1(new_n1228), .B2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1222), .A2(new_n1234), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1118), .A2(new_n989), .B1(new_n1220), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1219), .A2(new_n1236), .ZN(G381));
  AND2_X1   g1037(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1126), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(G375), .A2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1092), .A2(new_n990), .A3(new_n1019), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NOR4_X1   g1043(.A1(G384), .A2(G393), .A3(G381), .A4(G396), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1241), .A2(new_n1243), .A3(new_n1244), .ZN(G407));
  INV_X1    g1045(.A(G213), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1246), .A2(G343), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1241), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(G407), .A2(new_n1248), .A3(G213), .ZN(new_n1249));
  XOR2_X1   g1049(.A(new_n1249), .B(KEYINPUT124), .Z(G409));
  OAI211_X1 g1050(.A(G378), .B(new_n1207), .C1(new_n1213), .C2(new_n1215), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1217), .B(new_n1214), .C1(new_n1252), .C2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n989), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n1185), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1239), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1251), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1247), .ZN(new_n1259));
  INV_X1    g1059(.A(G384), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT60), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1218), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT125), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1262), .A2(new_n1263), .A3(new_n1122), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1263), .B1(new_n1262), .B2(new_n1122), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n706), .B1(new_n1218), .B2(new_n1261), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1236), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1260), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1262), .A2(new_n1122), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(KEYINPUT125), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1262), .A2(new_n1263), .A3(new_n1122), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1266), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(G384), .A3(new_n1236), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1269), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1258), .A2(new_n1259), .A3(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(KEYINPUT62), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1247), .B1(new_n1251), .B2(new_n1257), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1247), .A2(G2897), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1274), .A2(G384), .A3(new_n1236), .ZN(new_n1282));
  AOI21_X1  g1082(.A(G384), .B1(new_n1274), .B2(new_n1236), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT126), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT126), .B1(new_n1269), .B2(new_n1275), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1281), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1284), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1269), .A2(KEYINPUT126), .A3(new_n1275), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1288), .A2(new_n1289), .A3(G2897), .A4(new_n1247), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1291));
  OR2_X1    g1091(.A1(new_n1280), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT61), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT62), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1280), .A2(new_n1294), .A3(new_n1277), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1279), .A2(new_n1292), .A3(new_n1293), .A4(new_n1295), .ZN(new_n1296));
  XOR2_X1   g1096(.A(G393), .B(G396), .Z(new_n1297));
  AOI21_X1  g1097(.A(new_n1092), .B1(new_n990), .B2(new_n1019), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1297), .B1(new_n1243), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G390), .A2(G387), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1297), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(new_n1242), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1296), .A2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(KEYINPUT63), .B1(new_n1280), .B2(new_n1291), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1278), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1299), .A2(new_n1293), .A3(new_n1302), .ZN(new_n1307));
  AOI211_X1 g1107(.A(new_n1247), .B(new_n1276), .C1(new_n1251), .C2(new_n1257), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1307), .B1(new_n1308), .B2(KEYINPUT63), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1306), .A2(new_n1309), .A3(KEYINPUT127), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT127), .B1(new_n1306), .B2(new_n1309), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1304), .B1(new_n1310), .B2(new_n1311), .ZN(G405));
  NAND2_X1  g1112(.A1(new_n1303), .A2(new_n1276), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1299), .A2(new_n1277), .A3(new_n1302), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(G375), .A2(new_n1239), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1251), .ZN(new_n1317));
  XOR2_X1   g1117(.A(new_n1315), .B(new_n1317), .Z(G402));
endmodule


