//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1291,
    new_n1292, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1366, new_n1367, new_n1368;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n210), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n212), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n215), .B(new_n221), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G116), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n209), .A2(G33), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND4_X1  g0052(.A1(new_n247), .A2(new_n251), .A3(new_n219), .A4(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n250), .B1(new_n253), .B2(new_n249), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G283), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT77), .B(G97), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n210), .B(new_n255), .C1(new_n256), .C2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n252), .A2(new_n219), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT81), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n249), .A2(G20), .ZN(new_n260));
  AND3_X1   g0060(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n259), .B1(new_n258), .B2(new_n260), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n257), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n257), .B(KEYINPUT20), .C1(new_n261), .C2(new_n262), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n254), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G1), .A3(G13), .ZN(new_n269));
  INV_X1    g0069(.A(G45), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(G1), .ZN(new_n271));
  AND3_X1   g0071(.A1(new_n269), .A2(G274), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT5), .ZN(new_n273));
  OAI21_X1  g0073(.A(KEYINPUT78), .B1(new_n273), .B2(G41), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT78), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT5), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n273), .A2(G41), .ZN(new_n278));
  AND3_X1   g0078(.A1(new_n274), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n272), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G303), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(G264), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G257), .A2(G1698), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n282), .B(new_n284), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n269), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n287), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n276), .A2(KEYINPUT5), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n271), .A2(new_n294), .A3(new_n278), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(G270), .A3(new_n269), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n280), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G169), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n267), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT21), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT21), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(new_n267), .B2(new_n298), .ZN(new_n302));
  INV_X1    g0102(.A(new_n267), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n280), .A2(new_n293), .A3(G179), .A4(new_n296), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n297), .A2(G200), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n267), .B(new_n307), .C1(new_n308), .C2(new_n297), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n300), .A2(new_n302), .A3(new_n306), .A4(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT82), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n299), .A2(KEYINPUT21), .B1(new_n303), .B2(new_n305), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT82), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n312), .A2(new_n313), .A3(new_n302), .A4(new_n309), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT65), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(new_n210), .B2(G1), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n209), .A2(KEYINPUT65), .A3(G20), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n319), .A2(new_n248), .A3(new_n258), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT8), .B(G58), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT64), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G58), .ZN(new_n324));
  OR3_X1    g0124(.A1(new_n322), .A2(new_n324), .A3(KEYINPUT8), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n248), .B1(new_n323), .B2(new_n325), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n258), .ZN(new_n330));
  AND2_X1   g0130(.A1(G58), .A2(G68), .ZN(new_n331));
  OAI21_X1  g0131(.A(G20), .B1(new_n331), .B2(new_n201), .ZN(new_n332));
  INV_X1    g0132(.A(G159), .ZN(new_n333));
  NOR4_X1   g0133(.A1(new_n333), .A2(KEYINPUT72), .A3(G20), .A4(G33), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT72), .ZN(new_n335));
  NOR2_X1   g0135(.A1(G20), .A2(G33), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n335), .B1(new_n336), .B2(G159), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n332), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(G20), .B1(new_n282), .B2(new_n284), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT3), .B(G33), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n210), .A2(KEYINPUT7), .ZN(new_n341));
  OAI22_X1  g0141(.A1(new_n339), .A2(KEYINPUT7), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n338), .B1(new_n342), .B2(G68), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n330), .B1(new_n343), .B2(KEYINPUT16), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT16), .ZN(new_n345));
  INV_X1    g0145(.A(G68), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n283), .A2(KEYINPUT3), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n341), .B1(new_n347), .B2(KEYINPUT73), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT73), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n282), .A2(new_n284), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT7), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n340), .B2(G20), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n346), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n345), .B1(new_n354), .B2(new_n338), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n329), .B1(new_n344), .B2(new_n355), .ZN(new_n356));
  OR2_X1    g0156(.A1(G223), .A2(G1698), .ZN(new_n357));
  INV_X1    g0157(.A(G226), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G1698), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n282), .A2(new_n357), .A3(new_n284), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G33), .A2(G87), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n269), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(G1), .B1(new_n276), .B2(new_n270), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n363), .A2(new_n269), .A3(G274), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n269), .A2(G232), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G169), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(G179), .B2(new_n368), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT18), .B1(new_n356), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n337), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n336), .A2(new_n335), .A3(G159), .ZN(new_n374));
  XNOR2_X1  g0174(.A(G58), .B(G68), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n373), .A2(new_n374), .B1(new_n375), .B2(G20), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n341), .B1(new_n282), .B2(new_n284), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n281), .A2(G33), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n210), .B1(new_n347), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n377), .B1(new_n379), .B2(new_n352), .ZN(new_n380));
  OAI211_X1 g0180(.A(KEYINPUT16), .B(new_n376), .C1(new_n380), .C2(new_n346), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n282), .A2(new_n284), .A3(new_n349), .ZN(new_n382));
  OAI211_X1 g0182(.A(KEYINPUT7), .B(new_n210), .C1(new_n282), .C2(new_n349), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n382), .A2(new_n383), .B1(new_n339), .B2(KEYINPUT7), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n338), .B1(new_n384), .B2(G68), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n381), .B(new_n258), .C1(new_n385), .C2(KEYINPUT16), .ZN(new_n386));
  INV_X1    g0186(.A(new_n329), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT18), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n368), .A2(G179), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n369), .B2(new_n368), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n372), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(KEYINPUT74), .A2(KEYINPUT17), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(KEYINPUT74), .A2(KEYINPUT17), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n368), .A2(new_n308), .ZN(new_n398));
  INV_X1    g0198(.A(G200), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n362), .B2(new_n367), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n397), .B1(new_n356), .B2(new_n401), .ZN(new_n402));
  AND4_X1   g0202(.A1(new_n386), .A2(new_n387), .A3(new_n401), .A4(new_n394), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT75), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n386), .A2(new_n387), .A3(new_n401), .ZN(new_n405));
  INV_X1    g0205(.A(new_n397), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n356), .A2(new_n401), .A3(new_n394), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT75), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n393), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  OR2_X1    g0212(.A1(new_n412), .A2(KEYINPUT76), .ZN(new_n413));
  INV_X1    g0213(.A(new_n364), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n292), .A2(new_n363), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n414), .B1(G226), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(G222), .A2(G1698), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n288), .A2(G223), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n340), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n419), .B(new_n292), .C1(G77), .C2(new_n340), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n399), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n416), .A2(new_n420), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n421), .B1(G190), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT68), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT10), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n336), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n210), .A2(G33), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n426), .B1(new_n326), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n258), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT9), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n247), .A2(G50), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n320), .B2(G50), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n430), .B1(new_n429), .B2(new_n432), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n423), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n425), .A2(new_n436), .ZN(new_n437));
  OAI221_X1 g0237(.A(new_n423), .B1(new_n424), .B2(KEYINPUT10), .C1(new_n434), .C2(new_n435), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n422), .A2(G169), .ZN(new_n439));
  INV_X1    g0239(.A(G179), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n439), .B1(new_n440), .B2(new_n422), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n429), .A2(new_n432), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n437), .A2(new_n438), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n358), .A2(new_n288), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n232), .A2(G1698), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n282), .A2(new_n445), .A3(new_n284), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G33), .A2(G97), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n292), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n269), .A2(G238), .A3(new_n365), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n364), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT13), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n450), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n269), .B1(new_n447), .B2(new_n448), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n364), .A2(new_n451), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT13), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(new_n308), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT11), .ZN(new_n460));
  INV_X1    g0260(.A(G77), .ZN(new_n461));
  OAI22_X1  g0261(.A1(new_n427), .A2(new_n461), .B1(new_n210), .B2(G68), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT69), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n463), .B1(new_n336), .B2(G50), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n336), .A2(new_n463), .A3(G50), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n460), .B1(new_n467), .B2(new_n330), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT12), .B1(new_n247), .B2(G68), .ZN(new_n469));
  OR3_X1    g0269(.A1(new_n247), .A2(KEYINPUT12), .A3(G68), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n320), .A2(G68), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n466), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(new_n464), .ZN(new_n473));
  OAI211_X1 g0273(.A(KEYINPUT11), .B(new_n258), .C1(new_n473), .C2(new_n462), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n468), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n399), .B1(new_n454), .B2(new_n457), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n459), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n454), .A2(G179), .A3(new_n457), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT70), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n454), .A2(new_n457), .A3(KEYINPUT70), .A4(G179), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n458), .A2(G169), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT14), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT14), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n458), .A2(new_n485), .A3(G169), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT71), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n475), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n468), .A2(new_n471), .A3(new_n474), .A4(KEYINPUT71), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n477), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n340), .A2(G238), .A3(G1698), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n340), .A2(G232), .A3(new_n288), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n493), .B(new_n494), .C1(new_n206), .C2(new_n340), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n292), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n414), .B1(G244), .B2(new_n415), .ZN(new_n497));
  AOI21_X1  g0297(.A(G169), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT67), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n496), .A2(new_n497), .ZN(new_n500));
  OAI22_X1  g0300(.A1(new_n498), .A2(new_n499), .B1(new_n500), .B2(G179), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n496), .A2(KEYINPUT67), .A3(new_n440), .A4(new_n497), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n248), .A2(new_n461), .ZN(new_n503));
  XNOR2_X1  g0303(.A(new_n503), .B(KEYINPUT66), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n320), .A2(G77), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n210), .A2(new_n283), .ZN(new_n506));
  OAI22_X1  g0306(.A1(new_n321), .A2(new_n506), .B1(new_n210), .B2(new_n461), .ZN(new_n507));
  XNOR2_X1  g0307(.A(KEYINPUT15), .B(G87), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(new_n427), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n258), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n504), .A2(new_n505), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n501), .A2(new_n502), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n511), .B1(new_n500), .B2(G200), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n308), .B2(new_n500), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n444), .A2(new_n492), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n412), .A2(KEYINPUT76), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n413), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n209), .B(G45), .C1(new_n276), .C2(KEYINPUT5), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n273), .A2(G41), .ZN(new_n521));
  OAI211_X1 g0321(.A(G264), .B(new_n269), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT85), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT85), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n295), .A2(new_n524), .A3(G264), .A4(new_n269), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n282), .A2(new_n284), .A3(G250), .A4(new_n288), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n282), .A2(new_n284), .A3(G257), .A4(G1698), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G294), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n292), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n526), .A2(new_n280), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n369), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n523), .A2(new_n525), .B1(new_n530), .B2(new_n292), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(new_n440), .A3(new_n280), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n282), .A2(new_n284), .A3(new_n210), .A4(G87), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT22), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n340), .A2(KEYINPUT22), .A3(new_n210), .A4(G87), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n210), .A2(KEYINPUT23), .A3(G107), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G116), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT23), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n541), .A2(KEYINPUT83), .B1(new_n544), .B2(new_n210), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n206), .A3(G20), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT83), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n546), .A2(new_n547), .B1(KEYINPUT23), .B2(G107), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n539), .A2(new_n540), .A3(new_n545), .A4(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT24), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n330), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI22_X1  g0351(.A1(new_n541), .A2(KEYINPUT83), .B1(new_n543), .B2(new_n206), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n553));
  OAI22_X1  g0353(.A1(new_n546), .A2(new_n547), .B1(new_n553), .B2(G20), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n555), .A2(KEYINPUT24), .A3(new_n539), .A4(new_n540), .ZN(new_n556));
  OR3_X1    g0356(.A1(new_n247), .A2(KEYINPUT25), .A3(G107), .ZN(new_n557));
  OAI21_X1  g0357(.A(KEYINPUT25), .B1(new_n247), .B2(G107), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n557), .B(new_n558), .C1(new_n206), .C2(new_n253), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT84), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n253), .A2(new_n206), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT84), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n561), .A2(new_n562), .A3(new_n557), .A4(new_n558), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n551), .A2(new_n556), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(KEYINPUT86), .B1(new_n536), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n549), .A2(new_n550), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n566), .A2(new_n556), .A3(new_n258), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n560), .A2(new_n563), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT86), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(new_n535), .A4(new_n533), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n532), .A2(G200), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n564), .B(new_n572), .C1(new_n308), .C2(new_n532), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n565), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT87), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT87), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n565), .A2(new_n573), .A3(new_n571), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n508), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(new_n247), .ZN(new_n580));
  INV_X1    g0380(.A(G87), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n253), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(G87), .A2(G107), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n256), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT19), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n210), .B1(new_n448), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n340), .A2(new_n210), .A3(G68), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n585), .B1(new_n256), .B2(new_n427), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI211_X1 g0390(.A(new_n580), .B(new_n582), .C1(new_n590), .C2(new_n258), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n282), .A2(new_n284), .A3(G244), .A4(G1698), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n282), .A2(new_n284), .A3(G238), .A4(new_n288), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n593), .A3(new_n542), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n292), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n269), .A2(G274), .A3(new_n271), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT80), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n269), .A2(KEYINPUT80), .A3(G274), .A4(new_n271), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n269), .B(G250), .C1(G1), .C2(new_n270), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n595), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G200), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n591), .B(new_n603), .C1(new_n308), .C2(new_n602), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n590), .A2(new_n258), .ZN(new_n605));
  INV_X1    g0405(.A(new_n580), .ZN(new_n606));
  OR2_X1    g0406(.A1(new_n253), .A2(new_n508), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n602), .A2(new_n369), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n608), .B(new_n609), .C1(G179), .C2(new_n602), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n206), .A2(KEYINPUT6), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n256), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(G97), .A2(G107), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT6), .B1(new_n207), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(G20), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n336), .A2(G77), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n206), .B1(new_n351), .B2(new_n353), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n258), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n248), .A2(new_n205), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n253), .B2(new_n205), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n282), .A2(new_n284), .A3(G244), .A4(new_n288), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT4), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n340), .A2(KEYINPUT4), .A3(G244), .A4(new_n288), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n340), .A2(G250), .A3(G1698), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n627), .A2(new_n628), .A3(new_n255), .A4(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n292), .ZN(new_n631));
  OAI211_X1 g0431(.A(G257), .B(new_n269), .C1(new_n520), .C2(new_n521), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n274), .A2(new_n277), .A3(new_n278), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n632), .B1(new_n633), .B2(new_n596), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n369), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n634), .B1(new_n630), .B2(new_n292), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n440), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n624), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n636), .A2(G200), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n352), .A2(new_n379), .B1(new_n348), .B2(new_n350), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n617), .B(new_n616), .C1(new_n642), .C2(new_n206), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n622), .B1(new_n643), .B2(new_n258), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n638), .A2(G190), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n641), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n640), .A2(new_n646), .A3(KEYINPUT79), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n611), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(KEYINPUT79), .B1(new_n640), .B2(new_n646), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AND4_X1   g0450(.A1(new_n315), .A2(new_n519), .A3(new_n578), .A4(new_n650), .ZN(G372));
  NAND2_X1  g0451(.A1(new_n487), .A2(new_n491), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n477), .B2(new_n512), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n404), .A2(new_n410), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n372), .A2(new_n392), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT89), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n437), .A2(new_n438), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n655), .A2(KEYINPUT89), .A3(new_n656), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n659), .A2(new_n660), .B1(new_n442), .B2(new_n441), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n640), .A2(new_n646), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(new_n573), .A3(new_n611), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n569), .A2(new_n535), .A3(new_n533), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT88), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n664), .B(new_n665), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n300), .A2(new_n302), .A3(new_n306), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n663), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n604), .A2(new_n610), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n669), .B1(new_n670), .B2(new_n640), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n670), .A2(new_n669), .A3(new_n640), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n610), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n661), .B1(new_n518), .B2(new_n675), .ZN(G369));
  NAND2_X1  g0476(.A1(new_n312), .A2(new_n302), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G213), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n267), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n677), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT90), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n685), .B1(new_n311), .B2(new_n314), .ZN(new_n688));
  OAI21_X1  g0488(.A(G330), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n564), .A2(new_n684), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n578), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n664), .A2(new_n684), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n693), .A2(KEYINPUT91), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT91), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n691), .B1(new_n575), .B2(new_n577), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n697), .B1(new_n698), .B2(new_n694), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n690), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n666), .A2(new_n683), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n677), .A2(new_n684), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n702), .B1(new_n700), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n701), .A2(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n213), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n584), .A2(G116), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n217), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n565), .A2(new_n571), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT95), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(new_n667), .A3(new_n716), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n662), .A2(new_n573), .A3(new_n611), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT95), .B1(new_n677), .B2(new_n714), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n610), .ZN(new_n721));
  INV_X1    g0521(.A(new_n673), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(new_n671), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n683), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT29), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n684), .B1(new_n668), .B2(new_n674), .ZN(new_n726));
  XOR2_X1   g0526(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n578), .A2(new_n315), .A3(new_n650), .A4(new_n684), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n602), .A2(new_n440), .A3(new_n297), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n526), .A2(new_n280), .A3(new_n531), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n526), .A2(new_n531), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n733), .A2(new_n602), .A3(new_n304), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  AOI211_X1 g0535(.A(new_n735), .B(new_n634), .C1(new_n292), .C2(new_n630), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n732), .A2(new_n636), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n595), .A2(new_n600), .A3(new_n601), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n738), .A2(new_n305), .A3(new_n638), .A4(new_n534), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n735), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n684), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(KEYINPUT92), .B1(new_n741), .B2(KEYINPUT31), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT93), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n734), .A2(new_n736), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n297), .A2(new_n440), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n745), .A2(new_n636), .A3(new_n532), .A4(new_n602), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n740), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n683), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT31), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n743), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AOI211_X1 g0550(.A(KEYINPUT93), .B(KEYINPUT31), .C1(new_n747), .C2(new_n683), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n742), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(KEYINPUT93), .B1(new_n741), .B2(KEYINPUT31), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT92), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(new_n748), .B2(new_n749), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n748), .A2(new_n743), .A3(new_n749), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n753), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n729), .A2(new_n752), .A3(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n725), .A2(new_n728), .B1(G330), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n713), .B1(new_n759), .B2(G1), .ZN(G364));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n687), .A2(new_n688), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n219), .B1(G20), .B2(new_n369), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n210), .A2(G179), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n768), .A2(G190), .A3(G200), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n581), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G190), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G159), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n210), .A2(new_n440), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G200), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G190), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n771), .B1(new_n775), .B2(KEYINPUT32), .C1(new_n779), .C2(new_n346), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n775), .A2(KEYINPUT32), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n768), .A2(new_n308), .A3(G200), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n781), .B1(new_n206), .B2(new_n782), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n308), .A2(G179), .A3(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n210), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G97), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n777), .A2(new_n308), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n787), .B1(new_n789), .B2(new_n202), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n776), .A2(new_n772), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n776), .A2(G190), .A3(new_n399), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n340), .B1(new_n791), .B2(new_n461), .C1(new_n324), .C2(new_n792), .ZN(new_n793));
  OR4_X1    g0593(.A1(new_n780), .A2(new_n783), .A3(new_n790), .A4(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G322), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(G311), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n285), .B1(new_n791), .B2(new_n797), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n796), .B(new_n798), .C1(G329), .C2(new_n774), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n788), .A2(G326), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT33), .B(G317), .ZN(new_n801));
  INV_X1    g0601(.A(new_n769), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n778), .A2(new_n801), .B1(new_n802), .B2(G303), .ZN(new_n803));
  INV_X1    g0603(.A(new_n782), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n786), .A2(G294), .B1(new_n804), .B2(G283), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n799), .A2(new_n800), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n767), .B1(new_n794), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G13), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(G20), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n209), .B1(new_n809), .B2(G45), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n708), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n213), .A2(new_n340), .ZN(new_n813));
  INV_X1    g0613(.A(G355), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n813), .A2(new_n814), .B1(G116), .B2(new_n213), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n707), .A2(new_n340), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(new_n270), .B2(new_n218), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n242), .A2(new_n270), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n815), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n763), .A2(new_n766), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n812), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  OR3_X1    g0623(.A1(new_n765), .A2(new_n807), .A3(new_n823), .ZN(new_n824));
  OR3_X1    g0624(.A1(new_n687), .A2(G330), .A3(new_n688), .ZN(new_n825));
  INV_X1    g0625(.A(new_n812), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n825), .A2(new_n689), .A3(new_n826), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G396));
  NAND2_X1  g0629(.A1(new_n511), .A2(new_n683), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n512), .A2(new_n514), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n512), .B2(new_n830), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n726), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n684), .B(new_n832), .C1(new_n668), .C2(new_n674), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n758), .A2(G330), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n812), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n837), .B2(new_n836), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n766), .A2(new_n761), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n826), .B1(new_n461), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n791), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n788), .A2(G303), .B1(new_n842), .B2(G116), .ZN(new_n843));
  INV_X1    g0643(.A(G283), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n844), .B2(new_n779), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT96), .ZN(new_n846));
  INV_X1    g0646(.A(G294), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n285), .B1(new_n773), .B2(new_n797), .C1(new_n792), .C2(new_n847), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n787), .B1(new_n581), .B2(new_n782), .C1(new_n206), .C2(new_n769), .ZN(new_n849));
  OR3_X1    g0649(.A1(new_n846), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  OR2_X1    g0650(.A1(new_n850), .A2(KEYINPUT97), .ZN(new_n851));
  INV_X1    g0651(.A(new_n792), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n852), .A2(G143), .B1(new_n842), .B2(G159), .ZN(new_n853));
  INV_X1    g0653(.A(G150), .ZN(new_n854));
  INV_X1    g0654(.A(G137), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n853), .B1(new_n779), .B2(new_n854), .C1(new_n855), .C2(new_n789), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT34), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n804), .A2(G68), .ZN(new_n859));
  INV_X1    g0659(.A(G132), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n859), .B(new_n340), .C1(new_n860), .C2(new_n773), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n785), .A2(new_n324), .B1(new_n769), .B2(new_n202), .ZN(new_n862));
  NOR3_X1   g0662(.A1(new_n858), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n857), .B2(new_n856), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n850), .A2(KEYINPUT97), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n851), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n841), .B1(new_n762), .B2(new_n832), .C1(new_n866), .C2(new_n767), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n839), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(G384));
  NOR2_X1   g0669(.A1(new_n809), .A2(new_n209), .ZN(new_n870));
  INV_X1    g0670(.A(G330), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n343), .A2(KEYINPUT16), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n329), .B1(new_n872), .B2(new_n344), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n405), .B1(new_n873), .B2(new_n681), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n371), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT37), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n388), .A2(new_n391), .ZN(new_n877));
  INV_X1    g0677(.A(new_n681), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n388), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT37), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n877), .A2(new_n879), .A3(new_n880), .A4(new_n405), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  OR2_X1    g0682(.A1(new_n873), .A2(new_n681), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n882), .B1(new_n411), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(KEYINPUT38), .B(new_n882), .C1(new_n411), .C2(new_n883), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n489), .A2(new_n490), .A3(new_n683), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n492), .A2(new_n890), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n477), .B(new_n889), .C1(new_n487), .C2(new_n491), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n832), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n748), .B(KEYINPUT31), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n893), .B1(new_n729), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n888), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT40), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n405), .B1(new_n356), .B2(new_n371), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n356), .A2(new_n681), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT37), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n900), .A2(new_n881), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n407), .A2(new_n408), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n879), .B1(new_n656), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n885), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n897), .B1(new_n904), .B2(new_n887), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n896), .A2(new_n897), .B1(new_n895), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n518), .B1(new_n729), .B2(new_n894), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n871), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n907), .B2(new_n906), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT100), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n891), .A2(new_n892), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n512), .A2(new_n683), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n912), .B1(new_n835), .B2(new_n914), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n915), .A2(new_n888), .B1(new_n393), .B2(new_n681), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n652), .A2(new_n683), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT99), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT39), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n904), .A2(new_n887), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n904), .A2(new_n887), .A3(new_n919), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT99), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n919), .B1(new_n886), .B2(new_n887), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n917), .B(new_n920), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n916), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n519), .A2(new_n725), .A3(new_n728), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n926), .A2(new_n661), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n925), .B(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n870), .B1(new_n911), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n911), .B2(new_n928), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n613), .A2(new_n615), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT98), .Z(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT35), .ZN(new_n934));
  OAI211_X1 g0734(.A(G116), .B(new_n220), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n934), .B2(new_n933), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT36), .Z(new_n937));
  NOR3_X1   g0737(.A1(new_n217), .A2(new_n461), .A3(new_n331), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n346), .A2(G50), .ZN(new_n939));
  OAI211_X1 g0739(.A(G1), .B(new_n808), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n930), .A2(new_n937), .A3(new_n940), .ZN(G367));
  AND2_X1   g0741(.A1(new_n816), .A2(new_n238), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n821), .B1(new_n213), .B2(new_n508), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n769), .A2(new_n249), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n779), .A2(new_n847), .B1(KEYINPUT46), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(KEYINPUT46), .B2(new_n944), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(KEYINPUT106), .ZN(new_n948));
  INV_X1    g0748(.A(new_n256), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n786), .A2(G107), .B1(new_n804), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n797), .B2(new_n789), .ZN(new_n951));
  INV_X1    g0751(.A(G317), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n285), .B1(new_n773), .B2(new_n952), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n792), .A2(new_n286), .B1(new_n791), .B2(new_n844), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT106), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n955), .B1(new_n946), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n785), .A2(new_n346), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(G143), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n959), .B1(new_n792), .B2(new_n854), .C1(new_n960), .C2(new_n789), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT107), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n285), .B1(new_n804), .B2(G77), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT108), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(KEYINPUT108), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n802), .A2(G58), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n791), .A2(new_n202), .B1(new_n773), .B2(new_n855), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(G159), .B2(new_n778), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n964), .A2(new_n965), .A3(new_n966), .A4(new_n968), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n948), .A2(new_n957), .B1(new_n962), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT47), .Z(new_n971));
  OAI221_X1 g0771(.A(new_n812), .B1(new_n942), .B2(new_n943), .C1(new_n971), .C2(new_n767), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT109), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n591), .A2(new_n684), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT101), .Z(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(new_n610), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT102), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n611), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n977), .B2(new_n976), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n763), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n973), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n662), .B1(new_n644), .B2(new_n684), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n984), .A2(new_n715), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n683), .B1(new_n985), .B2(new_n640), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n703), .B1(new_n696), .B2(new_n699), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n640), .A2(new_n684), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n984), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n986), .B1(new_n991), .B2(KEYINPUT42), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(KEYINPUT42), .B2(new_n991), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT43), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n993), .B1(new_n994), .B2(new_n980), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n980), .A2(new_n994), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n993), .A2(new_n994), .A3(new_n980), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n701), .A2(new_n989), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n1000), .A2(KEYINPUT103), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1000), .B(KEYINPUT103), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n997), .A2(new_n998), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n810), .B(KEYINPUT105), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(KEYINPUT91), .B1(new_n693), .B2(new_n695), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n698), .A2(new_n697), .A3(new_n694), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n704), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n702), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(KEYINPUT44), .B1(new_n1012), .B2(new_n989), .ZN(new_n1013));
  OAI211_X1 g0813(.A(KEYINPUT44), .B(new_n989), .C1(new_n987), .C2(new_n702), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(KEYINPUT45), .B1(new_n705), .B2(new_n990), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT45), .ZN(new_n1017));
  NOR4_X1   g0817(.A1(new_n987), .A2(new_n1017), .A3(new_n702), .A4(new_n989), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n1013), .A2(new_n1015), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n701), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n689), .B(KEYINPUT104), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n696), .A2(new_n699), .A3(new_n703), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1010), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n689), .A2(KEYINPUT104), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1026), .A2(new_n1010), .A3(new_n1023), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1025), .A2(new_n759), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1018), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1017), .B1(new_n1012), .B2(new_n989), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT44), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n705), .B2(new_n990), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n1014), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1032), .A2(new_n1035), .A3(new_n701), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1021), .A2(new_n1029), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n759), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n708), .B(KEYINPUT41), .Z(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1007), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n983), .B1(new_n1005), .B2(new_n1041), .ZN(G387));
  AND2_X1   g0842(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1043), .A2(new_n759), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1028), .A2(new_n708), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1043), .A2(new_n1007), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n813), .A2(new_n710), .B1(G107), .B2(new_n213), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n710), .B(KEYINPUT110), .Z(new_n1049));
  OAI21_X1  g0849(.A(new_n270), .B1(new_n346), .B2(new_n461), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n321), .A2(G50), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT50), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1049), .B(new_n1053), .C1(new_n1052), .C2(new_n1051), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n817), .B1(new_n235), .B2(G45), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1048), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n812), .B1(new_n1056), .B2(new_n822), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n792), .A2(new_n202), .B1(new_n791), .B2(new_n346), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n285), .B(new_n1058), .C1(G150), .C2(new_n774), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n786), .A2(new_n579), .B1(new_n804), .B2(G97), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n788), .A2(G159), .B1(new_n802), .B2(G77), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n778), .A2(new_n325), .A3(new_n323), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n785), .A2(new_n844), .B1(new_n769), .B2(new_n847), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n852), .A2(G317), .B1(new_n842), .B2(G303), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n779), .B2(new_n797), .C1(new_n795), .C2(new_n789), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT48), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1064), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n1067), .B2(new_n1066), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT49), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n340), .B1(new_n774), .B2(G326), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n249), .B2(new_n782), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT111), .Z(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1063), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1057), .B1(new_n1076), .B2(new_n766), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n700), .B2(new_n764), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1047), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1046), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(G393));
  INV_X1    g0881(.A(KEYINPUT114), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT112), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1021), .A2(new_n1083), .A3(new_n1036), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1019), .A2(KEYINPUT112), .A3(new_n1020), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n1084), .A2(new_n1028), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1037), .A2(new_n708), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1082), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1087), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1084), .A2(new_n1028), .A3(new_n1085), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1089), .A2(KEYINPUT114), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n989), .A2(new_n763), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n285), .B1(new_n773), .B2(new_n795), .C1(new_n206), .C2(new_n782), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G283), .B2(new_n802), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT113), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n789), .A2(new_n952), .B1(new_n797), .B2(new_n792), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT52), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n785), .A2(new_n249), .B1(new_n791), .B2(new_n847), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(G303), .B2(new_n778), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1096), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n789), .A2(new_n854), .B1(new_n333), .B2(new_n792), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT51), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n340), .B1(new_n773), .B2(new_n960), .C1(new_n321), .C2(new_n791), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n778), .A2(G50), .B1(new_n804), .B2(G87), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n785), .A2(new_n461), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G68), .B2(new_n802), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1103), .A2(new_n1105), .A3(new_n1106), .A4(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n767), .B1(new_n1101), .B2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n817), .A2(new_n245), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n822), .B(new_n1111), .C1(new_n707), .C2(new_n949), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1110), .A2(new_n826), .A3(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1092), .A2(new_n1007), .B1(new_n1093), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1088), .A2(new_n1091), .A3(new_n1114), .ZN(G390));
  INV_X1    g0915(.A(new_n912), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n683), .B(new_n833), .C1(new_n720), .C2(new_n723), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1116), .B1(new_n1117), .B2(new_n913), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n917), .B1(new_n904), .B2(new_n887), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n758), .A2(G330), .A3(new_n832), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1121), .A2(new_n912), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n920), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n921), .A2(KEYINPUT99), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n888), .A2(KEYINPUT39), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n915), .A2(new_n917), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1120), .B(new_n1122), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n917), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n666), .A2(new_n667), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n718), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n683), .B1(new_n1132), .B2(new_n723), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n913), .B1(new_n1133), .B2(new_n832), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1130), .B1(new_n1134), .B2(new_n912), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1129), .A2(new_n1135), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n871), .B1(new_n729), .B2(new_n894), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n893), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1128), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1140), .A2(new_n1006), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n779), .A2(new_n855), .B1(new_n333), .B2(new_n785), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G128), .B2(new_n788), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n769), .A2(new_n854), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT53), .ZN(new_n1145));
  INV_X1    g0945(.A(G125), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n792), .A2(new_n860), .B1(new_n773), .B2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(KEYINPUT54), .B(G143), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1147), .B1(new_n842), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1143), .A2(new_n1145), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n340), .B1(new_n782), .B2(new_n202), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT116), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n792), .A2(new_n249), .B1(new_n773), .B2(new_n847), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n340), .B(new_n1154), .C1(new_n949), .C2(new_n842), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1155), .A2(new_n771), .A3(new_n859), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1107), .B1(G283), .B2(new_n788), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n206), .B2(new_n779), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n1151), .A2(new_n1153), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n766), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n826), .B1(new_n326), .B2(new_n840), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n1129), .B2(new_n761), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1141), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n519), .A2(new_n1137), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n926), .A2(new_n661), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1121), .A2(new_n912), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(KEYINPUT115), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT115), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1121), .A2(new_n1170), .A3(new_n912), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1169), .A2(new_n1139), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1134), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n913), .B1(new_n724), .B2(new_n832), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n1121), .B2(new_n912), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1116), .B1(new_n1137), .B2(new_n832), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1167), .B1(new_n1174), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1128), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1129), .A2(new_n1135), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1139), .B1(new_n1182), .B2(new_n1120), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n708), .B1(new_n1180), .B2(new_n1184), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1168), .A2(KEYINPUT115), .B1(new_n1138), .B2(new_n1137), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1134), .B1(new_n1186), .B2(new_n1171), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1166), .B1(new_n1187), .B2(new_n1178), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1188), .A2(new_n1140), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1164), .B1(new_n1185), .B2(new_n1189), .ZN(G378));
  AOI21_X1  g0990(.A(new_n826), .B1(new_n202), .B2(new_n840), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n778), .A2(G97), .B1(new_n842), .B2(new_n579), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT117), .Z(new_n1193));
  NAND2_X1  g0993(.A1(new_n285), .A2(new_n276), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n773), .A2(new_n844), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1194), .B(new_n1195), .C1(G107), .C2(new_n852), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n958), .B1(G77), .B2(new_n802), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n788), .A2(G116), .B1(new_n804), .B2(G58), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1193), .A2(new_n1196), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT58), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1194), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT118), .Z(new_n1204));
  NOR2_X1   g1004(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n1146), .A2(new_n789), .B1(new_n779), .B2(new_n860), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n852), .A2(G128), .B1(new_n842), .B2(G137), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n769), .B2(new_n1148), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1206), .B(new_n1208), .C1(G150), .C2(new_n786), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n804), .A2(G159), .ZN(new_n1212));
  AOI211_X1 g1012(.A(G33), .B(G41), .C1(new_n774), .C2(G124), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT59), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1214), .B1(new_n1215), .B2(new_n1209), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1204), .A2(new_n1205), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n442), .A2(new_n878), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n444), .B(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1219), .B(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1191), .B1(new_n767), .B2(new_n1217), .C1(new_n1222), .C2(new_n762), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT119), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n896), .A2(new_n897), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n905), .A2(new_n895), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1226), .A2(G330), .A3(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1228), .A2(new_n1221), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1222), .B1(new_n906), .B2(G330), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1225), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n925), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1228), .A2(new_n1221), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n906), .A2(G330), .A3(new_n1222), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n916), .A2(new_n924), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n1225), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1232), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1224), .B1(new_n1238), .B2(new_n1007), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1178), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1166), .B1(new_n1140), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT57), .B1(new_n1238), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1174), .A2(new_n1179), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1167), .B1(new_n1184), .B2(new_n1243), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1229), .A2(new_n1230), .A3(new_n1236), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n925), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1246));
  OAI21_X1  g1046(.A(KEYINPUT57), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n708), .B1(new_n1244), .B2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1239), .B1(new_n1242), .B2(new_n1248), .ZN(G375));
  OAI22_X1  g1049(.A1(new_n249), .A2(new_n779), .B1(new_n789), .B2(new_n847), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(G97), .B2(new_n802), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n792), .A2(new_n844), .B1(new_n791), .B2(new_n206), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n340), .B(new_n1252), .C1(G303), .C2(new_n774), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n786), .A2(new_n579), .B1(new_n804), .B2(G77), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1251), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT121), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n789), .A2(new_n860), .B1(new_n202), .B2(new_n785), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(G159), .B2(new_n802), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n285), .B1(new_n852), .B2(G137), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(G150), .A2(new_n842), .B1(new_n774), .B2(G128), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n778), .A2(new_n1149), .B1(new_n804), .B2(G58), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1257), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1265), .A2(new_n766), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n826), .B(new_n1266), .C1(new_n346), .C2(new_n840), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(KEYINPUT122), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n912), .A2(new_n761), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(KEYINPUT120), .B1(new_n1240), .B2(new_n1006), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT120), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1273), .B(new_n1007), .C1(new_n1187), .C2(new_n1178), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1271), .B1(new_n1272), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1240), .A2(new_n1167), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(new_n1188), .A3(new_n1040), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(G381));
  NAND2_X1  g1078(.A1(new_n1080), .A2(new_n828), .ZN(new_n1279));
  NOR4_X1   g1079(.A1(new_n1279), .A2(G378), .A3(G381), .A4(G384), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1041), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n982), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  OR2_X1    g1084(.A1(G390), .A2(G375), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT123), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NOR3_X1   g1088(.A1(new_n1284), .A2(new_n1285), .A3(KEYINPUT123), .ZN(new_n1289));
  OR2_X1    g1089(.A1(new_n1288), .A2(new_n1289), .ZN(G407));
  INV_X1    g1090(.A(G378), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n682), .ZN(new_n1292));
  OAI221_X1 g1092(.A(G213), .B1(G375), .B2(new_n1292), .C1(new_n1288), .C2(new_n1289), .ZN(G409));
  INV_X1    g1093(.A(KEYINPUT126), .ZN(new_n1294));
  OAI21_X1  g1094(.A(G396), .B1(new_n1046), .B2(new_n1079), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1294), .B1(new_n1279), .B2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(G390), .B2(G387), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT114), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1092), .A2(new_n1007), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1093), .A2(new_n1113), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1298), .A2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1283), .A2(new_n1302), .A3(new_n1091), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1297), .A2(new_n1303), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1279), .A2(new_n1295), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1294), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1304), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1297), .A2(new_n1303), .A3(new_n1306), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1174), .A2(new_n1167), .A3(KEYINPUT60), .A4(new_n1179), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n708), .ZN(new_n1312));
  OAI21_X1  g1112(.A(KEYINPUT60), .B1(new_n1240), .B2(new_n1167), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1312), .B1(new_n1276), .B2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1270), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n868), .B1(new_n1314), .B2(new_n1316), .ZN(new_n1317));
  NOR3_X1   g1117(.A1(new_n1187), .A2(new_n1166), .A3(new_n1178), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1318), .B1(KEYINPUT60), .B2(new_n1188), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1275), .B(G384), .C1(new_n1319), .C2(new_n1312), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n682), .A2(G213), .A3(G2897), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1317), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1321), .B1(new_n1317), .B2(new_n1320), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n682), .A2(G213), .ZN(new_n1325));
  OAI211_X1 g1125(.A(G378), .B(new_n1239), .C1(new_n1242), .C2(new_n1248), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1007), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(new_n1223), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1231), .A2(new_n925), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1236), .B1(new_n1235), .B2(new_n1225), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1241), .B(new_n1040), .C1(new_n1330), .C2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1329), .B1(new_n1332), .B2(KEYINPUT124), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT124), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1238), .A2(new_n1334), .A3(new_n1040), .A4(new_n1241), .ZN(new_n1335));
  AOI21_X1  g1135(.A(G378), .B1(new_n1333), .B2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1325), .B1(new_n1327), .B2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(KEYINPUT61), .B1(new_n1324), .B2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1320), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1313), .A2(new_n1276), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1340), .A2(new_n708), .A3(new_n1311), .ZN(new_n1341));
  AOI21_X1  g1141(.A(G384), .B1(new_n1341), .B2(new_n1275), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1339), .A2(new_n1342), .ZN(new_n1343));
  OAI211_X1 g1143(.A(new_n1325), .B(new_n1343), .C1(new_n1327), .C2(new_n1336), .ZN(new_n1344));
  AND2_X1   g1144(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1344), .B1(KEYINPUT125), .B2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1338), .A2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1332), .A2(KEYINPUT124), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1329), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1348), .A2(new_n1335), .A3(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1350), .A2(new_n1291), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(new_n1326), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT125), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1352), .A2(new_n1353), .A3(new_n1325), .A4(new_n1343), .ZN(new_n1354));
  AOI21_X1  g1154(.A(KEYINPUT62), .B1(new_n1354), .B2(KEYINPUT127), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1310), .B1(new_n1347), .B2(new_n1355), .ZN(new_n1356));
  AND3_X1   g1156(.A1(new_n1297), .A2(new_n1303), .A3(new_n1306), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1306), .B1(new_n1297), .B2(new_n1303), .ZN(new_n1358));
  NOR2_X1   g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1344), .A2(KEYINPUT125), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT63), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1360), .A2(new_n1361), .A3(new_n1354), .ZN(new_n1362));
  OR2_X1    g1162(.A1(new_n1344), .A2(new_n1361), .ZN(new_n1363));
  NAND4_X1  g1163(.A1(new_n1359), .A2(new_n1362), .A3(new_n1338), .A4(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1356), .A2(new_n1364), .ZN(G405));
  NAND2_X1  g1165(.A1(G375), .A2(new_n1291), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1366), .A2(new_n1326), .ZN(new_n1367));
  XNOR2_X1  g1167(.A(new_n1367), .B(new_n1343), .ZN(new_n1368));
  XNOR2_X1  g1168(.A(new_n1310), .B(new_n1368), .ZN(G402));
endmodule


