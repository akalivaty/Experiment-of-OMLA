

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(n1007), .A2(n606), .ZN(n616) );
  INV_X1 U551 ( .A(KEYINPUT97), .ZN(n658) );
  NOR2_X1 U552 ( .A1(G651), .A2(n564), .ZN(n786) );
  XOR2_X1 U553 ( .A(n518), .B(KEYINPUT17), .Z(n882) );
  XNOR2_X1 U554 ( .A(n754), .B(KEYINPUT40), .ZN(n755) );
  OR2_X1 U555 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U556 ( .A(n756), .B(n755), .ZN(G329) );
  XNOR2_X1 U557 ( .A(n527), .B(KEYINPUT87), .ZN(G164) );
  NOR2_X1 U558 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  NAND2_X1 U559 ( .A1(G138), .A2(n882), .ZN(n520) );
  INV_X1 U560 ( .A(G2105), .ZN(n522) );
  NOR2_X1 U561 ( .A1(G2104), .A2(n522), .ZN(n886) );
  NAND2_X1 U562 ( .A1(G126), .A2(n886), .ZN(n519) );
  NAND2_X1 U563 ( .A1(n520), .A2(n519), .ZN(n526) );
  NAND2_X1 U564 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  XNOR2_X1 U565 ( .A(n521), .B(KEYINPUT65), .ZN(n885) );
  NAND2_X1 U566 ( .A1(G114), .A2(n885), .ZN(n524) );
  AND2_X1 U567 ( .A1(n522), .A2(G2104), .ZN(n881) );
  NAND2_X1 U568 ( .A1(G102), .A2(n881), .ZN(n523) );
  NAND2_X1 U569 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U570 ( .A1(n885), .A2(G113), .ZN(n530) );
  NAND2_X1 U571 ( .A1(G101), .A2(n881), .ZN(n528) );
  XOR2_X1 U572 ( .A(KEYINPUT23), .B(n528), .Z(n529) );
  NAND2_X1 U573 ( .A1(n530), .A2(n529), .ZN(n534) );
  NAND2_X1 U574 ( .A1(G125), .A2(n886), .ZN(n532) );
  NAND2_X1 U575 ( .A1(G137), .A2(n882), .ZN(n531) );
  NAND2_X1 U576 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U577 ( .A1(n534), .A2(n533), .ZN(G160) );
  XOR2_X1 U578 ( .A(KEYINPUT0), .B(G543), .Z(n564) );
  NAND2_X1 U579 ( .A1(n786), .A2(G52), .ZN(n538) );
  INV_X1 U580 ( .A(G651), .ZN(n539) );
  NOR2_X1 U581 ( .A1(G543), .A2(n539), .ZN(n535) );
  XOR2_X1 U582 ( .A(KEYINPUT66), .B(n535), .Z(n536) );
  XNOR2_X1 U583 ( .A(KEYINPUT1), .B(n536), .ZN(n783) );
  NAND2_X1 U584 ( .A1(G64), .A2(n783), .ZN(n537) );
  NAND2_X1 U585 ( .A1(n538), .A2(n537), .ZN(n544) );
  NOR2_X1 U586 ( .A1(G651), .A2(G543), .ZN(n785) );
  NAND2_X1 U587 ( .A1(G90), .A2(n785), .ZN(n541) );
  NOR2_X1 U588 ( .A1(n564), .A2(n539), .ZN(n789) );
  NAND2_X1 U589 ( .A1(G77), .A2(n789), .ZN(n540) );
  NAND2_X1 U590 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U591 ( .A(KEYINPUT9), .B(n542), .Z(n543) );
  NOR2_X1 U592 ( .A1(n544), .A2(n543), .ZN(G171) );
  NAND2_X1 U593 ( .A1(n785), .A2(G89), .ZN(n545) );
  XNOR2_X1 U594 ( .A(KEYINPUT4), .B(n545), .ZN(n548) );
  NAND2_X1 U595 ( .A1(n789), .A2(G76), .ZN(n546) );
  XOR2_X1 U596 ( .A(KEYINPUT69), .B(n546), .Z(n547) );
  NAND2_X1 U597 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U598 ( .A(n549), .B(KEYINPUT5), .ZN(n554) );
  NAND2_X1 U599 ( .A1(n786), .A2(G51), .ZN(n551) );
  NAND2_X1 U600 ( .A1(G63), .A2(n783), .ZN(n550) );
  NAND2_X1 U601 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U602 ( .A(KEYINPUT6), .B(n552), .Z(n553) );
  NAND2_X1 U603 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U604 ( .A(n555), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U605 ( .A1(n786), .A2(G50), .ZN(n556) );
  XOR2_X1 U606 ( .A(KEYINPUT81), .B(n556), .Z(n558) );
  NAND2_X1 U607 ( .A1(G62), .A2(n783), .ZN(n557) );
  NAND2_X1 U608 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U609 ( .A(KEYINPUT82), .B(n559), .ZN(n563) );
  NAND2_X1 U610 ( .A1(G88), .A2(n785), .ZN(n561) );
  NAND2_X1 U611 ( .A1(G75), .A2(n789), .ZN(n560) );
  NAND2_X1 U612 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U613 ( .A1(n563), .A2(n562), .ZN(G166) );
  XOR2_X1 U614 ( .A(KEYINPUT88), .B(G166), .Z(G303) );
  XOR2_X1 U615 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U616 ( .A1(G49), .A2(n786), .ZN(n566) );
  NAND2_X1 U617 ( .A1(G87), .A2(n564), .ZN(n565) );
  NAND2_X1 U618 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U619 ( .A1(n783), .A2(n567), .ZN(n570) );
  NAND2_X1 U620 ( .A1(G74), .A2(G651), .ZN(n568) );
  XOR2_X1 U621 ( .A(KEYINPUT77), .B(n568), .Z(n569) );
  NAND2_X1 U622 ( .A1(n570), .A2(n569), .ZN(G288) );
  NAND2_X1 U623 ( .A1(G48), .A2(n786), .ZN(n579) );
  NAND2_X1 U624 ( .A1(n783), .A2(G61), .ZN(n571) );
  XNOR2_X1 U625 ( .A(n571), .B(KEYINPUT78), .ZN(n574) );
  NAND2_X1 U626 ( .A1(G73), .A2(n789), .ZN(n572) );
  XNOR2_X1 U627 ( .A(n572), .B(KEYINPUT2), .ZN(n573) );
  NAND2_X1 U628 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U629 ( .A1(G86), .A2(n785), .ZN(n575) );
  XNOR2_X1 U630 ( .A(KEYINPUT79), .B(n575), .ZN(n576) );
  NOR2_X1 U631 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U632 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U633 ( .A(n580), .B(KEYINPUT80), .ZN(G305) );
  NAND2_X1 U634 ( .A1(G85), .A2(n785), .ZN(n582) );
  NAND2_X1 U635 ( .A1(G72), .A2(n789), .ZN(n581) );
  NAND2_X1 U636 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U637 ( .A1(n786), .A2(G47), .ZN(n584) );
  NAND2_X1 U638 ( .A1(G60), .A2(n783), .ZN(n583) );
  NAND2_X1 U639 ( .A1(n584), .A2(n583), .ZN(n585) );
  OR2_X1 U640 ( .A1(n586), .A2(n585), .ZN(G290) );
  NAND2_X1 U641 ( .A1(n785), .A2(G81), .ZN(n587) );
  XNOR2_X1 U642 ( .A(n587), .B(KEYINPUT12), .ZN(n589) );
  NAND2_X1 U643 ( .A1(G68), .A2(n789), .ZN(n588) );
  NAND2_X1 U644 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U645 ( .A(KEYINPUT13), .B(n590), .Z(n594) );
  NAND2_X1 U646 ( .A1(n783), .A2(G56), .ZN(n591) );
  XNOR2_X1 U647 ( .A(n591), .B(KEYINPUT14), .ZN(n592) );
  XNOR2_X1 U648 ( .A(n592), .B(KEYINPUT67), .ZN(n593) );
  NOR2_X1 U649 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U650 ( .A1(n786), .A2(G43), .ZN(n595) );
  NAND2_X1 U651 ( .A1(n596), .A2(n595), .ZN(n1007) );
  INV_X1 U652 ( .A(G164), .ZN(n599) );
  NAND2_X1 U653 ( .A1(G160), .A2(G40), .ZN(n706) );
  INV_X1 U654 ( .A(n706), .ZN(n597) );
  INV_X1 U655 ( .A(G1384), .ZN(n705) );
  AND2_X1 U656 ( .A1(n597), .A2(n705), .ZN(n598) );
  NAND2_X1 U657 ( .A1(n599), .A2(n598), .ZN(n601) );
  INV_X1 U658 ( .A(KEYINPUT64), .ZN(n600) );
  XNOR2_X2 U659 ( .A(n601), .B(n600), .ZN(n642) );
  NAND2_X1 U660 ( .A1(G1996), .A2(n642), .ZN(n602) );
  XNOR2_X1 U661 ( .A(n602), .B(KEYINPUT26), .ZN(n604) );
  INV_X1 U662 ( .A(n642), .ZN(n663) );
  NAND2_X1 U663 ( .A1(G1341), .A2(n663), .ZN(n603) );
  NAND2_X1 U664 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U665 ( .A(n605), .B(KEYINPUT94), .ZN(n606) );
  NAND2_X1 U666 ( .A1(n783), .A2(G66), .ZN(n613) );
  NAND2_X1 U667 ( .A1(G92), .A2(n785), .ZN(n608) );
  NAND2_X1 U668 ( .A1(G79), .A2(n789), .ZN(n607) );
  NAND2_X1 U669 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U670 ( .A1(n786), .A2(G54), .ZN(n609) );
  XOR2_X1 U671 ( .A(KEYINPUT68), .B(n609), .Z(n610) );
  NOR2_X1 U672 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U673 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U674 ( .A(n614), .B(KEYINPUT15), .ZN(n1006) );
  NOR2_X1 U675 ( .A1(n616), .A2(n1006), .ZN(n615) );
  XNOR2_X1 U676 ( .A(n615), .B(KEYINPUT95), .ZN(n622) );
  NAND2_X1 U677 ( .A1(n616), .A2(n1006), .ZN(n620) );
  NOR2_X1 U678 ( .A1(G2067), .A2(n663), .ZN(n618) );
  NOR2_X1 U679 ( .A1(G1348), .A2(n642), .ZN(n617) );
  NOR2_X1 U680 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U681 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U682 ( .A1(n622), .A2(n621), .ZN(n634) );
  NAND2_X1 U683 ( .A1(n786), .A2(G53), .ZN(n624) );
  NAND2_X1 U684 ( .A1(G65), .A2(n783), .ZN(n623) );
  NAND2_X1 U685 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U686 ( .A1(G91), .A2(n785), .ZN(n626) );
  NAND2_X1 U687 ( .A1(G78), .A2(n789), .ZN(n625) );
  NAND2_X1 U688 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U689 ( .A1(n628), .A2(n627), .ZN(n798) );
  XOR2_X1 U690 ( .A(KEYINPUT27), .B(KEYINPUT93), .Z(n630) );
  NAND2_X1 U691 ( .A1(G2072), .A2(n642), .ZN(n629) );
  XNOR2_X1 U692 ( .A(n630), .B(n629), .ZN(n632) );
  INV_X1 U693 ( .A(G1956), .ZN(n925) );
  NOR2_X1 U694 ( .A1(n642), .A2(n925), .ZN(n631) );
  NOR2_X1 U695 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U696 ( .A1(n798), .A2(n635), .ZN(n633) );
  NAND2_X1 U697 ( .A1(n634), .A2(n633), .ZN(n638) );
  NOR2_X1 U698 ( .A1(n798), .A2(n635), .ZN(n636) );
  XOR2_X1 U699 ( .A(n636), .B(KEYINPUT28), .Z(n637) );
  NAND2_X1 U700 ( .A1(n638), .A2(n637), .ZN(n640) );
  XOR2_X1 U701 ( .A(KEYINPUT29), .B(KEYINPUT96), .Z(n639) );
  XNOR2_X1 U702 ( .A(n640), .B(n639), .ZN(n646) );
  XNOR2_X1 U703 ( .A(G2078), .B(KEYINPUT25), .ZN(n641) );
  XNOR2_X1 U704 ( .A(n641), .B(KEYINPUT92), .ZN(n947) );
  NAND2_X1 U705 ( .A1(n947), .A2(n642), .ZN(n644) );
  INV_X1 U706 ( .A(G1961), .ZN(n918) );
  NAND2_X1 U707 ( .A1(n663), .A2(n918), .ZN(n643) );
  NAND2_X1 U708 ( .A1(n644), .A2(n643), .ZN(n650) );
  NAND2_X1 U709 ( .A1(n650), .A2(G171), .ZN(n645) );
  NAND2_X1 U710 ( .A1(n646), .A2(n645), .ZN(n655) );
  NOR2_X1 U711 ( .A1(n663), .A2(G2084), .ZN(n660) );
  NAND2_X1 U712 ( .A1(G8), .A2(n663), .ZN(n729) );
  NOR2_X1 U713 ( .A1(G1966), .A2(n729), .ZN(n656) );
  NOR2_X1 U714 ( .A1(n660), .A2(n656), .ZN(n647) );
  NAND2_X1 U715 ( .A1(G8), .A2(n647), .ZN(n648) );
  XNOR2_X1 U716 ( .A(KEYINPUT30), .B(n648), .ZN(n649) );
  NOR2_X1 U717 ( .A1(G168), .A2(n649), .ZN(n652) );
  NOR2_X1 U718 ( .A1(G171), .A2(n650), .ZN(n651) );
  NOR2_X1 U719 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U720 ( .A(KEYINPUT31), .B(n653), .Z(n654) );
  NAND2_X1 U721 ( .A1(n655), .A2(n654), .ZN(n668) );
  INV_X1 U722 ( .A(n668), .ZN(n657) );
  NOR2_X1 U723 ( .A1(n657), .A2(n656), .ZN(n659) );
  XNOR2_X1 U724 ( .A(n659), .B(n658), .ZN(n662) );
  NAND2_X1 U725 ( .A1(G8), .A2(n660), .ZN(n661) );
  NAND2_X1 U726 ( .A1(n662), .A2(n661), .ZN(n674) );
  NOR2_X1 U727 ( .A1(n663), .A2(G2090), .ZN(n664) );
  XNOR2_X1 U728 ( .A(n664), .B(KEYINPUT98), .ZN(n666) );
  NOR2_X1 U729 ( .A1(n729), .A2(G1971), .ZN(n665) );
  NOR2_X1 U730 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U731 ( .A1(n667), .A2(G303), .ZN(n670) );
  NAND2_X1 U732 ( .A1(G286), .A2(n668), .ZN(n669) );
  NAND2_X1 U733 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U734 ( .A1(G8), .A2(n671), .ZN(n672) );
  XNOR2_X1 U735 ( .A(KEYINPUT32), .B(n672), .ZN(n673) );
  NAND2_X1 U736 ( .A1(n674), .A2(n673), .ZN(n725) );
  NOR2_X1 U737 ( .A1(G1976), .A2(G288), .ZN(n681) );
  NOR2_X1 U738 ( .A1(G303), .A2(G1971), .ZN(n675) );
  NOR2_X1 U739 ( .A1(n681), .A2(n675), .ZN(n1016) );
  XOR2_X1 U740 ( .A(n1016), .B(KEYINPUT99), .Z(n676) );
  NAND2_X1 U741 ( .A1(n725), .A2(n676), .ZN(n679) );
  INV_X1 U742 ( .A(n729), .ZN(n677) );
  NAND2_X1 U743 ( .A1(G1976), .A2(G288), .ZN(n1002) );
  AND2_X1 U744 ( .A1(n677), .A2(n1002), .ZN(n678) );
  AND2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U746 ( .A1(KEYINPUT33), .A2(n680), .ZN(n685) );
  NAND2_X1 U747 ( .A1(KEYINPUT33), .A2(n681), .ZN(n682) );
  XNOR2_X1 U748 ( .A(KEYINPUT100), .B(n682), .ZN(n683) );
  NOR2_X1 U749 ( .A1(n729), .A2(n683), .ZN(n684) );
  NOR2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n722) );
  XNOR2_X1 U751 ( .A(G1981), .B(G305), .ZN(n686) );
  XNOR2_X1 U752 ( .A(n686), .B(KEYINPUT101), .ZN(n997) );
  NAND2_X1 U753 ( .A1(G107), .A2(n885), .ZN(n688) );
  NAND2_X1 U754 ( .A1(G95), .A2(n881), .ZN(n687) );
  NAND2_X1 U755 ( .A1(n688), .A2(n687), .ZN(n692) );
  NAND2_X1 U756 ( .A1(G119), .A2(n886), .ZN(n690) );
  NAND2_X1 U757 ( .A1(G131), .A2(n882), .ZN(n689) );
  NAND2_X1 U758 ( .A1(n690), .A2(n689), .ZN(n691) );
  OR2_X1 U759 ( .A1(n692), .A2(n691), .ZN(n863) );
  NAND2_X1 U760 ( .A1(G1991), .A2(n863), .ZN(n703) );
  NAND2_X1 U761 ( .A1(G105), .A2(n881), .ZN(n693) );
  XOR2_X1 U762 ( .A(KEYINPUT38), .B(n693), .Z(n699) );
  NAND2_X1 U763 ( .A1(n885), .A2(G117), .ZN(n694) );
  XNOR2_X1 U764 ( .A(n694), .B(KEYINPUT90), .ZN(n696) );
  NAND2_X1 U765 ( .A1(G129), .A2(n886), .ZN(n695) );
  NAND2_X1 U766 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U767 ( .A(KEYINPUT91), .B(n697), .Z(n698) );
  NOR2_X1 U768 ( .A1(n699), .A2(n698), .ZN(n701) );
  NAND2_X1 U769 ( .A1(n882), .A2(G141), .ZN(n700) );
  NAND2_X1 U770 ( .A1(n701), .A2(n700), .ZN(n877) );
  NAND2_X1 U771 ( .A1(G1996), .A2(n877), .ZN(n702) );
  NAND2_X1 U772 ( .A1(n703), .A2(n702), .ZN(n980) );
  INV_X1 U773 ( .A(n980), .ZN(n704) );
  XOR2_X1 U774 ( .A(G1986), .B(G290), .Z(n1003) );
  NAND2_X1 U775 ( .A1(n704), .A2(n1003), .ZN(n708) );
  AND2_X1 U776 ( .A1(n599), .A2(n705), .ZN(n707) );
  NOR2_X1 U777 ( .A1(n707), .A2(n706), .ZN(n741) );
  NAND2_X1 U778 ( .A1(n708), .A2(n741), .ZN(n719) );
  XNOR2_X1 U779 ( .A(G2067), .B(KEYINPUT37), .ZN(n738) );
  NAND2_X1 U780 ( .A1(G104), .A2(n881), .ZN(n710) );
  NAND2_X1 U781 ( .A1(G140), .A2(n882), .ZN(n709) );
  NAND2_X1 U782 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U783 ( .A(KEYINPUT34), .B(n711), .ZN(n716) );
  NAND2_X1 U784 ( .A1(G116), .A2(n885), .ZN(n713) );
  NAND2_X1 U785 ( .A1(G128), .A2(n886), .ZN(n712) );
  NAND2_X1 U786 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U787 ( .A(n714), .B(KEYINPUT35), .Z(n715) );
  NOR2_X1 U788 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U789 ( .A(KEYINPUT36), .B(n717), .Z(n718) );
  XNOR2_X1 U790 ( .A(KEYINPUT89), .B(n718), .ZN(n862) );
  NOR2_X1 U791 ( .A1(n738), .A2(n862), .ZN(n985) );
  NAND2_X1 U792 ( .A1(n985), .A2(n741), .ZN(n736) );
  NAND2_X1 U793 ( .A1(n719), .A2(n736), .ZN(n748) );
  INV_X1 U794 ( .A(n748), .ZN(n720) );
  AND2_X1 U795 ( .A1(n997), .A2(n720), .ZN(n721) );
  NAND2_X1 U796 ( .A1(n722), .A2(n721), .ZN(n753) );
  NOR2_X1 U797 ( .A1(G2090), .A2(G303), .ZN(n723) );
  NAND2_X1 U798 ( .A1(G8), .A2(n723), .ZN(n724) );
  NAND2_X1 U799 ( .A1(n725), .A2(n724), .ZN(n726) );
  AND2_X1 U800 ( .A1(n726), .A2(n729), .ZN(n746) );
  NOR2_X1 U801 ( .A1(G1981), .A2(G305), .ZN(n727) );
  XOR2_X1 U802 ( .A(n727), .B(KEYINPUT24), .Z(n728) );
  NOR2_X1 U803 ( .A1(n729), .A2(n728), .ZN(n744) );
  NOR2_X1 U804 ( .A1(G1996), .A2(n877), .ZN(n974) );
  NOR2_X1 U805 ( .A1(G1986), .A2(G290), .ZN(n730) );
  NOR2_X1 U806 ( .A1(G1991), .A2(n863), .ZN(n979) );
  NOR2_X1 U807 ( .A1(n730), .A2(n979), .ZN(n731) );
  XNOR2_X1 U808 ( .A(n731), .B(KEYINPUT102), .ZN(n732) );
  NOR2_X1 U809 ( .A1(n980), .A2(n732), .ZN(n733) );
  NOR2_X1 U810 ( .A1(n974), .A2(n733), .ZN(n735) );
  XOR2_X1 U811 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n734) );
  XNOR2_X1 U812 ( .A(n735), .B(n734), .ZN(n737) );
  NAND2_X1 U813 ( .A1(n737), .A2(n736), .ZN(n739) );
  NAND2_X1 U814 ( .A1(n738), .A2(n862), .ZN(n988) );
  NAND2_X1 U815 ( .A1(n739), .A2(n988), .ZN(n740) );
  XNOR2_X1 U816 ( .A(KEYINPUT104), .B(n740), .ZN(n742) );
  NAND2_X1 U817 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U818 ( .A(n743), .B(KEYINPUT105), .ZN(n747) );
  OR2_X1 U819 ( .A1(n744), .A2(n747), .ZN(n745) );
  NOR2_X1 U820 ( .A1(n746), .A2(n745), .ZN(n751) );
  INV_X1 U821 ( .A(n747), .ZN(n749) );
  AND2_X1 U822 ( .A1(n749), .A2(n748), .ZN(n750) );
  OR2_X1 U823 ( .A1(n751), .A2(n750), .ZN(n752) );
  AND2_X1 U824 ( .A1(n753), .A2(n752), .ZN(n756) );
  INV_X1 U825 ( .A(KEYINPUT106), .ZN(n754) );
  AND2_X1 U826 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U827 ( .A(G57), .ZN(G237) );
  INV_X1 U828 ( .A(n798), .ZN(G299) );
  NAND2_X1 U829 ( .A1(G7), .A2(G661), .ZN(n757) );
  XNOR2_X1 U830 ( .A(n757), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U831 ( .A(G223), .ZN(n825) );
  NAND2_X1 U832 ( .A1(n825), .A2(G567), .ZN(n758) );
  XOR2_X1 U833 ( .A(KEYINPUT11), .B(n758), .Z(G234) );
  INV_X1 U834 ( .A(G860), .ZN(n782) );
  OR2_X1 U835 ( .A1(n1007), .A2(n782), .ZN(G153) );
  INV_X1 U836 ( .A(G171), .ZN(G301) );
  NAND2_X1 U837 ( .A1(G868), .A2(G301), .ZN(n760) );
  OR2_X1 U838 ( .A1(n1006), .A2(G868), .ZN(n759) );
  NAND2_X1 U839 ( .A1(n760), .A2(n759), .ZN(G284) );
  INV_X1 U840 ( .A(G868), .ZN(n804) );
  NOR2_X1 U841 ( .A1(G286), .A2(n804), .ZN(n762) );
  NOR2_X1 U842 ( .A1(G868), .A2(G299), .ZN(n761) );
  NOR2_X1 U843 ( .A1(n762), .A2(n761), .ZN(G297) );
  NAND2_X1 U844 ( .A1(n782), .A2(G559), .ZN(n763) );
  NAND2_X1 U845 ( .A1(n763), .A2(n1006), .ZN(n764) );
  XNOR2_X1 U846 ( .A(n764), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U847 ( .A1(n1006), .A2(G868), .ZN(n765) );
  NOR2_X1 U848 ( .A1(G559), .A2(n765), .ZN(n766) );
  XNOR2_X1 U849 ( .A(n766), .B(KEYINPUT70), .ZN(n768) );
  NOR2_X1 U850 ( .A1(n1007), .A2(G868), .ZN(n767) );
  NOR2_X1 U851 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U852 ( .A(KEYINPUT71), .B(n769), .Z(G282) );
  XOR2_X1 U853 ( .A(G2100), .B(KEYINPUT74), .Z(n780) );
  NAND2_X1 U854 ( .A1(n881), .A2(G99), .ZN(n770) );
  XNOR2_X1 U855 ( .A(n770), .B(KEYINPUT72), .ZN(n772) );
  NAND2_X1 U856 ( .A1(G111), .A2(n885), .ZN(n771) );
  NAND2_X1 U857 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U858 ( .A(n773), .B(KEYINPUT73), .ZN(n775) );
  NAND2_X1 U859 ( .A1(G135), .A2(n882), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n778) );
  NAND2_X1 U861 ( .A1(n886), .A2(G123), .ZN(n776) );
  XOR2_X1 U862 ( .A(KEYINPUT18), .B(n776), .Z(n777) );
  NOR2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n981) );
  XNOR2_X1 U864 ( .A(G2096), .B(n981), .ZN(n779) );
  NAND2_X1 U865 ( .A1(n780), .A2(n779), .ZN(G156) );
  NAND2_X1 U866 ( .A1(G559), .A2(n1006), .ZN(n781) );
  XOR2_X1 U867 ( .A(n1007), .B(n781), .Z(n802) );
  NAND2_X1 U868 ( .A1(n782), .A2(n802), .ZN(n795) );
  NAND2_X1 U869 ( .A1(n783), .A2(G67), .ZN(n784) );
  XNOR2_X1 U870 ( .A(n784), .B(KEYINPUT76), .ZN(n794) );
  NAND2_X1 U871 ( .A1(G93), .A2(n785), .ZN(n788) );
  NAND2_X1 U872 ( .A1(G55), .A2(n786), .ZN(n787) );
  NAND2_X1 U873 ( .A1(n788), .A2(n787), .ZN(n792) );
  NAND2_X1 U874 ( .A1(G80), .A2(n789), .ZN(n790) );
  XNOR2_X1 U875 ( .A(KEYINPUT75), .B(n790), .ZN(n791) );
  NOR2_X1 U876 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U877 ( .A1(n794), .A2(n793), .ZN(n805) );
  XNOR2_X1 U878 ( .A(n795), .B(n805), .ZN(G145) );
  XNOR2_X1 U879 ( .A(KEYINPUT19), .B(G288), .ZN(n796) );
  XNOR2_X1 U880 ( .A(n796), .B(n805), .ZN(n797) );
  XNOR2_X1 U881 ( .A(G290), .B(n797), .ZN(n800) );
  XNOR2_X1 U882 ( .A(n798), .B(G305), .ZN(n799) );
  XNOR2_X1 U883 ( .A(n800), .B(n799), .ZN(n801) );
  XNOR2_X1 U884 ( .A(G166), .B(n801), .ZN(n897) );
  XNOR2_X1 U885 ( .A(n802), .B(n897), .ZN(n803) );
  NOR2_X1 U886 ( .A1(n804), .A2(n803), .ZN(n807) );
  NOR2_X1 U887 ( .A1(G868), .A2(n805), .ZN(n806) );
  NOR2_X1 U888 ( .A1(n807), .A2(n806), .ZN(G295) );
  NAND2_X1 U889 ( .A1(G2084), .A2(G2078), .ZN(n808) );
  XOR2_X1 U890 ( .A(KEYINPUT20), .B(n808), .Z(n809) );
  NAND2_X1 U891 ( .A1(G2090), .A2(n809), .ZN(n810) );
  XNOR2_X1 U892 ( .A(KEYINPUT21), .B(n810), .ZN(n811) );
  NAND2_X1 U893 ( .A1(n811), .A2(G2072), .ZN(n812) );
  XOR2_X1 U894 ( .A(KEYINPUT83), .B(n812), .Z(G158) );
  XNOR2_X1 U895 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U896 ( .A1(G132), .A2(G82), .ZN(n813) );
  XNOR2_X1 U897 ( .A(n813), .B(KEYINPUT84), .ZN(n814) );
  XNOR2_X1 U898 ( .A(n814), .B(KEYINPUT22), .ZN(n815) );
  NOR2_X1 U899 ( .A1(G218), .A2(n815), .ZN(n816) );
  NAND2_X1 U900 ( .A1(G96), .A2(n816), .ZN(n833) );
  NAND2_X1 U901 ( .A1(G2106), .A2(n833), .ZN(n817) );
  XNOR2_X1 U902 ( .A(KEYINPUT85), .B(n817), .ZN(n822) );
  NAND2_X1 U903 ( .A1(G69), .A2(G120), .ZN(n818) );
  NOR2_X1 U904 ( .A1(G237), .A2(n818), .ZN(n819) );
  NAND2_X1 U905 ( .A1(G108), .A2(n819), .ZN(n832) );
  NAND2_X1 U906 ( .A1(G567), .A2(n832), .ZN(n820) );
  XOR2_X1 U907 ( .A(KEYINPUT86), .B(n820), .Z(n821) );
  NOR2_X1 U908 ( .A1(n822), .A2(n821), .ZN(G319) );
  INV_X1 U909 ( .A(G319), .ZN(n824) );
  NAND2_X1 U910 ( .A1(G483), .A2(G661), .ZN(n823) );
  NOR2_X1 U911 ( .A1(n824), .A2(n823), .ZN(n831) );
  NAND2_X1 U912 ( .A1(n831), .A2(G36), .ZN(G176) );
  NAND2_X1 U913 ( .A1(n825), .A2(G2106), .ZN(n826) );
  XOR2_X1 U914 ( .A(KEYINPUT109), .B(n826), .Z(G217) );
  NAND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n827) );
  XOR2_X1 U916 ( .A(KEYINPUT110), .B(n827), .Z(n828) );
  NAND2_X1 U917 ( .A1(n828), .A2(G661), .ZN(n829) );
  XOR2_X1 U918 ( .A(KEYINPUT111), .B(n829), .Z(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U920 ( .A1(n831), .A2(n830), .ZN(G188) );
  INV_X1 U922 ( .A(G132), .ZN(G219) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G82), .ZN(G220) );
  INV_X1 U925 ( .A(G69), .ZN(G235) );
  NOR2_X1 U926 ( .A1(n833), .A2(n832), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  XOR2_X1 U928 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n835) );
  XNOR2_X1 U929 ( .A(G2678), .B(KEYINPUT43), .ZN(n834) );
  XNOR2_X1 U930 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U931 ( .A(KEYINPUT42), .B(G2090), .Z(n837) );
  XNOR2_X1 U932 ( .A(G2067), .B(G2072), .ZN(n836) );
  XNOR2_X1 U933 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U934 ( .A(n839), .B(n838), .Z(n841) );
  XNOR2_X1 U935 ( .A(G2100), .B(G2096), .ZN(n840) );
  XNOR2_X1 U936 ( .A(n841), .B(n840), .ZN(n843) );
  XOR2_X1 U937 ( .A(G2084), .B(G2078), .Z(n842) );
  XNOR2_X1 U938 ( .A(n843), .B(n842), .ZN(G227) );
  XOR2_X1 U939 ( .A(G1986), .B(G1976), .Z(n845) );
  XNOR2_X1 U940 ( .A(G1961), .B(G1971), .ZN(n844) );
  XNOR2_X1 U941 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U942 ( .A(n846), .B(G2474), .Z(n848) );
  XNOR2_X1 U943 ( .A(G1966), .B(G1981), .ZN(n847) );
  XNOR2_X1 U944 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U945 ( .A(KEYINPUT41), .B(G1991), .Z(n850) );
  XNOR2_X1 U946 ( .A(G1996), .B(G1956), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(n851) );
  XNOR2_X1 U948 ( .A(n852), .B(n851), .ZN(G229) );
  NAND2_X1 U949 ( .A1(n886), .A2(G124), .ZN(n853) );
  XNOR2_X1 U950 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U951 ( .A1(G100), .A2(n881), .ZN(n854) );
  NAND2_X1 U952 ( .A1(n855), .A2(n854), .ZN(n859) );
  NAND2_X1 U953 ( .A1(G112), .A2(n885), .ZN(n857) );
  NAND2_X1 U954 ( .A1(G136), .A2(n882), .ZN(n856) );
  NAND2_X1 U955 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U956 ( .A1(n859), .A2(n858), .ZN(G162) );
  XOR2_X1 U957 ( .A(KEYINPUT116), .B(KEYINPUT115), .Z(n861) );
  XNOR2_X1 U958 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(n866) );
  XNOR2_X1 U960 ( .A(G164), .B(n862), .ZN(n864) );
  XNOR2_X1 U961 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U962 ( .A(n866), .B(n865), .ZN(n879) );
  NAND2_X1 U963 ( .A1(G106), .A2(n881), .ZN(n868) );
  NAND2_X1 U964 ( .A1(G142), .A2(n882), .ZN(n867) );
  NAND2_X1 U965 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U966 ( .A(n869), .B(KEYINPUT45), .ZN(n874) );
  NAND2_X1 U967 ( .A1(G118), .A2(n885), .ZN(n871) );
  NAND2_X1 U968 ( .A1(G130), .A2(n886), .ZN(n870) );
  NAND2_X1 U969 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U970 ( .A(KEYINPUT114), .B(n872), .Z(n873) );
  NAND2_X1 U971 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U972 ( .A(n875), .B(n981), .ZN(n876) );
  XNOR2_X1 U973 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U974 ( .A(n879), .B(n878), .ZN(n880) );
  XOR2_X1 U975 ( .A(n880), .B(G162), .Z(n893) );
  NAND2_X1 U976 ( .A1(G103), .A2(n881), .ZN(n884) );
  NAND2_X1 U977 ( .A1(G139), .A2(n882), .ZN(n883) );
  NAND2_X1 U978 ( .A1(n884), .A2(n883), .ZN(n891) );
  NAND2_X1 U979 ( .A1(G115), .A2(n885), .ZN(n888) );
  NAND2_X1 U980 ( .A1(G127), .A2(n886), .ZN(n887) );
  NAND2_X1 U981 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U982 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U983 ( .A1(n891), .A2(n890), .ZN(n969) );
  XNOR2_X1 U984 ( .A(G160), .B(n969), .ZN(n892) );
  XNOR2_X1 U985 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U986 ( .A1(G37), .A2(n894), .ZN(G395) );
  XNOR2_X1 U987 ( .A(n1007), .B(G286), .ZN(n896) );
  XNOR2_X1 U988 ( .A(G171), .B(n1006), .ZN(n895) );
  XNOR2_X1 U989 ( .A(n896), .B(n895), .ZN(n898) );
  XNOR2_X1 U990 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U991 ( .A1(G37), .A2(n899), .ZN(G397) );
  XNOR2_X1 U992 ( .A(G2451), .B(G2427), .ZN(n909) );
  XOR2_X1 U993 ( .A(KEYINPUT107), .B(G2443), .Z(n901) );
  XNOR2_X1 U994 ( .A(G2435), .B(G2438), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n905) );
  XOR2_X1 U996 ( .A(G2454), .B(G2430), .Z(n903) );
  XNOR2_X1 U997 ( .A(G1348), .B(G1341), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U999 ( .A(n905), .B(n904), .Z(n907) );
  XNOR2_X1 U1000 ( .A(G2446), .B(KEYINPUT108), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1002 ( .A(n909), .B(n908), .ZN(n910) );
  NAND2_X1 U1003 ( .A1(n910), .A2(G14), .ZN(n917) );
  NAND2_X1 U1004 ( .A1(G319), .A2(n917), .ZN(n914) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n911) );
  XOR2_X1 U1006 ( .A(KEYINPUT49), .B(n911), .Z(n912) );
  XNOR2_X1 U1007 ( .A(n912), .B(KEYINPUT117), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(n914), .A2(n913), .ZN(n916) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1010 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(G108), .ZN(G238) );
  INV_X1 U1013 ( .A(G96), .ZN(G221) );
  INV_X1 U1014 ( .A(n917), .ZN(G401) );
  XNOR2_X1 U1015 ( .A(G5), .B(n918), .ZN(n933) );
  XNOR2_X1 U1016 ( .A(G6), .B(G1981), .ZN(n919) );
  XNOR2_X1 U1017 ( .A(n919), .B(KEYINPUT127), .ZN(n924) );
  XOR2_X1 U1018 ( .A(G1348), .B(KEYINPUT59), .Z(n920) );
  XNOR2_X1 U1019 ( .A(G4), .B(n920), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(G19), .B(G1341), .ZN(n921) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n928) );
  XOR2_X1 U1023 ( .A(KEYINPUT126), .B(n925), .Z(n926) );
  XNOR2_X1 U1024 ( .A(G20), .B(n926), .ZN(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1026 ( .A(KEYINPUT60), .B(n929), .Z(n931) );
  XNOR2_X1 U1027 ( .A(G1966), .B(G21), .ZN(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n940) );
  XNOR2_X1 U1030 ( .A(G1971), .B(G22), .ZN(n935) );
  XNOR2_X1 U1031 ( .A(G23), .B(G1976), .ZN(n934) );
  NOR2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n937) );
  XOR2_X1 U1033 ( .A(G1986), .B(G24), .Z(n936) );
  NAND2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1035 ( .A(KEYINPUT58), .B(n938), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1037 ( .A(n941), .B(KEYINPUT61), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(G16), .B(KEYINPUT125), .ZN(n942) );
  NAND2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1040 ( .A1(G11), .A2(n944), .ZN(n968) );
  XOR2_X1 U1041 ( .A(G1991), .B(G25), .Z(n945) );
  NAND2_X1 U1042 ( .A1(n945), .A2(G28), .ZN(n956) );
  XOR2_X1 U1043 ( .A(G1996), .B(KEYINPUT119), .Z(n946) );
  XNOR2_X1 U1044 ( .A(G32), .B(n946), .ZN(n949) );
  XOR2_X1 U1045 ( .A(n947), .B(G27), .Z(n948) );
  NOR2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(KEYINPUT120), .B(n950), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(G2067), .B(G26), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(G33), .B(G2072), .ZN(n951) );
  NOR2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1053 ( .A(KEYINPUT53), .B(n957), .Z(n961) );
  XNOR2_X1 U1054 ( .A(KEYINPUT54), .B(G34), .ZN(n958) );
  XNOR2_X1 U1055 ( .A(n958), .B(KEYINPUT121), .ZN(n959) );
  XNOR2_X1 U1056 ( .A(G2084), .B(n959), .ZN(n960) );
  NAND2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(G35), .B(G2090), .ZN(n962) );
  NOR2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1060 ( .A(KEYINPUT55), .B(n964), .Z(n965) );
  NOR2_X1 U1061 ( .A1(G29), .A2(n965), .ZN(n966) );
  XNOR2_X1 U1062 ( .A(n966), .B(KEYINPUT122), .ZN(n967) );
  NOR2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n996) );
  XOR2_X1 U1064 ( .A(G2072), .B(n969), .Z(n971) );
  XOR2_X1 U1065 ( .A(G164), .B(G2078), .Z(n970) );
  NOR2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(KEYINPUT50), .B(n972), .ZN(n977) );
  XOR2_X1 U1068 ( .A(G2090), .B(G162), .Z(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1070 ( .A(KEYINPUT51), .B(n975), .Z(n976) );
  NAND2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n990) );
  XOR2_X1 U1072 ( .A(G2084), .B(G160), .Z(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n983) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(n986), .B(KEYINPUT118), .ZN(n987) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1080 ( .A(KEYINPUT52), .B(n991), .ZN(n993) );
  INV_X1 U1081 ( .A(KEYINPUT55), .ZN(n992) );
  NAND2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1083 ( .A1(n994), .A2(G29), .ZN(n995) );
  NAND2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n1023) );
  XOR2_X1 U1085 ( .A(G16), .B(KEYINPUT56), .Z(n1021) );
  XNOR2_X1 U1086 ( .A(G1966), .B(G168), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(n999), .B(KEYINPUT57), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(G1971), .A2(G303), .ZN(n1000) );
  NAND2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1018) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(G1956), .B(G299), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1011) );
  XOR2_X1 U1094 ( .A(G1348), .B(n1006), .Z(n1009) );
  XNOR2_X1 U1095 ( .A(n1007), .B(G1341), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1014) );
  XOR2_X1 U1098 ( .A(G1961), .B(G301), .Z(n1012) );
  XNOR2_X1 U1099 ( .A(KEYINPUT123), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1103 ( .A(KEYINPUT124), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1104 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1105 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1106 ( .A(n1024), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

