

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  NOR2_X1 U322 ( .A1(n512), .A2(n417), .ZN(n569) );
  XOR2_X1 U323 ( .A(n375), .B(KEYINPUT77), .Z(n290) );
  NOR2_X1 U324 ( .A1(n470), .A2(n402), .ZN(n403) );
  INV_X1 U325 ( .A(G78GAT), .ZN(n380) );
  OR2_X1 U326 ( .A1(n459), .A2(n525), .ZN(n416) );
  XNOR2_X1 U327 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U328 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U329 ( .A(n451), .B(n450), .ZN(n526) );
  INV_X1 U330 ( .A(G169GAT), .ZN(n454) );
  XOR2_X1 U331 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n292) );
  XNOR2_X1 U332 ( .A(G8GAT), .B(KEYINPUT30), .ZN(n291) );
  XNOR2_X1 U333 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U334 ( .A(G50GAT), .B(G36GAT), .Z(n294) );
  XOR2_X1 U335 ( .A(G15GAT), .B(G1GAT), .Z(n379) );
  XNOR2_X1 U336 ( .A(n379), .B(KEYINPUT67), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U338 ( .A(n296), .B(n295), .Z(n298) );
  NAND2_X1 U339 ( .A1(G229GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U340 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U341 ( .A(G197GAT), .B(G22GAT), .Z(n300) );
  XNOR2_X1 U342 ( .A(G169GAT), .B(G141GAT), .ZN(n299) );
  XNOR2_X1 U343 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U344 ( .A(n302), .B(n301), .Z(n310) );
  XOR2_X1 U345 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n304) );
  XNOR2_X1 U346 ( .A(G43GAT), .B(G29GAT), .ZN(n303) );
  XNOR2_X1 U347 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U348 ( .A(KEYINPUT69), .B(n305), .Z(n364) );
  XOR2_X1 U349 ( .A(KEYINPUT70), .B(KEYINPUT65), .Z(n307) );
  XNOR2_X1 U350 ( .A(G113GAT), .B(KEYINPUT66), .ZN(n306) );
  XNOR2_X1 U351 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U352 ( .A(n364), .B(n308), .ZN(n309) );
  XNOR2_X1 U353 ( .A(n310), .B(n309), .ZN(n570) );
  XOR2_X1 U354 ( .A(KEYINPUT87), .B(KEYINPUT4), .Z(n312) );
  XNOR2_X1 U355 ( .A(KEYINPUT90), .B(KEYINPUT88), .ZN(n311) );
  XNOR2_X1 U356 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U357 ( .A(KEYINPUT1), .B(KEYINPUT92), .Z(n314) );
  XNOR2_X1 U358 ( .A(KEYINPUT5), .B(KEYINPUT6), .ZN(n313) );
  XNOR2_X1 U359 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U360 ( .A(n316), .B(n315), .Z(n326) );
  XOR2_X1 U361 ( .A(G127GAT), .B(G134GAT), .Z(n318) );
  XNOR2_X1 U362 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n317) );
  XNOR2_X1 U363 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U364 ( .A(G113GAT), .B(n319), .ZN(n450) );
  XOR2_X1 U365 ( .A(KEYINPUT83), .B(KEYINPUT3), .Z(n321) );
  XNOR2_X1 U366 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n320) );
  XNOR2_X1 U367 ( .A(n321), .B(n320), .ZN(n429) );
  XOR2_X1 U368 ( .A(KEYINPUT89), .B(n429), .Z(n323) );
  NAND2_X1 U369 ( .A1(G225GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U370 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U371 ( .A(n450), .B(n324), .Z(n325) );
  XNOR2_X1 U372 ( .A(n326), .B(n325), .ZN(n334) );
  XOR2_X1 U373 ( .A(KEYINPUT91), .B(G57GAT), .Z(n328) );
  XNOR2_X1 U374 ( .A(G1GAT), .B(G148GAT), .ZN(n327) );
  XNOR2_X1 U375 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U376 ( .A(G85GAT), .B(G155GAT), .Z(n330) );
  XNOR2_X1 U377 ( .A(G29GAT), .B(G162GAT), .ZN(n329) );
  XNOR2_X1 U378 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U379 ( .A(n332), .B(n331), .Z(n333) );
  XNOR2_X1 U380 ( .A(n334), .B(n333), .ZN(n512) );
  XOR2_X1 U381 ( .A(KEYINPUT21), .B(G218GAT), .Z(n336) );
  XNOR2_X1 U382 ( .A(KEYINPUT81), .B(KEYINPUT82), .ZN(n335) );
  XNOR2_X1 U383 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U384 ( .A(G197GAT), .B(n337), .ZN(n434) );
  XNOR2_X1 U385 ( .A(G8GAT), .B(G183GAT), .ZN(n338) );
  XNOR2_X1 U386 ( .A(n338), .B(G211GAT), .ZN(n369) );
  XOR2_X1 U387 ( .A(G36GAT), .B(G190GAT), .Z(n353) );
  XOR2_X1 U388 ( .A(n369), .B(n353), .Z(n340) );
  NAND2_X1 U389 ( .A1(G226GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U391 ( .A(n341), .B(KEYINPUT93), .Z(n345) );
  XOR2_X1 U392 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n343) );
  XNOR2_X1 U393 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n342) );
  XNOR2_X1 U394 ( .A(n343), .B(n342), .ZN(n439) );
  XNOR2_X1 U395 ( .A(n439), .B(KEYINPUT94), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U397 ( .A(n434), .B(n346), .Z(n350) );
  XOR2_X1 U398 ( .A(G92GAT), .B(G64GAT), .Z(n348) );
  XNOR2_X1 U399 ( .A(G204GAT), .B(KEYINPUT72), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U401 ( .A(G176GAT), .B(n349), .ZN(n397) );
  XNOR2_X1 U402 ( .A(n350), .B(n397), .ZN(n459) );
  XOR2_X1 U403 ( .A(KEYINPUT75), .B(KEYINPUT64), .Z(n352) );
  XNOR2_X1 U404 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n351) );
  XNOR2_X1 U405 ( .A(n352), .B(n351), .ZN(n363) );
  XOR2_X1 U406 ( .A(KEYINPUT11), .B(n353), .Z(n355) );
  XOR2_X1 U407 ( .A(G99GAT), .B(G85GAT), .Z(n394) );
  XNOR2_X1 U408 ( .A(G218GAT), .B(n394), .ZN(n354) );
  XNOR2_X1 U409 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U410 ( .A(KEYINPUT10), .B(G92GAT), .Z(n357) );
  NAND2_X1 U411 ( .A1(G232GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U413 ( .A(n359), .B(n358), .Z(n361) );
  XOR2_X1 U414 ( .A(G50GAT), .B(G162GAT), .Z(n419) );
  XNOR2_X1 U415 ( .A(n419), .B(G106GAT), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n363), .B(n362), .ZN(n365) );
  XNOR2_X1 U418 ( .A(n365), .B(n364), .ZN(n561) );
  INV_X1 U419 ( .A(n561), .ZN(n470) );
  XOR2_X1 U420 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n367) );
  XNOR2_X1 U421 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n367), .B(n366), .ZN(n385) );
  XOR2_X1 U423 ( .A(G22GAT), .B(G155GAT), .Z(n425) );
  INV_X1 U424 ( .A(n425), .ZN(n368) );
  NAND2_X1 U425 ( .A1(n369), .A2(n368), .ZN(n372) );
  INV_X1 U426 ( .A(n369), .ZN(n370) );
  NAND2_X1 U427 ( .A1(n370), .A2(n425), .ZN(n371) );
  NAND2_X1 U428 ( .A1(n372), .A2(n371), .ZN(n374) );
  NAND2_X1 U429 ( .A1(G231GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U430 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U431 ( .A(KEYINPUT71), .B(KEYINPUT13), .Z(n377) );
  XNOR2_X1 U432 ( .A(G71GAT), .B(G57GAT), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n377), .B(n376), .ZN(n390) );
  XNOR2_X1 U434 ( .A(n390), .B(KEYINPUT76), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n290), .B(n378), .ZN(n383) );
  XNOR2_X1 U436 ( .A(n379), .B(G127GAT), .ZN(n381) );
  XOR2_X1 U437 ( .A(n385), .B(n384), .Z(n578) );
  XOR2_X1 U438 ( .A(KEYINPUT109), .B(n578), .Z(n557) );
  XOR2_X1 U439 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n387) );
  NAND2_X1 U440 ( .A1(G230GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U441 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U442 ( .A(n388), .B(KEYINPUT32), .Z(n392) );
  XNOR2_X1 U443 ( .A(G106GAT), .B(G78GAT), .ZN(n389) );
  XNOR2_X1 U444 ( .A(n389), .B(G148GAT), .ZN(n418) );
  XNOR2_X1 U445 ( .A(n418), .B(n390), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U447 ( .A(n393), .B(KEYINPUT73), .Z(n396) );
  XNOR2_X1 U448 ( .A(G120GAT), .B(n394), .ZN(n395) );
  XNOR2_X1 U449 ( .A(n396), .B(n395), .ZN(n398) );
  XNOR2_X1 U450 ( .A(n398), .B(n397), .ZN(n573) );
  XNOR2_X1 U451 ( .A(n573), .B(KEYINPUT41), .ZN(n551) );
  NOR2_X1 U452 ( .A1(n570), .A2(n551), .ZN(n400) );
  XOR2_X1 U453 ( .A(KEYINPUT46), .B(KEYINPUT110), .Z(n399) );
  XNOR2_X1 U454 ( .A(n400), .B(n399), .ZN(n401) );
  NAND2_X1 U455 ( .A1(n557), .A2(n401), .ZN(n402) );
  NAND2_X1 U456 ( .A1(n403), .A2(KEYINPUT47), .ZN(n407) );
  INV_X1 U457 ( .A(n403), .ZN(n405) );
  INV_X1 U458 ( .A(KEYINPUT47), .ZN(n404) );
  NAND2_X1 U459 ( .A1(n405), .A2(n404), .ZN(n406) );
  NAND2_X1 U460 ( .A1(n407), .A2(n406), .ZN(n414) );
  XNOR2_X1 U461 ( .A(KEYINPUT36), .B(n561), .ZN(n581) );
  NOR2_X1 U462 ( .A1(n581), .A2(n578), .ZN(n408) );
  XNOR2_X1 U463 ( .A(n408), .B(KEYINPUT111), .ZN(n409) );
  XNOR2_X1 U464 ( .A(KEYINPUT45), .B(n409), .ZN(n410) );
  NOR2_X1 U465 ( .A1(n573), .A2(n410), .ZN(n411) );
  XNOR2_X1 U466 ( .A(KEYINPUT112), .B(n411), .ZN(n412) );
  NAND2_X1 U467 ( .A1(n412), .A2(n570), .ZN(n413) );
  NAND2_X1 U468 ( .A1(n414), .A2(n413), .ZN(n415) );
  XOR2_X1 U469 ( .A(KEYINPUT48), .B(n415), .Z(n525) );
  XNOR2_X1 U470 ( .A(KEYINPUT54), .B(n416), .ZN(n417) );
  XOR2_X1 U471 ( .A(n419), .B(n418), .Z(n421) );
  NAND2_X1 U472 ( .A1(G228GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U473 ( .A(n421), .B(n420), .ZN(n433) );
  XOR2_X1 U474 ( .A(G204GAT), .B(G211GAT), .Z(n423) );
  XNOR2_X1 U475 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n422) );
  XNOR2_X1 U476 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U477 ( .A(n424), .B(KEYINPUT85), .Z(n427) );
  XNOR2_X1 U478 ( .A(n425), .B(KEYINPUT23), .ZN(n426) );
  XNOR2_X1 U479 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U480 ( .A(n428), .B(KEYINPUT86), .Z(n431) );
  XNOR2_X1 U481 ( .A(n429), .B(KEYINPUT84), .ZN(n430) );
  XNOR2_X1 U482 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U483 ( .A(n433), .B(n432), .ZN(n435) );
  XNOR2_X1 U484 ( .A(n435), .B(n434), .ZN(n466) );
  NAND2_X1 U485 ( .A1(n569), .A2(n466), .ZN(n436) );
  XNOR2_X1 U486 ( .A(n436), .B(KEYINPUT55), .ZN(n452) );
  XOR2_X1 U487 ( .A(G71GAT), .B(KEYINPUT78), .Z(n438) );
  XNOR2_X1 U488 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n449) );
  XOR2_X1 U490 ( .A(G99GAT), .B(G190GAT), .Z(n441) );
  XNOR2_X1 U491 ( .A(n439), .B(KEYINPUT79), .ZN(n440) );
  XNOR2_X1 U492 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U493 ( .A(G183GAT), .B(G176GAT), .Z(n443) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U495 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U496 ( .A(n445), .B(n444), .Z(n447) );
  XNOR2_X1 U497 ( .A(G43GAT), .B(KEYINPUT80), .ZN(n446) );
  XNOR2_X1 U498 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U499 ( .A(n449), .B(n448), .ZN(n451) );
  NAND2_X1 U500 ( .A1(n452), .A2(n526), .ZN(n560) );
  NOR2_X1 U501 ( .A1(n570), .A2(n560), .ZN(n453) );
  XNOR2_X1 U502 ( .A(n454), .B(n453), .ZN(G1348GAT) );
  XNOR2_X1 U503 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n475) );
  NOR2_X1 U504 ( .A1(n570), .A2(n573), .ZN(n455) );
  XOR2_X1 U505 ( .A(KEYINPUT74), .B(n455), .Z(n487) );
  INV_X1 U506 ( .A(n459), .ZN(n515) );
  NAND2_X1 U507 ( .A1(n526), .A2(n515), .ZN(n456) );
  NAND2_X1 U508 ( .A1(n456), .A2(n466), .ZN(n457) );
  XNOR2_X1 U509 ( .A(n457), .B(KEYINPUT95), .ZN(n458) );
  XNOR2_X1 U510 ( .A(KEYINPUT25), .B(n458), .ZN(n462) );
  XOR2_X1 U511 ( .A(KEYINPUT27), .B(n459), .Z(n465) );
  NOR2_X1 U512 ( .A1(n466), .A2(n526), .ZN(n460) );
  XNOR2_X1 U513 ( .A(n460), .B(KEYINPUT26), .ZN(n568) );
  NAND2_X1 U514 ( .A1(n465), .A2(n568), .ZN(n461) );
  NAND2_X1 U515 ( .A1(n462), .A2(n461), .ZN(n463) );
  XOR2_X1 U516 ( .A(KEYINPUT96), .B(n463), .Z(n464) );
  NOR2_X1 U517 ( .A1(n512), .A2(n464), .ZN(n469) );
  NAND2_X1 U518 ( .A1(n512), .A2(n465), .ZN(n524) );
  XNOR2_X1 U519 ( .A(KEYINPUT28), .B(n466), .ZN(n528) );
  INV_X1 U520 ( .A(n528), .ZN(n518) );
  OR2_X1 U521 ( .A1(n518), .A2(n526), .ZN(n467) );
  NOR2_X1 U522 ( .A1(n524), .A2(n467), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n469), .A2(n468), .ZN(n483) );
  NOR2_X1 U524 ( .A1(n578), .A2(n470), .ZN(n471) );
  XOR2_X1 U525 ( .A(KEYINPUT16), .B(n471), .Z(n472) );
  NOR2_X1 U526 ( .A1(n483), .A2(n472), .ZN(n473) );
  XNOR2_X1 U527 ( .A(KEYINPUT97), .B(n473), .ZN(n500) );
  NOR2_X1 U528 ( .A1(n487), .A2(n500), .ZN(n480) );
  NAND2_X1 U529 ( .A1(n480), .A2(n512), .ZN(n474) );
  XNOR2_X1 U530 ( .A(n475), .B(n474), .ZN(G1324GAT) );
  NAND2_X1 U531 ( .A1(n480), .A2(n515), .ZN(n476) );
  XNOR2_X1 U532 ( .A(n476), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U533 ( .A(KEYINPUT98), .B(KEYINPUT35), .Z(n478) );
  NAND2_X1 U534 ( .A1(n480), .A2(n526), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U536 ( .A(G15GAT), .B(n479), .ZN(G1326GAT) );
  XOR2_X1 U537 ( .A(G22GAT), .B(KEYINPUT99), .Z(n482) );
  NAND2_X1 U538 ( .A1(n480), .A2(n518), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(G1327GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT37), .B(KEYINPUT100), .Z(n486) );
  NOR2_X1 U541 ( .A1(n581), .A2(n483), .ZN(n484) );
  NAND2_X1 U542 ( .A1(n578), .A2(n484), .ZN(n485) );
  XNOR2_X1 U543 ( .A(n486), .B(n485), .ZN(n511) );
  NOR2_X1 U544 ( .A1(n511), .A2(n487), .ZN(n488) );
  XNOR2_X1 U545 ( .A(KEYINPUT38), .B(n488), .ZN(n496) );
  NAND2_X1 U546 ( .A1(n496), .A2(n512), .ZN(n491) );
  XNOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n489), .B(KEYINPUT39), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  NAND2_X1 U550 ( .A1(n496), .A2(n515), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n492), .B(KEYINPUT102), .ZN(n493) );
  XNOR2_X1 U552 ( .A(G36GAT), .B(n493), .ZN(G1329GAT) );
  NAND2_X1 U553 ( .A1(n496), .A2(n526), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n494), .B(KEYINPUT40), .ZN(n495) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  NAND2_X1 U556 ( .A1(n518), .A2(n496), .ZN(n497) );
  XNOR2_X1 U557 ( .A(G50GAT), .B(n497), .ZN(G1331GAT) );
  INV_X1 U558 ( .A(n570), .ZN(n498) );
  NOR2_X1 U559 ( .A1(n551), .A2(n498), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n499), .B(KEYINPUT103), .ZN(n510) );
  NOR2_X1 U561 ( .A1(n500), .A2(n510), .ZN(n507) );
  NAND2_X1 U562 ( .A1(n512), .A2(n507), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n501), .B(KEYINPUT42), .ZN(n502) );
  XNOR2_X1 U564 ( .A(G57GAT), .B(n502), .ZN(G1332GAT) );
  NAND2_X1 U565 ( .A1(n507), .A2(n515), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n503), .B(KEYINPUT104), .ZN(n504) );
  XNOR2_X1 U567 ( .A(G64GAT), .B(n504), .ZN(G1333GAT) );
  XOR2_X1 U568 ( .A(G71GAT), .B(KEYINPUT105), .Z(n506) );
  NAND2_X1 U569 ( .A1(n507), .A2(n526), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n506), .B(n505), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(G78GAT), .B(KEYINPUT43), .Z(n509) );
  NAND2_X1 U572 ( .A1(n507), .A2(n518), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(KEYINPUT106), .ZN(n514) );
  NOR2_X1 U575 ( .A1(n511), .A2(n510), .ZN(n519) );
  NAND2_X1 U576 ( .A1(n519), .A2(n512), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n514), .B(n513), .ZN(G1336GAT) );
  NAND2_X1 U578 ( .A1(n519), .A2(n515), .ZN(n516) );
  XNOR2_X1 U579 ( .A(n516), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U580 ( .A1(n526), .A2(n519), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n517), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U582 ( .A(G106GAT), .B(KEYINPUT107), .ZN(n523) );
  XOR2_X1 U583 ( .A(KEYINPUT108), .B(KEYINPUT44), .Z(n521) );
  NAND2_X1 U584 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n523), .B(n522), .ZN(G1339GAT) );
  NOR2_X1 U587 ( .A1(n525), .A2(n524), .ZN(n540) );
  NAND2_X1 U588 ( .A1(n540), .A2(n526), .ZN(n527) );
  XNOR2_X1 U589 ( .A(KEYINPUT113), .B(n527), .ZN(n529) );
  NAND2_X1 U590 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U591 ( .A(KEYINPUT114), .B(n530), .ZN(n537) );
  NOR2_X1 U592 ( .A1(n570), .A2(n537), .ZN(n531) );
  XOR2_X1 U593 ( .A(G113GAT), .B(n531), .Z(G1340GAT) );
  NOR2_X1 U594 ( .A1(n537), .A2(n551), .ZN(n533) );
  XNOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  XNOR2_X1 U597 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n535) );
  NOR2_X1 U598 ( .A1(n557), .A2(n537), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XNOR2_X1 U601 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n539) );
  NOR2_X1 U602 ( .A1(n561), .A2(n537), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  NAND2_X1 U604 ( .A1(n540), .A2(n568), .ZN(n549) );
  NOR2_X1 U605 ( .A1(n570), .A2(n549), .ZN(n541) );
  XOR2_X1 U606 ( .A(G141GAT), .B(n541), .Z(G1344GAT) );
  NOR2_X1 U607 ( .A1(n551), .A2(n549), .ZN(n546) );
  XOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n543) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U611 ( .A(KEYINPUT52), .B(n544), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  NOR2_X1 U613 ( .A1(n578), .A2(n549), .ZN(n547) );
  XOR2_X1 U614 ( .A(KEYINPUT118), .B(n547), .Z(n548) );
  XNOR2_X1 U615 ( .A(G155GAT), .B(n548), .ZN(G1346GAT) );
  NOR2_X1 U616 ( .A1(n561), .A2(n549), .ZN(n550) );
  XOR2_X1 U617 ( .A(G162GAT), .B(n550), .Z(G1347GAT) );
  NOR2_X1 U618 ( .A1(n551), .A2(n560), .ZN(n556) );
  XOR2_X1 U619 ( .A(KEYINPUT57), .B(KEYINPUT120), .Z(n553) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(KEYINPUT119), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U622 ( .A(KEYINPUT56), .B(n554), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(G1349GAT) );
  NOR2_X1 U624 ( .A1(n557), .A2(n560), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G183GAT), .B(KEYINPUT121), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1350GAT) );
  NOR2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n565) );
  XOR2_X1 U628 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n563) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(KEYINPUT123), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U631 ( .A(n565), .B(n564), .Z(G1351GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n567) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n572) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n580) );
  NOR2_X1 U636 ( .A1(n570), .A2(n580), .ZN(n571) );
  XOR2_X1 U637 ( .A(n572), .B(n571), .Z(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n576) );
  INV_X1 U639 ( .A(n580), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U642 ( .A(G204GAT), .B(n577), .Z(G1353GAT) );
  OR2_X1 U643 ( .A1(n578), .A2(n580), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(G218GAT), .B(n584), .Z(G1355GAT) );
endmodule

