//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT15), .ZN(new_n203));
  OR2_X1    g002(.A1(KEYINPUT88), .A2(G43gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(KEYINPUT88), .A2(G43gat), .ZN(new_n205));
  AOI21_X1  g004(.A(G50gat), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT89), .ZN(new_n207));
  INV_X1    g006(.A(G50gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(new_n208), .B2(G43gat), .ZN(new_n209));
  INV_X1    g008(.A(G43gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n210), .A2(KEYINPUT89), .A3(G50gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n203), .B1(new_n206), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT15), .B1(new_n208), .B2(G43gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n210), .A2(G50gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  INV_X1    g017(.A(G36gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n220), .A2(KEYINPUT14), .B1(new_n221), .B2(new_n219), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  AND3_X1   g022(.A1(new_n213), .A2(new_n223), .A3(KEYINPUT90), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT90), .B1(new_n213), .B2(new_n223), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n214), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT86), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n228), .A2(new_n229), .B1(new_n221), .B2(new_n219), .ZN(new_n230));
  OAI211_X1 g029(.A(KEYINPUT86), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n227), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n215), .A2(new_n216), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT87), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n228), .A2(new_n229), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n219), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n237), .A3(new_n231), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n214), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT87), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n240), .A3(new_n233), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n235), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n202), .B1(new_n226), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n213), .A2(new_n223), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT90), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n213), .A2(new_n223), .A3(KEYINPUT90), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n235), .A2(new_n241), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n249), .A3(KEYINPUT91), .ZN(new_n250));
  XOR2_X1   g049(.A(KEYINPUT92), .B(KEYINPUT17), .Z(new_n251));
  NAND3_X1  g050(.A1(new_n243), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G15gat), .B(G22gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT16), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n253), .B1(new_n254), .B2(G1gat), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n255), .B1(G1gat), .B2(new_n253), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(G8gat), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n242), .B1(new_n246), .B2(new_n247), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n257), .B1(new_n258), .B2(KEYINPUT17), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G229gat), .A2(G233gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n250), .A3(new_n257), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT93), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT18), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n260), .A2(KEYINPUT93), .A3(new_n261), .A4(new_n262), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT94), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n260), .A2(KEYINPUT18), .A3(new_n261), .A4(new_n262), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n261), .B(KEYINPUT13), .Z(new_n271));
  INV_X1    g070(.A(new_n262), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n257), .B1(new_n243), .B2(new_n250), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n268), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G113gat), .B(G141gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT85), .B(G197gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  XOR2_X1   g079(.A(KEYINPUT11), .B(G169gat), .Z(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT12), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n269), .A2(new_n277), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT18), .B1(new_n263), .B2(new_n264), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n275), .B1(new_n286), .B2(new_n267), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT94), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n288), .B1(new_n286), .B2(new_n267), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n287), .B1(new_n289), .B2(new_n283), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT95), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT40), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT4), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT2), .ZN(new_n296));
  INV_X1    g095(.A(G155gat), .ZN(new_n297));
  INV_X1    g096(.A(G162gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(new_n297), .B2(new_n298), .ZN(new_n300));
  INV_X1    g099(.A(G141gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G148gat), .ZN(new_n302));
  INV_X1    g101(.A(G148gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G141gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n303), .A2(G141gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT73), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n300), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  XOR2_X1   g108(.A(G155gat), .B(G162gat), .Z(new_n310));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n311));
  XNOR2_X1  g110(.A(G141gat), .B(G148gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n296), .A2(KEYINPUT71), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT71), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT2), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n310), .B(new_n311), .C1(new_n312), .C2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n301), .A2(G148gat), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n313), .B(new_n315), .C1(new_n307), .C2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n311), .B1(new_n320), .B2(new_n310), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n309), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT67), .ZN(new_n323));
  INV_X1    g122(.A(G113gat), .ZN(new_n324));
  INV_X1    g123(.A(G120gat), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT1), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G113gat), .A2(G120gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G134gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G127gat), .ZN(new_n330));
  INV_X1    g129(.A(G127gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G134gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n326), .A2(new_n327), .B1(new_n330), .B2(new_n332), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n323), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n328), .A2(new_n333), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n326), .A2(new_n327), .A3(new_n330), .A4(new_n332), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(KEYINPUT67), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n295), .B1(new_n322), .B2(new_n340), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n300), .A2(new_n306), .A3(new_n308), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n310), .B1(new_n312), .B2(new_n316), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT72), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n342), .B1(new_n344), .B2(new_n317), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n334), .A2(new_n335), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(KEYINPUT4), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n346), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT3), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n348), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n322), .A2(KEYINPUT3), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n341), .B(new_n347), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT39), .ZN(new_n353));
  NAND2_X1  g152(.A1(G225gat), .A2(G233gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G57gat), .B(G85gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n357), .B(KEYINPUT75), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT74), .B(KEYINPUT0), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G1gat), .B(G29gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n356), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n322), .A2(new_n348), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n346), .B(new_n309), .C1(new_n318), .C2(new_n321), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n365), .A3(new_n354), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT39), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(new_n355), .B2(new_n352), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n294), .B1(new_n363), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n365), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n344), .A2(new_n317), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n346), .B1(new_n371), .B2(new_n309), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n355), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n334), .A2(new_n323), .A3(new_n335), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT67), .B1(new_n337), .B2(new_n338), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(KEYINPUT4), .A3(new_n345), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n365), .A2(new_n295), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n378), .A3(new_n354), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n350), .A2(new_n351), .ZN(new_n380));
  OAI211_X1 g179(.A(KEYINPUT5), .B(new_n373), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n322), .A2(KEYINPUT3), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n345), .A2(new_n349), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(new_n383), .A3(new_n348), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n355), .A2(KEYINPUT5), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n384), .A2(new_n347), .A3(new_n341), .A4(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n362), .B1(new_n381), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n352), .A2(new_n355), .ZN(new_n389));
  INV_X1    g188(.A(new_n367), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n391), .A2(KEYINPUT40), .A3(new_n362), .A4(new_n356), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n369), .A2(new_n388), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G8gat), .B(G36gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT70), .ZN(new_n395));
  XNOR2_X1  g194(.A(G64gat), .B(G92gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n395), .B(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(G226gat), .A2(G233gat), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(G169gat), .A2(G176gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT23), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT23), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n403), .B1(G169gat), .B2(G176gat), .ZN(new_n404));
  OAI211_X1 g203(.A(KEYINPUT64), .B(new_n402), .C1(new_n404), .C2(new_n401), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT25), .ZN(new_n406));
  NOR3_X1   g205(.A1(new_n403), .A2(G169gat), .A3(G176gat), .ZN(new_n407));
  INV_X1    g206(.A(new_n401), .ZN(new_n408));
  INV_X1    g207(.A(G169gat), .ZN(new_n409));
  INV_X1    g208(.A(G176gat), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT23), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n407), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n413), .A2(G190gat), .ZN(new_n414));
  INV_X1    g213(.A(G190gat), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n415), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n416));
  OR2_X1    g215(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n406), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n405), .A2(new_n412), .A3(new_n418), .A4(KEYINPUT25), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT27), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(G183gat), .ZN(new_n424));
  INV_X1    g223(.A(G183gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT27), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n426), .A3(new_n415), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT28), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT27), .B(G183gat), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(KEYINPUT28), .A3(new_n415), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(new_n431), .A3(KEYINPUT65), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT65), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n427), .A2(new_n433), .A3(new_n428), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT26), .ZN(new_n435));
  NAND2_X1  g234(.A1(G183gat), .A2(G190gat), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT26), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n437), .B1(G169gat), .B2(G176gat), .ZN(new_n438));
  AND2_X1   g237(.A1(G169gat), .A2(G176gat), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n435), .B(new_n436), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT66), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n401), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n443), .B(KEYINPUT66), .C1(new_n439), .C2(new_n438), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n432), .A2(new_n434), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n422), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT29), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n400), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AND2_X1   g247(.A1(KEYINPUT68), .A2(G218gat), .ZN(new_n449));
  NOR2_X1   g248(.A1(KEYINPUT68), .A2(G218gat), .ZN(new_n450));
  OAI21_X1  g249(.A(G211gat), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT22), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(G197gat), .B(G204gat), .ZN(new_n454));
  INV_X1    g253(.A(G211gat), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(G218gat), .ZN(new_n456));
  INV_X1    g255(.A(G218gat), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n457), .A2(G211gat), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT69), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G211gat), .B(G218gat), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT69), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n453), .A2(new_n454), .A3(new_n459), .A4(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n453), .A2(new_n454), .B1(new_n462), .B2(new_n459), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n399), .B1(new_n422), .B2(new_n445), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n448), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n466), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n442), .A2(new_n444), .A3(new_n434), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n470), .A2(new_n432), .B1(new_n420), .B2(new_n421), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n399), .B1(new_n471), .B2(KEYINPUT29), .ZN(new_n472));
  INV_X1    g271(.A(new_n467), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n398), .B1(new_n468), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n466), .B1(new_n448), .B2(new_n467), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n469), .A3(new_n473), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n477), .A3(new_n397), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n475), .A2(KEYINPUT30), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT30), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n476), .A2(new_n477), .A3(new_n480), .A4(new_n397), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT82), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n393), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n369), .A2(new_n388), .A3(new_n392), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n479), .A2(new_n481), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT82), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(G228gat), .A2(G233gat), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n447), .B1(new_n464), .B2(new_n465), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT3), .B1(new_n490), .B2(KEYINPUT78), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n453), .A2(new_n454), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n462), .A2(new_n459), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT29), .B1(new_n494), .B2(new_n463), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT78), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n345), .B1(new_n491), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT29), .B1(new_n345), .B2(new_n349), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n499), .A2(new_n469), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n489), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT80), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT3), .B1(new_n490), .B2(KEYINPUT79), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT79), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n495), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n345), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(G228gat), .B(G233gat), .C1(new_n499), .C2(new_n469), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n505), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n349), .B1(new_n495), .B2(new_n504), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n322), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n499), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n489), .B1(new_n512), .B2(new_n466), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n513), .A3(KEYINPUT80), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n501), .A2(new_n508), .A3(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G78gat), .B(G106gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT31), .B(G50gat), .ZN(new_n517));
  XOR2_X1   g316(.A(new_n516), .B(new_n517), .Z(new_n518));
  NAND2_X1  g317(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n518), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n501), .A2(new_n508), .A3(new_n514), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT81), .B(G22gat), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n519), .A2(new_n523), .A3(new_n521), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n381), .A2(new_n386), .ZN(new_n528));
  INV_X1    g327(.A(new_n362), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT76), .B(KEYINPUT6), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n528), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n379), .A2(new_n380), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n373), .A2(KEYINPUT5), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n386), .B(new_n362), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n530), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n532), .B(new_n478), .C1(new_n536), .C2(new_n387), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n476), .A2(new_n477), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n397), .B1(new_n539), .B2(KEYINPUT37), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT37), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n476), .A2(new_n477), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT38), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT38), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n540), .A2(new_n545), .A3(new_n542), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT83), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT83), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n540), .A2(new_n548), .A3(new_n545), .A4(new_n542), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n538), .A2(new_n544), .A3(new_n547), .A4(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n488), .A2(new_n527), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT84), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT84), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n488), .A2(new_n553), .A3(new_n550), .A4(new_n527), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n535), .A2(KEYINPUT77), .A3(new_n530), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT77), .B1(new_n535), .B2(new_n530), .ZN(new_n556));
  NOR3_X1   g355(.A1(new_n555), .A2(new_n556), .A3(new_n387), .ZN(new_n557));
  INV_X1    g356(.A(new_n532), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n486), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n519), .A2(new_n523), .A3(new_n521), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n523), .B1(new_n519), .B2(new_n521), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G227gat), .A2(G233gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n471), .A2(new_n376), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n446), .A2(new_n340), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT32), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n564), .A2(new_n565), .A3(new_n563), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT34), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT34), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n564), .A2(new_n565), .A3(new_n571), .A4(new_n563), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n564), .A2(new_n565), .ZN(new_n574));
  INV_X1    g373(.A(new_n563), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT33), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G15gat), .B(G43gat), .Z(new_n579));
  XNOR2_X1  g378(.A(G71gat), .B(G99gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n573), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n581), .B1(new_n566), .B2(KEYINPUT33), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n583), .A2(new_n570), .A3(new_n572), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n568), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n582), .A2(new_n584), .A3(new_n568), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(KEYINPUT36), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT36), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n582), .A2(new_n584), .A3(new_n568), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n589), .B1(new_n590), .B2(new_n585), .ZN(new_n591));
  AOI22_X1  g390(.A1(new_n559), .A2(new_n562), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n552), .A2(new_n554), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n590), .A2(new_n585), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n594), .B1(new_n560), .B2(new_n561), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT35), .B1(new_n595), .B2(new_n559), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n532), .B1(new_n536), .B2(new_n387), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n527), .A2(new_n594), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n293), .B1(new_n593), .B2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G99gat), .B(G106gat), .Z(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G85gat), .A2(G92gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT7), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  INV_X1    g405(.A(G85gat), .ZN(new_n607));
  INV_X1    g406(.A(G92gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n603), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n603), .B1(new_n605), .B2(new_n609), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n613), .B1(new_n258), .B2(KEYINPUT17), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n252), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n243), .A2(new_n250), .A3(new_n613), .ZN(new_n616));
  AND2_X1   g415(.A1(G232gat), .A2(G233gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT41), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G190gat), .B(G218gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT98), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n620), .A2(new_n622), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n617), .A2(KEYINPUT41), .ZN(new_n625));
  XOR2_X1   g424(.A(G134gat), .B(G162gat), .Z(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  OR3_X1    g427(.A1(new_n623), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n628), .B1(new_n623), .B2(new_n624), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT96), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G71gat), .B(G78gat), .Z(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(G57gat), .B(G64gat), .Z(new_n637));
  NAND3_X1  g436(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(KEYINPUT9), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n635), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT21), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(G231gat), .A2(G233gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(G127gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n257), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n647), .B1(new_n642), .B2(new_n641), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n646), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G183gat), .B(G211gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT97), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(new_n297), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n651), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n649), .B(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n631), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(G230gat), .A2(G233gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT100), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n641), .B1(new_n611), .B2(new_n612), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT10), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n605), .A2(new_n609), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n602), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n663), .A2(new_n638), .A3(new_n640), .A4(new_n610), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n660), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n664), .A2(new_n661), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n659), .B1(new_n667), .B2(KEYINPUT99), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT99), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n665), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(G120gat), .B(G148gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT101), .ZN(new_n673));
  XNOR2_X1  g472(.A(G176gat), .B(G204gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n664), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n675), .B1(new_n676), .B2(new_n659), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n659), .ZN(new_n679));
  MUX2_X1   g478(.A(new_n676), .B(new_n667), .S(new_n679), .Z(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n675), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n657), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n601), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n557), .A2(new_n558), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g487(.A1(new_n685), .A2(new_n482), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT16), .B(G8gat), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n691), .B(KEYINPUT42), .Z(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(G8gat), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT102), .Z(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(G1325gat));
  AOI21_X1  g494(.A(G15gat), .B1(new_n685), .B2(new_n594), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n696), .B(KEYINPUT103), .Z(new_n697));
  NAND2_X1  g496(.A1(new_n588), .A2(new_n591), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n685), .A2(G15gat), .A3(new_n699), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n697), .A2(new_n700), .ZN(G1326gat));
  NOR2_X1   g500(.A1(new_n684), .A2(new_n527), .ZN(new_n702));
  XOR2_X1   g501(.A(KEYINPUT43), .B(G22gat), .Z(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1327gat));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n287), .A2(new_n289), .A3(new_n283), .ZN(new_n706));
  AOI221_X4 g505(.A(new_n275), .B1(new_n288), .B2(new_n284), .C1(new_n267), .C2(new_n286), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n682), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n655), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n554), .A2(new_n592), .ZN(new_n712));
  AOI22_X1  g511(.A1(new_n484), .A2(new_n487), .B1(new_n525), .B2(new_n526), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n553), .B1(new_n713), .B2(new_n550), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n600), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n631), .ZN(new_n716));
  NAND2_X1  g515(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n719));
  AOI21_X1  g518(.A(new_n719), .B1(new_n715), .B2(new_n716), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n711), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT105), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n723), .B(new_n711), .C1(new_n718), .C2(new_n720), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n686), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n705), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n724), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n631), .B1(new_n593), .B2(new_n600), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n730), .B2(new_n719), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n723), .B1(new_n731), .B2(new_n711), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(KEYINPUT106), .A3(new_n686), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n727), .A2(new_n734), .A3(G29gat), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n631), .A2(new_n710), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n601), .A2(new_n736), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n737), .A2(G29gat), .A3(new_n726), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT45), .Z(new_n739));
  NAND2_X1  g538(.A1(new_n735), .A2(new_n739), .ZN(G1328gat));
  OAI21_X1  g539(.A(G36gat), .B1(new_n725), .B2(new_n486), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n737), .A2(G36gat), .A3(new_n486), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT46), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(G1329gat));
  NAND2_X1  g543(.A1(new_n204), .A2(new_n205), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n721), .B2(new_n698), .ZN(new_n746));
  INV_X1    g545(.A(new_n594), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n737), .A2(new_n747), .A3(new_n745), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n746), .A2(KEYINPUT47), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n733), .A2(new_n699), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n748), .B1(new_n751), .B2(new_n745), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n752), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT48), .ZN(new_n755));
  OAI21_X1  g554(.A(G50gat), .B1(new_n721), .B2(new_n527), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n527), .A2(G50gat), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n601), .A2(new_n736), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n755), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n208), .B1(new_n733), .B2(new_n562), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n758), .A2(new_n762), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n755), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n754), .B(new_n760), .C1(new_n761), .C2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n722), .A2(new_n562), .A3(new_n724), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n765), .B1(new_n767), .B2(G50gat), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT108), .B1(new_n768), .B2(new_n759), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n766), .A2(new_n769), .ZN(G1331gat));
  NOR3_X1   g569(.A1(new_n657), .A2(new_n291), .A3(new_n709), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n715), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n726), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n773), .B(G57gat), .Z(G1332gat));
  XOR2_X1   g573(.A(new_n772), .B(KEYINPUT109), .Z(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(new_n486), .ZN(new_n776));
  NOR2_X1   g575(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n777));
  AND2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n776), .B2(new_n777), .ZN(G1333gat));
  OAI21_X1  g579(.A(G71gat), .B1(new_n775), .B2(new_n698), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n747), .A2(G71gat), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n772), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n783), .B(new_n784), .ZN(G1334gat));
  NOR2_X1   g584(.A1(new_n775), .A2(new_n527), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n786), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g586(.A1(new_n708), .A2(new_n655), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n788), .B(KEYINPUT110), .Z(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n730), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT111), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n715), .A2(new_n716), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n788), .B(KEYINPUT110), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n796), .A3(KEYINPUT51), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n790), .A2(new_n791), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n792), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n799), .A2(new_n607), .A3(new_n686), .A4(new_n682), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n794), .A2(new_n709), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n731), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n686), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n800), .B1(new_n804), .B2(new_n607), .ZN(G1336gat));
  NOR3_X1   g604(.A1(new_n709), .A2(new_n486), .A3(G92gat), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(KEYINPUT112), .ZN(new_n807));
  INV_X1    g606(.A(new_n798), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n790), .A2(new_n791), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT113), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n802), .A2(new_n482), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G92gat), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n814), .B(new_n807), .C1(new_n808), .C2(new_n809), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n811), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT52), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n799), .A2(KEYINPUT114), .A3(new_n806), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT114), .B1(new_n799), .B2(new_n806), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n818), .B(new_n813), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n817), .A2(new_n821), .ZN(G1337gat));
  INV_X1    g621(.A(G99gat), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n799), .A2(new_n823), .A3(new_n594), .A4(new_n682), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n802), .A2(new_n699), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n824), .B1(new_n826), .B2(new_n823), .ZN(G1338gat));
  OR2_X1    g626(.A1(new_n808), .A2(new_n809), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n527), .A2(G106gat), .A3(new_n709), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n802), .A2(new_n562), .ZN(new_n830));
  AOI22_X1  g629(.A1(new_n828), .A2(new_n829), .B1(new_n830), .B2(G106gat), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(G106gat), .ZN(new_n833));
  XNOR2_X1  g632(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n799), .A2(new_n829), .ZN(new_n836));
  OAI22_X1  g635(.A1(new_n831), .A2(new_n832), .B1(new_n835), .B2(new_n836), .ZN(G1339gat));
  NAND2_X1  g636(.A1(new_n683), .A2(new_n708), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n268), .A2(new_n283), .A3(new_n276), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n261), .B1(new_n260), .B2(new_n262), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n272), .A2(new_n273), .A3(new_n271), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n282), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n665), .A2(new_n666), .A3(new_n659), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT54), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n846), .B1(new_n668), .B2(new_n670), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n667), .A2(new_n848), .A3(new_n679), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n675), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n844), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n846), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n850), .B1(new_n671), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT116), .B1(new_n853), .B2(KEYINPUT55), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT116), .ZN(new_n855));
  NOR4_X1   g654(.A1(new_n847), .A2(new_n850), .A3(new_n855), .A4(new_n844), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n678), .B(new_n851), .C1(new_n854), .C2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n716), .A2(new_n843), .A3(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n858), .B1(new_n706), .B2(new_n707), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n839), .A2(new_n682), .A3(new_n842), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n716), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n861), .A2(KEYINPUT117), .A3(new_n863), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n860), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n838), .B1(new_n868), .B2(new_n656), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870));
  INV_X1    g669(.A(new_n595), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n869), .A2(new_n870), .A3(new_n686), .A4(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n857), .B1(new_n285), .B2(new_n290), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n865), .B1(new_n873), .B2(new_n862), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n867), .A2(new_n874), .A3(new_n631), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n656), .B1(new_n875), .B2(new_n859), .ZN(new_n876));
  INV_X1    g675(.A(new_n838), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n686), .B(new_n871), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT118), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n872), .A2(new_n879), .A3(new_n486), .A4(new_n291), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n324), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n869), .A2(new_n686), .A3(new_n486), .A4(new_n871), .ZN(new_n882));
  OR3_X1    g681(.A1(new_n882), .A2(new_n324), .A3(new_n293), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n881), .A2(new_n883), .A3(KEYINPUT119), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1340gat));
  NOR3_X1   g687(.A1(new_n882), .A2(new_n325), .A3(new_n709), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n872), .A2(new_n879), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n486), .A3(new_n682), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n889), .B1(new_n891), .B2(new_n325), .ZN(G1341gat));
  NOR3_X1   g691(.A1(new_n882), .A2(new_n331), .A3(new_n655), .ZN(new_n893));
  AND4_X1   g692(.A1(new_n486), .A2(new_n872), .A3(new_n656), .A4(new_n879), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n894), .A2(KEYINPUT120), .ZN(new_n895));
  AOI21_X1  g694(.A(G127gat), .B1(new_n894), .B2(KEYINPUT120), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(G1342gat));
  NOR3_X1   g696(.A1(new_n631), .A2(G134gat), .A3(new_n482), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n872), .A2(new_n879), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT56), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n872), .A2(new_n879), .A3(new_n901), .A4(new_n898), .ZN(new_n902));
  OAI21_X1  g701(.A(G134gat), .B1(new_n882), .B2(new_n631), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n900), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n900), .A2(KEYINPUT121), .A3(new_n902), .A4(new_n903), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1343gat));
  NOR2_X1   g707(.A1(new_n699), .A2(new_n527), .ZN(new_n909));
  AND4_X1   g708(.A1(new_n686), .A2(new_n869), .A3(new_n486), .A4(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n293), .A2(G141gat), .ZN(new_n911));
  AOI21_X1  g710(.A(KEYINPUT58), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n699), .A2(new_n726), .A3(new_n482), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n291), .A2(new_n292), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n671), .A2(new_n852), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n917));
  INV_X1    g716(.A(new_n850), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT122), .B1(new_n847), .B2(new_n850), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n919), .A2(new_n920), .A3(new_n844), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n921), .B(new_n678), .C1(new_n854), .C2(new_n856), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT123), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n916), .A2(KEYINPUT55), .A3(new_n918), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n855), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n853), .A2(KEYINPUT116), .A3(KEYINPUT55), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n927), .A2(new_n928), .A3(new_n678), .A4(new_n921), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n923), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT95), .B1(new_n285), .B2(new_n290), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n915), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n631), .B1(new_n932), .B2(new_n862), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n656), .B1(new_n933), .B2(new_n859), .ZN(new_n934));
  OAI211_X1 g733(.A(KEYINPUT57), .B(new_n562), .C1(new_n934), .C2(new_n877), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n562), .B1(new_n876), .B2(new_n877), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT57), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI211_X1 g737(.A(new_n293), .B(new_n914), .C1(new_n935), .C2(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n912), .B1(new_n939), .B2(new_n301), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n876), .A2(new_n877), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n941), .A2(new_n726), .ZN(new_n942));
  AND4_X1   g741(.A1(new_n486), .A2(new_n942), .A3(new_n909), .A4(new_n911), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n914), .B1(new_n935), .B2(new_n938), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n291), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n943), .B1(new_n945), .B2(G141gat), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT58), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n940), .B1(new_n946), .B2(new_n947), .ZN(G1344gat));
  NAND3_X1  g747(.A1(new_n910), .A2(new_n303), .A3(new_n682), .ZN(new_n949));
  AOI211_X1 g748(.A(KEYINPUT59), .B(new_n303), .C1(new_n944), .C2(new_n682), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT59), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n293), .A2(new_n683), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT124), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n937), .B(new_n562), .C1(new_n953), .C2(new_n934), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n936), .A2(KEYINPUT57), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n954), .A2(new_n682), .A3(new_n913), .A4(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n951), .B1(new_n956), .B2(G148gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n949), .B1(new_n950), .B2(new_n957), .ZN(G1345gat));
  NAND3_X1  g757(.A1(new_n910), .A2(new_n297), .A3(new_n656), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n944), .A2(new_n656), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n960), .B2(new_n297), .ZN(G1346gat));
  NOR3_X1   g760(.A1(new_n631), .A2(G162gat), .A3(new_n482), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n942), .A2(new_n909), .A3(new_n962), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n944), .A2(new_n716), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n963), .B1(new_n964), .B2(new_n298), .ZN(G1347gat));
  NOR2_X1   g764(.A1(new_n686), .A2(new_n486), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n871), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n941), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(G169gat), .B1(new_n968), .B2(new_n291), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n293), .A2(new_n409), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n969), .B1(new_n968), .B2(new_n970), .ZN(G1348gat));
  NAND2_X1  g770(.A1(new_n968), .A2(new_n682), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g772(.A1(new_n968), .A2(new_n656), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n974), .A2(new_n430), .ZN(new_n975));
  NAND2_X1  g774(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n974), .A2(new_n425), .ZN(new_n977));
  AND3_X1   g776(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n976), .B1(new_n975), .B2(new_n977), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n978), .A2(new_n979), .ZN(G1350gat));
  NAND2_X1  g779(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n981));
  XNOR2_X1  g780(.A(KEYINPUT61), .B(G190gat), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n968), .A2(new_n716), .ZN(new_n983));
  MUX2_X1   g782(.A(new_n981), .B(new_n982), .S(new_n983), .Z(G1351gat));
  INV_X1    g783(.A(new_n936), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n966), .A2(new_n698), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g787(.A(G197gat), .B1(new_n988), .B2(new_n291), .ZN(new_n989));
  AND2_X1   g788(.A1(new_n954), .A2(new_n955), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n990), .A2(new_n986), .ZN(new_n991));
  INV_X1    g790(.A(G197gat), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n293), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n989), .B1(new_n991), .B2(new_n993), .ZN(G1352gat));
  INV_X1    g793(.A(G204gat), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n682), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g795(.A(KEYINPUT62), .B1(new_n987), .B2(new_n996), .ZN(new_n997));
  OR3_X1    g796(.A1(new_n987), .A2(KEYINPUT62), .A3(new_n996), .ZN(new_n998));
  AND3_X1   g797(.A1(new_n990), .A2(new_n682), .A3(new_n986), .ZN(new_n999));
  OAI211_X1 g798(.A(new_n997), .B(new_n998), .C1(new_n999), .C2(new_n995), .ZN(G1353gat));
  NAND4_X1  g799(.A1(new_n954), .A2(new_n656), .A3(new_n955), .A4(new_n986), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1001), .A2(G211gat), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1002), .A2(KEYINPUT63), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT63), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n1001), .A2(new_n1004), .A3(G211gat), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n656), .A2(new_n455), .ZN(new_n1006));
  NOR2_X1   g805(.A1(new_n987), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n1007), .A2(KEYINPUT126), .ZN(new_n1008));
  AND2_X1   g807(.A1(new_n1007), .A2(KEYINPUT126), .ZN(new_n1009));
  OAI211_X1 g808(.A(new_n1003), .B(new_n1005), .C1(new_n1008), .C2(new_n1009), .ZN(G1354gat));
  OR2_X1    g809(.A1(new_n449), .A2(new_n450), .ZN(new_n1011));
  NAND4_X1  g810(.A1(new_n990), .A2(new_n1011), .A3(new_n716), .A4(new_n986), .ZN(new_n1012));
  OAI211_X1 g811(.A(KEYINPUT127), .B(new_n457), .C1(new_n987), .C2(new_n631), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n457), .B1(new_n987), .B2(new_n631), .ZN(new_n1014));
  INV_X1    g813(.A(KEYINPUT127), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AND3_X1   g815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1016), .ZN(G1355gat));
endmodule


