//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n576, new_n577, new_n578, new_n579,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n593, new_n594, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n632,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  OR2_X1    g040(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(KEYINPUT3), .A3(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n468), .A2(G137), .A3(new_n471), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n465), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT70), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n465), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n471), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n481));
  INV_X1    g056(.A(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT3), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n473), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n481), .B1(new_n485), .B2(G125), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n473), .A2(new_n483), .A3(new_n481), .A4(G125), .ZN(new_n487));
  INV_X1    g062(.A(G113), .ZN(new_n488));
  OR3_X1    g063(.A1(new_n488), .A2(new_n482), .A3(KEYINPUT68), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT68), .B1(new_n488), .B2(new_n482), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n480), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n479), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G160));
  OAI221_X1 g069(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n471), .C2(G112), .ZN(new_n495));
  XOR2_X1   g070(.A(new_n495), .B(KEYINPUT71), .Z(new_n496));
  INV_X1    g071(.A(G124), .ZN(new_n497));
  INV_X1    g072(.A(new_n473), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(new_n480), .ZN(new_n500));
  INV_X1    g075(.A(G136), .ZN(new_n501));
  INV_X1    g076(.A(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  OAI221_X1 g078(.A(new_n496), .B1(new_n497), .B2(new_n500), .C1(new_n501), .C2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G162));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(G114), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(G2105), .ZN(new_n508));
  AND2_X1   g083(.A1(G126), .A2(G2105), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n468), .A2(new_n473), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT72), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n468), .A2(new_n512), .A3(new_n473), .A4(new_n509), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n508), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n468), .A2(new_n473), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n471), .A2(G138), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT4), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT4), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n485), .A2(new_n518), .A3(G138), .A4(new_n471), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n514), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(G164));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  AND2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G543), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT5), .B(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G88), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n523), .A2(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n528), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G651), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n531), .A2(new_n534), .ZN(G303));
  INV_X1    g110(.A(G303), .ZN(G166));
  XOR2_X1   g111(.A(KEYINPUT5), .B(G543), .Z(new_n537));
  NOR2_X1   g112(.A1(new_n524), .A2(new_n525), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G89), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n540), .A2(KEYINPUT74), .A3(new_n542), .ZN(new_n546));
  INV_X1    g121(.A(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n538), .A2(new_n547), .ZN(new_n548));
  AND2_X1   g123(.A1(G63), .A2(G651), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n548), .A2(G51), .B1(new_n528), .B2(new_n549), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(KEYINPUT73), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(KEYINPUT73), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n545), .A2(new_n546), .B1(new_n551), .B2(new_n552), .ZN(G168));
  NAND2_X1  g128(.A1(new_n539), .A2(G90), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n548), .A2(G52), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n533), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT75), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n558), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n560), .A2(new_n561), .A3(new_n555), .A4(new_n554), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G171));
  AOI22_X1  g138(.A1(new_n528), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n533), .ZN(new_n565));
  INV_X1    g140(.A(G43), .ZN(new_n566));
  INV_X1    g141(.A(G81), .ZN(new_n567));
  OAI22_X1  g142(.A1(new_n566), .A2(new_n527), .B1(new_n529), .B2(new_n567), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n568), .A2(KEYINPUT76), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n568), .A2(KEYINPUT76), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n565), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G860), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT77), .ZN(G153));
  NAND4_X1  g149(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XNOR2_X1  g150(.A(KEYINPUT78), .B(KEYINPUT8), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT79), .ZN(new_n577));
  NAND2_X1  g152(.A1(G1), .A2(G3), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(G319), .A2(G483), .A3(G661), .A4(new_n579), .ZN(G188));
  INV_X1    g155(.A(G53), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT9), .B1(new_n527), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT9), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n548), .A2(new_n583), .A3(G53), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  OR3_X1    g160(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT80), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n529), .A2(KEYINPUT80), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n586), .A2(new_n587), .A3(G91), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n528), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(new_n533), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n585), .A2(new_n588), .A3(new_n590), .ZN(G299));
  INV_X1    g166(.A(G171), .ZN(G301));
  NAND2_X1  g167(.A1(new_n545), .A2(new_n546), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n551), .A2(new_n552), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(G286));
  NAND3_X1  g170(.A1(new_n586), .A2(new_n587), .A3(G87), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n528), .A2(G74), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(new_n548), .B2(G49), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(G288));
  NAND3_X1  g176(.A1(new_n586), .A2(new_n587), .A3(G86), .ZN(new_n602));
  NAND2_X1  g177(.A1(G73), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G61), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n537), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(G651), .B1(new_n548), .B2(G48), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n602), .A2(new_n606), .ZN(G305));
  NAND2_X1  g182(.A1(new_n539), .A2(G85), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT82), .B(G47), .ZN(new_n610));
  OAI221_X1 g185(.A(new_n608), .B1(new_n533), .B2(new_n609), .C1(new_n527), .C2(new_n610), .ZN(G290));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NOR2_X1   g187(.A1(G301), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n586), .A2(new_n587), .A3(G92), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT10), .A4(G92), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n537), .B2(new_n620), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n621), .A2(G651), .B1(new_n548), .B2(G54), .ZN(new_n622));
  AND3_X1   g197(.A1(new_n618), .A2(KEYINPUT83), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(KEYINPUT83), .B1(new_n618), .B2(new_n622), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n613), .B1(new_n626), .B2(new_n612), .ZN(G284));
  AOI21_X1  g202(.A(new_n613), .B1(new_n626), .B2(new_n612), .ZN(G321));
  NAND2_X1  g203(.A1(G299), .A2(new_n612), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G168), .B2(new_n612), .ZN(G297));
  OAI21_X1  g205(.A(new_n629), .B1(G168), .B2(new_n612), .ZN(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n626), .B1(new_n632), .B2(G860), .ZN(G148));
  OAI21_X1  g208(.A(KEYINPUT84), .B1(new_n572), .B2(G868), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n626), .A2(new_n632), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G868), .ZN(new_n636));
  MUX2_X1   g211(.A(KEYINPUT84), .B(new_n634), .S(new_n636), .Z(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g213(.A(new_n500), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G123), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT85), .ZN(new_n641));
  OAI221_X1 g216(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n471), .C2(G111), .ZN(new_n642));
  INV_X1    g217(.A(G135), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n642), .B1(new_n503), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n646), .A2(G2096), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(G2096), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n464), .A2(new_n485), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT12), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT13), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2100), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n647), .A2(new_n648), .A3(new_n652), .ZN(G156));
  XOR2_X1   g228(.A(KEYINPUT15), .B(G2435), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2438), .ZN(new_n655));
  XOR2_X1   g230(.A(G2427), .B(G2430), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT86), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(KEYINPUT14), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2451), .B(G2454), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n660), .B(new_n664), .Z(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(G14), .A3(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G401));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2072), .B(G2078), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT18), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n673), .A2(new_n674), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n678), .A2(new_n672), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT87), .B(KEYINPUT17), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n674), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n673), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n679), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n681), .A2(new_n682), .A3(new_n672), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n677), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(G2096), .Z(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT88), .B(G2100), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G227));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1971), .B(G1976), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT19), .ZN(new_n695));
  XOR2_X1   g270(.A(G1956), .B(G2474), .Z(new_n696));
  XOR2_X1   g271(.A(G1961), .B(G1966), .Z(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT20), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n696), .A2(new_n697), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT89), .ZN(new_n703));
  OR3_X1    g278(.A1(new_n695), .A2(new_n698), .A3(new_n701), .ZN(new_n704));
  AND3_X1   g279(.A1(new_n700), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(G1991), .B(G1996), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n707), .A2(new_n708), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n693), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n711), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n713), .A2(new_n692), .A3(new_n709), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(G229));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G23), .ZN(new_n718));
  INV_X1    g293(.A(new_n599), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(new_n717), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT33), .B(G1976), .Z(new_n721));
  XOR2_X1   g296(.A(new_n720), .B(new_n721), .Z(new_n722));
  XOR2_X1   g297(.A(KEYINPUT91), .B(G16), .Z(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n724), .A2(G22), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G166), .B2(new_n724), .ZN(new_n726));
  INV_X1    g301(.A(G1971), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  MUX2_X1   g303(.A(G6), .B(G305), .S(G16), .Z(new_n729));
  XOR2_X1   g304(.A(KEYINPUT32), .B(G1981), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  AND3_X1   g306(.A1(new_n722), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT34), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT92), .Z(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G25), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT90), .Z(new_n738));
  OAI221_X1 g313(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n471), .C2(G107), .ZN(new_n739));
  INV_X1    g314(.A(G131), .ZN(new_n740));
  INV_X1    g315(.A(G119), .ZN(new_n741));
  OAI221_X1 g316(.A(new_n739), .B1(new_n503), .B2(new_n740), .C1(new_n741), .C2(new_n500), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n738), .B1(new_n742), .B2(G29), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT35), .B(G1991), .Z(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  MUX2_X1   g320(.A(G24), .B(G290), .S(new_n724), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1986), .ZN(new_n747));
  AOI211_X1 g322(.A(new_n745), .B(new_n747), .C1(new_n732), .C2(new_n733), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n735), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT36), .ZN(new_n750));
  NOR2_X1   g325(.A1(G29), .A2(G35), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G162), .B2(G29), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT29), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G2090), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n736), .A2(G27), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G164), .B2(new_n736), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT98), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G2078), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n723), .A2(G19), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT94), .Z(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n572), .B2(new_n723), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1341), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT26), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n464), .A2(G105), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G141), .ZN(new_n768));
  INV_X1    g343(.A(G129), .ZN(new_n769));
  OAI221_X1 g344(.A(new_n767), .B1(new_n503), .B2(new_n768), .C1(new_n769), .C2(new_n500), .ZN(new_n770));
  MUX2_X1   g345(.A(G32), .B(new_n770), .S(G29), .Z(new_n771));
  XOR2_X1   g346(.A(KEYINPUT27), .B(G1996), .Z(new_n772));
  NAND2_X1  g347(.A1(new_n717), .A2(G5), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G171), .B2(new_n717), .ZN(new_n774));
  OAI22_X1  g349(.A1(new_n771), .A2(new_n772), .B1(new_n774), .B2(G1961), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n762), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT30), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n777), .A2(G28), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n736), .B1(new_n777), .B2(G28), .ZN(new_n779));
  AND2_X1   g354(.A1(KEYINPUT31), .A2(G11), .ZN(new_n780));
  NOR2_X1   g355(.A1(KEYINPUT31), .A2(G11), .ZN(new_n781));
  OAI22_X1  g356(.A1(new_n778), .A2(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n645), .B2(G29), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT25), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G139), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n485), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n788));
  OAI221_X1 g363(.A(new_n786), .B1(new_n787), .B2(new_n503), .C1(new_n471), .C2(new_n788), .ZN(new_n789));
  MUX2_X1   g364(.A(G33), .B(new_n789), .S(G29), .Z(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G2072), .Z(new_n791));
  AOI22_X1  g366(.A1(new_n771), .A2(new_n772), .B1(new_n774), .B2(G1961), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n776), .A2(new_n783), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  NOR3_X1   g368(.A1(new_n754), .A2(new_n758), .A3(new_n793), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT97), .B(KEYINPUT28), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n736), .A2(G26), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  OAI221_X1 g372(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n471), .C2(G116), .ZN(new_n798));
  INV_X1    g373(.A(G140), .ZN(new_n799));
  INV_X1    g374(.A(G128), .ZN(new_n800));
  OAI221_X1 g375(.A(new_n798), .B1(new_n503), .B2(new_n799), .C1(new_n800), .C2(new_n500), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT95), .ZN(new_n802));
  AND3_X1   g377(.A1(new_n802), .A2(KEYINPUT96), .A3(G29), .ZN(new_n803));
  AOI21_X1  g378(.A(KEYINPUT96), .B1(new_n802), .B2(G29), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n797), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(G2067), .Z(new_n806));
  NOR2_X1   g381(.A1(G4), .A2(G16), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n626), .B2(G16), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT93), .B(G1348), .Z(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n808), .A2(new_n810), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n736), .B1(KEYINPUT24), .B2(G34), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(KEYINPUT24), .B2(G34), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n493), .B2(G29), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G2084), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n723), .A2(G20), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT23), .ZN(new_n818));
  INV_X1    g393(.A(G299), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(new_n717), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(G1956), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n717), .A2(G21), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G168), .B2(new_n717), .ZN(new_n823));
  INV_X1    g398(.A(G1966), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n816), .A2(new_n821), .A3(new_n825), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n811), .A2(new_n812), .A3(new_n826), .ZN(new_n827));
  AND3_X1   g402(.A1(new_n794), .A2(new_n806), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n750), .A2(new_n828), .ZN(G150));
  INV_X1    g404(.A(G150), .ZN(G311));
  NOR2_X1   g405(.A1(new_n625), .A2(new_n632), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G55), .ZN(new_n834));
  INV_X1    g409(.A(G93), .ZN(new_n835));
  OAI22_X1  g410(.A1(new_n834), .A2(new_n527), .B1(new_n529), .B2(new_n835), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n528), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n837), .A2(new_n533), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n571), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n833), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT39), .ZN(new_n843));
  AOI21_X1  g418(.A(G860), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n843), .B2(new_n842), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n840), .A2(G860), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT100), .B(KEYINPUT37), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n845), .A2(new_n848), .ZN(G145));
  XNOR2_X1  g424(.A(new_n504), .B(new_n493), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n646), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT101), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n511), .A2(new_n513), .ZN(new_n853));
  INV_X1    g428(.A(new_n508), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI211_X1 g430(.A(KEYINPUT101), .B(new_n508), .C1(new_n511), .C2(new_n513), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n520), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n802), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n742), .ZN(new_n859));
  OAI221_X1 g434(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n471), .C2(G118), .ZN(new_n860));
  INV_X1    g435(.A(G142), .ZN(new_n861));
  INV_X1    g436(.A(G130), .ZN(new_n862));
  OAI221_X1 g437(.A(new_n860), .B1(new_n503), .B2(new_n861), .C1(new_n862), .C2(new_n500), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT102), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n650), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n789), .B(new_n770), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n859), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n859), .A2(new_n867), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n851), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n859), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n865), .B(new_n866), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n851), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n859), .A2(new_n867), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(G37), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n870), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g454(.A(new_n635), .B(new_n841), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n618), .A2(new_n622), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(G299), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n819), .A2(new_n618), .A3(new_n622), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(KEYINPUT41), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT103), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n883), .A2(new_n888), .A3(new_n884), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n889), .A2(new_n887), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n881), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n885), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n893), .B1(new_n894), .B2(new_n881), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT42), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n893), .B(new_n897), .C1(new_n894), .C2(new_n881), .ZN(new_n898));
  XNOR2_X1  g473(.A(G303), .B(new_n599), .ZN(new_n899));
  XNOR2_X1  g474(.A(G305), .B(G290), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n899), .B(new_n900), .Z(new_n901));
  AND3_X1   g476(.A1(new_n896), .A2(new_n898), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n901), .B1(new_n896), .B2(new_n898), .ZN(new_n903));
  OAI21_X1  g478(.A(G868), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(G868), .B2(new_n839), .ZN(G295));
  OAI21_X1  g480(.A(new_n904), .B1(G868), .B2(new_n839), .ZN(G331));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT106), .B1(G301), .B2(G168), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n909));
  NAND3_X1  g484(.A1(G286), .A2(new_n909), .A3(G171), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT105), .B1(G286), .B2(G171), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n913));
  NAND3_X1  g488(.A1(G301), .A2(G168), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n911), .A2(new_n915), .A3(new_n841), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n841), .B1(new_n911), .B2(new_n915), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n891), .B(new_n890), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n901), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n911), .A2(new_n915), .ZN(new_n920));
  INV_X1    g495(.A(new_n841), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n911), .A2(new_n915), .A3(new_n841), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n894), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n918), .A2(new_n919), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n919), .B1(new_n918), .B2(new_n924), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n927), .A2(G37), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n926), .B1(new_n928), .B2(KEYINPUT107), .ZN(new_n929));
  XNOR2_X1  g504(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n927), .B2(G37), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n922), .A2(new_n923), .B1(new_n889), .B2(new_n886), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n916), .A2(new_n917), .A3(new_n885), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n901), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(new_n925), .A3(new_n877), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n907), .B1(new_n933), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n930), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n918), .A2(new_n924), .ZN(new_n942));
  OAI211_X1 g517(.A(KEYINPUT107), .B(new_n877), .C1(new_n942), .C2(new_n919), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(new_n932), .A3(new_n925), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n941), .B1(new_n944), .B2(new_n940), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n939), .B1(new_n907), .B2(new_n945), .ZN(G397));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n947));
  INV_X1    g522(.A(new_n520), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n512), .B1(new_n499), .B2(new_n509), .ZN(new_n949));
  INV_X1    g524(.A(new_n513), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n854), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT101), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n514), .A2(new_n852), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n948), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n947), .B1(new_n954), .B2(G1384), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n476), .A2(new_n492), .A3(G40), .A4(new_n478), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n802), .B(G2067), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n957), .B1(new_n958), .B2(new_n770), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n959), .B(KEYINPUT124), .Z(new_n960));
  NOR3_X1   g535(.A1(new_n955), .A2(G1996), .A3(new_n956), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT46), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n963), .B(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n957), .A2(G1996), .A3(new_n770), .ZN(new_n966));
  OR2_X1    g541(.A1(new_n966), .A2(KEYINPUT109), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(KEYINPUT109), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n770), .A2(G1996), .ZN(new_n969));
  OR2_X1    g544(.A1(new_n958), .A2(new_n969), .ZN(new_n970));
  AOI22_X1  g545(.A1(new_n967), .A2(new_n968), .B1(new_n970), .B2(new_n957), .ZN(new_n971));
  INV_X1    g546(.A(new_n744), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n742), .A2(new_n972), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n802), .A2(G2067), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n957), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n742), .A2(new_n972), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n957), .B1(new_n977), .B2(new_n973), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n971), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(G290), .A2(G1986), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n957), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT48), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n965), .A2(new_n976), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1384), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT45), .B1(new_n857), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n956), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n947), .A2(G1384), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n987), .B1(G164), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n824), .B1(new_n986), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n857), .A2(new_n992), .A3(new_n985), .ZN(new_n993));
  INV_X1    g568(.A(G2084), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n521), .A2(new_n985), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n956), .B1(new_n995), .B2(KEYINPUT50), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n993), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n991), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(G8), .ZN(new_n999));
  INV_X1    g574(.A(G8), .ZN(new_n1000));
  NOR2_X1   g575(.A1(G168), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT51), .B1(new_n1001), .B2(KEYINPUT116), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1003), .ZN(new_n1005));
  OAI211_X1 g580(.A(G8), .B(new_n1005), .C1(new_n998), .C2(G286), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n998), .A2(new_n1001), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT62), .ZN(new_n1010));
  NAND2_X1  g585(.A1(G303), .A2(G8), .ZN(new_n1011));
  XOR2_X1   g586(.A(new_n1011), .B(KEYINPUT55), .Z(new_n1012));
  NAND2_X1  g587(.A1(new_n995), .A2(new_n947), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n987), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT110), .B1(new_n954), .B2(new_n989), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n857), .A2(new_n1016), .A3(new_n988), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1014), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1018), .A2(G1971), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n993), .A2(new_n996), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1020), .A2(G2090), .ZN(new_n1021));
  OAI211_X1 g596(.A(G8), .B(new_n1012), .C1(new_n1019), .C2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g597(.A(KEYINPUT112), .B(G86), .Z(new_n1023));
  OAI21_X1  g598(.A(new_n606), .B1(new_n529), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(G1981), .ZN(new_n1025));
  INV_X1    g600(.A(G1981), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n602), .A2(new_n1026), .A3(new_n606), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1025), .A2(KEYINPUT49), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT49), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n857), .A2(new_n987), .A3(new_n985), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(G8), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n719), .A2(G1976), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(G8), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT52), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1976), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT52), .B1(G288), .B2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1038), .A2(G8), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT111), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1031), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(new_n1000), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1042), .A2(new_n1043), .A3(new_n1033), .A4(new_n1038), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1036), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n992), .B1(new_n857), .B2(new_n985), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n987), .B1(new_n995), .B2(KEYINPUT50), .ZN(new_n1047));
  OR3_X1    g622(.A1(new_n1046), .A2(new_n1047), .A3(KEYINPUT113), .ZN(new_n1048));
  INV_X1    g623(.A(G2090), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT113), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n956), .B1(new_n995), .B2(new_n947), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n727), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1000), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1022), .B(new_n1045), .C1(new_n1056), .C2(new_n1012), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1004), .A2(new_n1006), .B1(new_n1001), .B2(new_n998), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT62), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G2078), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT53), .B1(new_n1018), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G1961), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1020), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n990), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1067), .A2(G2078), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(new_n955), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(G171), .B1(new_n1063), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT117), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(G171), .C1(new_n1063), .C2(new_n1070), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1010), .A2(new_n1058), .A3(new_n1061), .A4(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT63), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n998), .A2(G8), .A3(G168), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1077), .B1(new_n1057), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(G8), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1012), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1078), .A2(new_n1077), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1082), .A2(new_n1022), .A3(new_n1045), .A4(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1079), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1022), .ZN(new_n1086));
  OR2_X1    g661(.A1(G288), .A2(G1976), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1027), .B1(new_n1087), .B2(new_n1030), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1086), .A2(new_n1045), .B1(new_n1042), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1076), .A2(new_n1085), .A3(new_n1089), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n857), .A2(new_n1016), .A3(new_n988), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1016), .B1(new_n857), .B2(new_n988), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1062), .B(new_n1053), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1067), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT119), .B(G2078), .Z(new_n1095));
  NAND4_X1  g670(.A1(new_n492), .A2(KEYINPUT53), .A3(G40), .A4(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n476), .A2(KEYINPUT118), .A3(new_n478), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT118), .B1(new_n476), .B2(new_n478), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n986), .A2(new_n1100), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1052), .A2(new_n1101), .B1(new_n1020), .B2(new_n1064), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1094), .A2(new_n1102), .A3(G301), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT120), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1094), .A2(new_n1102), .A3(new_n1105), .A4(G301), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1072), .A2(new_n1074), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT56), .B(G2072), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1052), .A2(new_n1053), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT114), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1018), .A2(new_n1115), .A3(new_n1112), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1118), .A2(G1956), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(G299), .B(KEYINPUT57), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1117), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1122), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1124));
  AOI21_X1  g699(.A(G1348), .B1(new_n993), .B2(new_n996), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1031), .A2(G2067), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT115), .ZN(new_n1127));
  OR3_X1    g702(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1127), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1130), .A2(new_n625), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1123), .B1(new_n1124), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT60), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1133), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n626), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1128), .A2(new_n1133), .A3(new_n1129), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1136), .A2(new_n626), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1135), .B1(new_n1137), .B2(new_n1134), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  AOI211_X1 g714(.A(new_n1119), .B(new_n1121), .C1(new_n1114), .C2(new_n1116), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1139), .B1(new_n1124), .B2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT58), .B(G1341), .ZN(new_n1142));
  OAI22_X1  g717(.A1(new_n1054), .A2(G1996), .B1(new_n1041), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n572), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT59), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1119), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1123), .B(KEYINPUT61), .C1(new_n1122), .C2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1138), .A2(new_n1141), .A3(new_n1145), .A4(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1111), .B1(new_n1132), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1100), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n955), .B(new_n1150), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n1065), .ZN(new_n1152));
  OAI21_X1  g727(.A(KEYINPUT121), .B1(new_n1063), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1094), .A2(new_n1102), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1153), .A2(G171), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT122), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1153), .A2(new_n1158), .A3(G171), .A4(new_n1155), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1094), .A2(G301), .A3(new_n1069), .A4(new_n1065), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT54), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(KEYINPUT123), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n1165));
  AOI211_X1 g740(.A(new_n1165), .B(new_n1162), .C1(new_n1157), .C2(new_n1159), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1090), .B1(new_n1149), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(KEYINPUT108), .B1(G290), .B2(G1986), .ZN(new_n1169));
  NAND2_X1  g744(.A1(G290), .A2(G1986), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1169), .B(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n957), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n979), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n984), .B1(new_n1168), .B2(new_n1173), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n1176));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n1177));
  AOI21_X1  g751(.A(new_n1177), .B1(new_n690), .B2(G319), .ZN(new_n1178));
  AOI211_X1 g752(.A(KEYINPUT125), .B(new_n459), .C1(new_n688), .C2(new_n689), .ZN(new_n1179));
  OAI21_X1  g753(.A(new_n670), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n1181));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g756(.A(KEYINPUT126), .B(new_n670), .C1(new_n1178), .C2(new_n1179), .ZN(new_n1183));
  AND2_X1   g757(.A1(new_n715), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g758(.A1(new_n878), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  OAI21_X1  g759(.A(new_n1176), .B1(new_n945), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g760(.A1(new_n1182), .A2(new_n715), .A3(new_n1183), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n873), .A2(new_n875), .ZN(new_n1188));
  AOI21_X1  g762(.A(G37), .B1(new_n1188), .B2(new_n851), .ZN(new_n1189));
  AOI21_X1  g763(.A(new_n1187), .B1(new_n1189), .B2(new_n876), .ZN(new_n1190));
  AOI21_X1  g764(.A(new_n930), .B1(new_n929), .B2(new_n932), .ZN(new_n1191));
  OAI211_X1 g765(.A(new_n1190), .B(KEYINPUT127), .C1(new_n1191), .C2(new_n941), .ZN(new_n1192));
  AND2_X1   g766(.A1(new_n1186), .A2(new_n1192), .ZN(G308));
  NAND2_X1  g767(.A1(new_n1186), .A2(new_n1192), .ZN(G225));
endmodule


