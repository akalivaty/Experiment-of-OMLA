

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795;

  OR2_X1 U381 ( .A1(n373), .A2(n369), .ZN(n622) );
  XNOR2_X1 U382 ( .A(n579), .B(n425), .ZN(n746) );
  NOR2_X1 U383 ( .A1(n746), .A2(n580), .ZN(n581) );
  INV_X1 U384 ( .A(G953), .ZN(n782) );
  NAND2_X2 U385 ( .A1(n709), .A2(n661), .ZN(n379) );
  XNOR2_X2 U386 ( .A(n622), .B(KEYINPUT1), .ZN(n574) );
  AND2_X2 U387 ( .A1(n701), .A2(n573), .ZN(n596) );
  AND2_X2 U388 ( .A1(n419), .A2(n361), .ZN(n414) );
  NAND2_X2 U389 ( .A1(n439), .A2(n654), .ZN(n444) );
  BUF_X2 U390 ( .A(n765), .Z(n766) );
  NOR2_X1 U391 ( .A1(G953), .A2(G237), .ZN(n502) );
  INV_X1 U392 ( .A(n379), .ZN(n662) );
  NAND2_X1 U393 ( .A1(n403), .A2(n402), .ZN(n401) );
  NAND2_X1 U394 ( .A1(n653), .A2(n651), .ZN(n781) );
  XNOR2_X1 U395 ( .A(n779), .B(n460), .ZN(n493) );
  XNOR2_X1 U396 ( .A(KEYINPUT69), .B(KEYINPUT4), .ZN(n458) );
  XNOR2_X1 U397 ( .A(KEYINPUT67), .B(G101), .ZN(n459) );
  NAND2_X2 U398 ( .A1(n395), .A2(n393), .ZN(n694) );
  AND2_X2 U399 ( .A1(n376), .A2(n378), .ZN(n395) );
  NAND2_X1 U400 ( .A1(n394), .A2(n662), .ZN(n393) );
  NAND2_X1 U401 ( .A1(n377), .A2(n366), .ZN(n376) );
  NAND2_X1 U402 ( .A1(n379), .A2(KEYINPUT65), .ZN(n378) );
  NAND2_X1 U403 ( .A1(n401), .A2(n400), .ZN(n377) );
  INV_X1 U404 ( .A(n781), .ZN(n400) );
  NAND2_X1 U405 ( .A1(n410), .A2(n362), .ZN(n398) );
  OR2_X1 U406 ( .A1(n582), .A2(n535), .ZN(n734) );
  XNOR2_X1 U407 ( .A(n521), .B(n368), .ZN(n779) );
  XNOR2_X1 U408 ( .A(n388), .B(n457), .ZN(n521) );
  XNOR2_X1 U409 ( .A(KEYINPUT88), .B(G110), .ZN(n428) );
  XNOR2_X1 U410 ( .A(G107), .B(G104), .ZN(n429) );
  XNOR2_X1 U411 ( .A(G116), .B(KEYINPUT3), .ZN(n384) );
  NOR2_X1 U412 ( .A1(n568), .A2(n567), .ZN(n591) );
  INV_X1 U413 ( .A(G237), .ZN(n440) );
  XNOR2_X1 U414 ( .A(KEYINPUT15), .B(G902), .ZN(n654) );
  XNOR2_X1 U415 ( .A(n458), .B(G137), .ZN(n368) );
  AND2_X1 U416 ( .A1(n720), .A2(n721), .ZN(n715) );
  XNOR2_X1 U417 ( .A(KEYINPUT86), .B(KEYINPUT0), .ZN(n456) );
  NAND2_X1 U418 ( .A1(n731), .A2(n421), .ZN(n420) );
  INV_X1 U419 ( .A(n447), .ZN(n421) );
  NOR2_X2 U420 ( .A1(n415), .A2(n414), .ZN(n413) );
  NAND2_X1 U421 ( .A1(n407), .A2(n404), .ZN(n415) );
  AND2_X1 U422 ( .A1(n405), .A2(n416), .ZN(n404) );
  NAND2_X1 U423 ( .A1(n389), .A2(KEYINPUT79), .ZN(n402) );
  NOR2_X1 U424 ( .A1(n781), .A2(KEYINPUT65), .ZN(n392) );
  XNOR2_X1 U425 ( .A(n646), .B(KEYINPUT70), .ZN(n647) );
  NOR2_X1 U426 ( .A1(n386), .A2(n385), .ZN(n648) );
  NOR2_X1 U427 ( .A1(n611), .A2(n546), .ZN(n620) );
  NAND2_X1 U428 ( .A1(n375), .A2(n374), .ZN(n373) );
  XNOR2_X1 U429 ( .A(G113), .B(KEYINPUT72), .ZN(n426) );
  XNOR2_X1 U430 ( .A(n482), .B(n481), .ZN(n720) );
  NAND2_X1 U431 ( .A1(n683), .A2(n371), .ZN(n482) );
  BUF_X2 U432 ( .A(n574), .Z(n712) );
  INV_X1 U433 ( .A(n559), .ZN(n380) );
  NAND2_X1 U434 ( .A1(n361), .A2(n406), .ZN(n405) );
  INV_X1 U435 ( .A(n423), .ZN(n406) );
  NAND2_X1 U436 ( .A1(n417), .A2(n456), .ZN(n416) );
  INV_X1 U437 ( .A(n455), .ZN(n417) );
  INV_X1 U438 ( .A(KEYINPUT79), .ZN(n367) );
  NAND2_X1 U439 ( .A1(G237), .A2(G234), .ZN(n448) );
  XNOR2_X1 U440 ( .A(n638), .B(n637), .ZN(n385) );
  XNOR2_X1 U441 ( .A(KEYINPUT80), .B(KEYINPUT46), .ZN(n637) );
  NOR2_X1 U442 ( .A1(n645), .A2(n639), .ZN(n387) );
  INV_X1 U443 ( .A(KEYINPUT68), .ZN(n594) );
  NAND2_X1 U444 ( .A1(n412), .A2(n411), .ZN(n410) );
  NAND2_X1 U445 ( .A1(n372), .A2(n371), .ZN(n370) );
  XNOR2_X1 U446 ( .A(G122), .B(G104), .ZN(n496) );
  XOR2_X1 U447 ( .A(KEYINPUT96), .B(KEYINPUT12), .Z(n497) );
  XNOR2_X1 U448 ( .A(n499), .B(n498), .ZN(n500) );
  INV_X1 U449 ( .A(KEYINPUT11), .ZN(n498) );
  XNOR2_X1 U450 ( .A(G143), .B(G113), .ZN(n499) );
  XNOR2_X1 U451 ( .A(G146), .B(G125), .ZN(n474) );
  INV_X1 U452 ( .A(n419), .ZN(n412) );
  XNOR2_X1 U453 ( .A(KEYINPUT16), .B(G122), .ZN(n430) );
  XNOR2_X1 U454 ( .A(G140), .B(KEYINPUT92), .ZN(n469) );
  INV_X1 U455 ( .A(G134), .ZN(n457) );
  XNOR2_X1 U456 ( .A(G116), .B(G122), .ZN(n513) );
  NAND2_X1 U457 ( .A1(n391), .A2(n390), .ZN(n394) );
  NAND2_X1 U458 ( .A1(n396), .A2(KEYINPUT2), .ZN(n390) );
  NAND2_X1 U459 ( .A1(n392), .A2(n401), .ZN(n391) );
  AND2_X1 U460 ( .A1(n620), .A2(n609), .ZN(n621) );
  NOR2_X1 U461 ( .A1(n616), .A2(n615), .ZN(n629) );
  XNOR2_X1 U462 ( .A(n493), .B(n464), .ZN(n689) );
  NAND2_X1 U463 ( .A1(n665), .A2(G953), .ZN(n698) );
  XNOR2_X1 U464 ( .A(n382), .B(KEYINPUT31), .ZN(n762) );
  NAND2_X1 U465 ( .A1(n399), .A2(n383), .ZN(n382) );
  INV_X1 U466 ( .A(n727), .ZN(n383) );
  XNOR2_X1 U467 ( .A(n557), .B(n556), .ZN(n568) );
  XNOR2_X1 U468 ( .A(n648), .B(n647), .ZN(n660) );
  AND2_X1 U469 ( .A1(n455), .A2(n418), .ZN(n361) );
  AND2_X1 U470 ( .A1(n536), .A2(n721), .ZN(n362) );
  NOR2_X1 U471 ( .A1(n739), .A2(n746), .ZN(n363) );
  AND2_X1 U472 ( .A1(n765), .A2(n659), .ZN(n364) );
  AND2_X1 U473 ( .A1(n412), .A2(n409), .ZN(n365) );
  INV_X1 U474 ( .A(G902), .ZN(n371) );
  AND2_X1 U475 ( .A1(n704), .A2(KEYINPUT65), .ZN(n366) );
  INV_X1 U476 ( .A(KEYINPUT65), .ZN(n396) );
  NAND2_X1 U477 ( .A1(n766), .A2(n367), .ZN(n403) );
  NAND2_X1 U478 ( .A1(n408), .A2(n361), .ZN(n407) );
  XNOR2_X2 U479 ( .A(G143), .B(G128), .ZN(n388) );
  NOR2_X1 U480 ( .A1(n689), .A2(n370), .ZN(n369) );
  INV_X1 U481 ( .A(n466), .ZN(n372) );
  NAND2_X1 U482 ( .A1(n466), .A2(G902), .ZN(n374) );
  NAND2_X1 U483 ( .A1(n689), .A2(n466), .ZN(n375) );
  NAND2_X1 U484 ( .A1(n364), .A2(n653), .ZN(n709) );
  NAND2_X1 U485 ( .A1(n381), .A2(n380), .ZN(n565) );
  INV_X1 U486 ( .A(n762), .ZN(n381) );
  XNOR2_X1 U487 ( .A(n384), .B(G119), .ZN(n427) );
  NAND2_X1 U488 ( .A1(n387), .A2(n640), .ZN(n386) );
  XNOR2_X1 U489 ( .A(n388), .B(n459), .ZN(n435) );
  NAND2_X1 U490 ( .A1(n765), .A2(n603), .ZN(n389) );
  XNOR2_X2 U491 ( .A(n602), .B(n601), .ZN(n765) );
  NOR2_X2 U492 ( .A1(n398), .A2(n397), .ZN(n537) );
  INV_X1 U493 ( .A(n413), .ZN(n397) );
  NAND2_X1 U494 ( .A1(n413), .A2(n410), .ZN(n580) );
  INV_X1 U495 ( .A(n580), .ZN(n399) );
  XNOR2_X1 U496 ( .A(n477), .B(n476), .ZN(n683) );
  XNOR2_X2 U497 ( .A(n494), .B(G472), .ZN(n609) );
  NOR2_X1 U498 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U499 ( .A1(n424), .A2(n423), .ZN(n422) );
  INV_X1 U500 ( .A(n424), .ZN(n408) );
  INV_X1 U501 ( .A(n422), .ZN(n409) );
  NOR2_X1 U502 ( .A1(n422), .A2(n418), .ZN(n411) );
  INV_X1 U503 ( .A(n456), .ZN(n418) );
  NOR2_X1 U504 ( .A1(n550), .A2(n420), .ZN(n419) );
  NAND2_X1 U505 ( .A1(n446), .A2(n447), .ZN(n423) );
  NAND2_X1 U506 ( .A1(n550), .A2(n447), .ZN(n424) );
  XOR2_X1 U507 ( .A(n578), .B(n577), .Z(n425) );
  XNOR2_X1 U508 ( .A(n566), .B(KEYINPUT105), .ZN(n567) );
  XNOR2_X1 U509 ( .A(n501), .B(n500), .ZN(n504) );
  INV_X1 U510 ( .A(KEYINPUT48), .ZN(n646) );
  INV_X1 U511 ( .A(n617), .ZN(n585) );
  XNOR2_X1 U512 ( .A(n427), .B(n426), .ZN(n491) );
  XNOR2_X1 U513 ( .A(n429), .B(n428), .ZN(n461) );
  XNOR2_X1 U514 ( .A(n461), .B(n430), .ZN(n431) );
  XNOR2_X1 U515 ( .A(n491), .B(n431), .ZN(n772) );
  XNOR2_X1 U516 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n433) );
  NAND2_X1 U517 ( .A1(n782), .A2(G224), .ZN(n432) );
  XNOR2_X1 U518 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U519 ( .A(n435), .B(n434), .ZN(n437) );
  XNOR2_X1 U520 ( .A(n458), .B(n474), .ZN(n436) );
  XNOR2_X1 U521 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U522 ( .A(n772), .B(n438), .ZN(n674) );
  INV_X1 U523 ( .A(n674), .ZN(n439) );
  NAND2_X1 U524 ( .A1(n371), .A2(n440), .ZN(n445) );
  NAND2_X1 U525 ( .A1(n445), .A2(G210), .ZN(n442) );
  INV_X1 U526 ( .A(KEYINPUT89), .ZN(n441) );
  XNOR2_X1 U527 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X2 U528 ( .A(n444), .B(n443), .ZN(n550) );
  NAND2_X1 U529 ( .A1(n445), .A2(G214), .ZN(n731) );
  INV_X1 U530 ( .A(n731), .ZN(n446) );
  XNOR2_X1 U531 ( .A(KEYINPUT66), .B(KEYINPUT19), .ZN(n447) );
  NOR2_X1 U532 ( .A1(G898), .A2(n782), .ZN(n773) );
  XNOR2_X1 U533 ( .A(n448), .B(KEYINPUT14), .ZN(n452) );
  NAND2_X1 U534 ( .A1(n452), .A2(G902), .ZN(n449) );
  XOR2_X1 U535 ( .A(KEYINPUT90), .B(n449), .Z(n542) );
  NAND2_X1 U536 ( .A1(n773), .A2(n542), .ZN(n451) );
  INV_X1 U537 ( .A(KEYINPUT91), .ZN(n450) );
  XNOR2_X1 U538 ( .A(n451), .B(n450), .ZN(n454) );
  NAND2_X1 U539 ( .A1(G952), .A2(n452), .ZN(n744) );
  NOR2_X1 U540 ( .A1(n744), .A2(G953), .ZN(n545) );
  INV_X1 U541 ( .A(n545), .ZN(n453) );
  NAND2_X1 U542 ( .A1(n454), .A2(n453), .ZN(n455) );
  XNOR2_X1 U543 ( .A(n459), .B(G146), .ZN(n460) );
  XNOR2_X1 U544 ( .A(G140), .B(G131), .ZN(n505) );
  NAND2_X1 U545 ( .A1(n782), .A2(G227), .ZN(n462) );
  XNOR2_X1 U546 ( .A(n505), .B(n462), .ZN(n463) );
  XNOR2_X1 U547 ( .A(n461), .B(n463), .ZN(n464) );
  INV_X1 U548 ( .A(KEYINPUT71), .ZN(n465) );
  XNOR2_X1 U549 ( .A(n465), .B(G469), .ZN(n466) );
  XOR2_X1 U550 ( .A(G110), .B(G119), .Z(n468) );
  XNOR2_X1 U551 ( .A(G128), .B(G137), .ZN(n467) );
  XNOR2_X1 U552 ( .A(n468), .B(n467), .ZN(n472) );
  XOR2_X1 U553 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n470) );
  XNOR2_X1 U554 ( .A(n470), .B(n469), .ZN(n471) );
  XOR2_X1 U555 ( .A(n472), .B(n471), .Z(n477) );
  NAND2_X1 U556 ( .A1(G234), .A2(n782), .ZN(n473) );
  XOR2_X1 U557 ( .A(KEYINPUT8), .B(n473), .Z(n519) );
  NAND2_X1 U558 ( .A1(n519), .A2(G221), .ZN(n475) );
  XNOR2_X1 U559 ( .A(n474), .B(KEYINPUT10), .ZN(n506) );
  XNOR2_X1 U560 ( .A(n475), .B(n506), .ZN(n476) );
  NAND2_X1 U561 ( .A1(G234), .A2(n654), .ZN(n478) );
  XNOR2_X1 U562 ( .A(KEYINPUT20), .B(n478), .ZN(n483) );
  NAND2_X1 U563 ( .A1(G217), .A2(n483), .ZN(n480) );
  XNOR2_X1 U564 ( .A(KEYINPUT93), .B(KEYINPUT25), .ZN(n479) );
  XNOR2_X1 U565 ( .A(n480), .B(n479), .ZN(n481) );
  NAND2_X1 U566 ( .A1(n483), .A2(G221), .ZN(n484) );
  XNOR2_X1 U567 ( .A(n484), .B(KEYINPUT21), .ZN(n486) );
  INV_X1 U568 ( .A(KEYINPUT94), .ZN(n485) );
  XNOR2_X1 U569 ( .A(n486), .B(n485), .ZN(n721) );
  NAND2_X1 U570 ( .A1(n622), .A2(n715), .ZN(n614) );
  NAND2_X1 U571 ( .A1(n502), .A2(G210), .ZN(n487) );
  XNOR2_X1 U572 ( .A(n487), .B(KEYINPUT5), .ZN(n489) );
  XNOR2_X1 U573 ( .A(G131), .B(KEYINPUT95), .ZN(n488) );
  XNOR2_X1 U574 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U575 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U576 ( .A(n493), .B(n492), .ZN(n695) );
  OR2_X1 U577 ( .A1(n695), .A2(G902), .ZN(n494) );
  NOR2_X1 U578 ( .A1(n614), .A2(n609), .ZN(n495) );
  AND2_X1 U579 ( .A1(n399), .A2(n495), .ZN(n559) );
  XNOR2_X1 U580 ( .A(n497), .B(n496), .ZN(n501) );
  NAND2_X1 U581 ( .A1(n502), .A2(G214), .ZN(n503) );
  XNOR2_X1 U582 ( .A(n504), .B(n503), .ZN(n507) );
  XNOR2_X1 U583 ( .A(n506), .B(n505), .ZN(n778) );
  XNOR2_X1 U584 ( .A(n507), .B(n778), .ZN(n668) );
  NAND2_X1 U585 ( .A1(n668), .A2(n371), .ZN(n512) );
  XOR2_X1 U586 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n509) );
  XNOR2_X1 U587 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n508) );
  XNOR2_X1 U588 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U589 ( .A(G475), .B(n510), .ZN(n511) );
  XNOR2_X1 U590 ( .A(n512), .B(n511), .ZN(n582) );
  XOR2_X1 U591 ( .A(KEYINPUT100), .B(G107), .Z(n514) );
  XNOR2_X1 U592 ( .A(n514), .B(n513), .ZN(n518) );
  XOR2_X1 U593 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n516) );
  XNOR2_X1 U594 ( .A(KEYINPUT7), .B(KEYINPUT102), .ZN(n515) );
  XNOR2_X1 U595 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U596 ( .A(n518), .B(n517), .Z(n523) );
  NAND2_X1 U597 ( .A1(G217), .A2(n519), .ZN(n520) );
  XNOR2_X1 U598 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U599 ( .A(n523), .B(n522), .ZN(n664) );
  NAND2_X1 U600 ( .A1(n664), .A2(n371), .ZN(n526) );
  INV_X1 U601 ( .A(KEYINPUT103), .ZN(n524) );
  XNOR2_X1 U602 ( .A(n524), .B(G478), .ZN(n525) );
  XNOR2_X1 U603 ( .A(n526), .B(n525), .ZN(n535) );
  INV_X1 U604 ( .A(n535), .ZN(n583) );
  AND2_X1 U605 ( .A1(n582), .A2(n583), .ZN(n757) );
  NAND2_X1 U606 ( .A1(n559), .A2(n757), .ZN(n527) );
  XNOR2_X1 U607 ( .A(n527), .B(G104), .ZN(G6) );
  OR2_X1 U608 ( .A1(n582), .A2(n583), .ZN(n560) );
  INV_X1 U609 ( .A(n560), .ZN(n761) );
  NAND2_X1 U610 ( .A1(n559), .A2(n761), .ZN(n532) );
  XOR2_X1 U611 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n529) );
  XNOR2_X1 U612 ( .A(G107), .B(KEYINPUT113), .ZN(n528) );
  XNOR2_X1 U613 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U614 ( .A(KEYINPUT26), .B(n530), .Z(n531) );
  XNOR2_X1 U615 ( .A(n532), .B(n531), .ZN(G9) );
  AND2_X1 U616 ( .A1(n609), .A2(n715), .ZN(n533) );
  NAND2_X1 U617 ( .A1(n712), .A2(n533), .ZN(n727) );
  NAND2_X1 U618 ( .A1(n762), .A2(n757), .ZN(n534) );
  XNOR2_X1 U619 ( .A(n534), .B(G113), .ZN(G15) );
  INV_X1 U620 ( .A(n734), .ZN(n536) );
  XNOR2_X1 U621 ( .A(n537), .B(KEYINPUT22), .ZN(n553) );
  BUF_X1 U622 ( .A(n553), .Z(n538) );
  INV_X1 U623 ( .A(n538), .ZN(n541) );
  OR2_X1 U624 ( .A1(n609), .A2(n720), .ZN(n539) );
  OR2_X1 U625 ( .A1(n712), .A2(n539), .ZN(n540) );
  OR2_X1 U626 ( .A1(n541), .A2(n540), .ZN(n573) );
  XNOR2_X1 U627 ( .A(n573), .B(G110), .ZN(G12) );
  XNOR2_X1 U628 ( .A(n609), .B(KEYINPUT6), .ZN(n575) );
  NAND2_X1 U629 ( .A1(n542), .A2(G953), .ZN(n543) );
  NOR2_X1 U630 ( .A1(G900), .A2(n543), .ZN(n544) );
  NOR2_X1 U631 ( .A1(n545), .A2(n544), .ZN(n611) );
  INV_X1 U632 ( .A(n720), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n721), .A2(n569), .ZN(n546) );
  AND2_X1 U634 ( .A1(n757), .A2(n620), .ZN(n547) );
  NAND2_X1 U635 ( .A1(n731), .A2(n547), .ZN(n548) );
  OR2_X1 U636 ( .A1(n575), .A2(n548), .ZN(n604) );
  OR2_X1 U637 ( .A1(n604), .A2(n712), .ZN(n549) );
  XNOR2_X1 U638 ( .A(n549), .B(KEYINPUT43), .ZN(n552) );
  BUF_X1 U639 ( .A(n550), .Z(n551) );
  NAND2_X1 U640 ( .A1(n552), .A2(n551), .ZN(n658) );
  XNOR2_X1 U641 ( .A(n658), .B(G140), .ZN(G42) );
  AND2_X2 U642 ( .A1(n553), .A2(n575), .ZN(n571) );
  XNOR2_X1 U643 ( .A(n571), .B(KEYINPUT82), .ZN(n555) );
  NOR2_X1 U644 ( .A1(n712), .A2(n569), .ZN(n554) );
  NAND2_X1 U645 ( .A1(n555), .A2(n554), .ZN(n557) );
  INV_X1 U646 ( .A(KEYINPUT106), .ZN(n556) );
  BUF_X1 U647 ( .A(n568), .Z(n558) );
  XOR2_X1 U648 ( .A(n558), .B(G101), .Z(G3) );
  INV_X1 U649 ( .A(n757), .ZN(n561) );
  NAND2_X1 U650 ( .A1(n561), .A2(n560), .ZN(n563) );
  INV_X1 U651 ( .A(KEYINPUT104), .ZN(n562) );
  XNOR2_X1 U652 ( .A(n563), .B(n562), .ZN(n735) );
  INV_X1 U653 ( .A(n735), .ZN(n564) );
  NAND2_X1 U654 ( .A1(n565), .A2(n564), .ZN(n566) );
  AND2_X1 U655 ( .A1(n712), .A2(n569), .ZN(n570) );
  NAND2_X1 U656 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X2 U657 ( .A(n572), .B(KEYINPUT32), .ZN(n701) );
  NAND2_X1 U658 ( .A1(n574), .A2(n715), .ZN(n576) );
  XNOR2_X1 U659 ( .A(KEYINPUT107), .B(KEYINPUT33), .ZN(n578) );
  INV_X1 U660 ( .A(KEYINPUT87), .ZN(n577) );
  XNOR2_X1 U661 ( .A(n581), .B(KEYINPUT34), .ZN(n586) );
  INV_X1 U662 ( .A(n582), .ZN(n584) );
  OR2_X1 U663 ( .A1(n584), .A2(n583), .ZN(n617) );
  NAND2_X1 U664 ( .A1(n586), .A2(n585), .ZN(n588) );
  XNOR2_X1 U665 ( .A(KEYINPUT73), .B(KEYINPUT35), .ZN(n587) );
  XNOR2_X2 U666 ( .A(n588), .B(n587), .ZN(n702) );
  NAND2_X1 U667 ( .A1(n596), .A2(n702), .ZN(n589) );
  NAND2_X1 U668 ( .A1(n589), .A2(KEYINPUT44), .ZN(n590) );
  NAND2_X1 U669 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U670 ( .A(n592), .B(KEYINPUT83), .ZN(n600) );
  INV_X1 U671 ( .A(KEYINPUT44), .ZN(n593) );
  NAND2_X1 U672 ( .A1(n702), .A2(n593), .ZN(n595) );
  XNOR2_X1 U673 ( .A(n595), .B(n594), .ZN(n598) );
  XNOR2_X1 U674 ( .A(n596), .B(KEYINPUT84), .ZN(n597) );
  NAND2_X1 U675 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U676 ( .A1(n600), .A2(n599), .ZN(n602) );
  XNOR2_X1 U677 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n601) );
  INV_X1 U678 ( .A(n654), .ZN(n603) );
  INV_X1 U679 ( .A(n765), .ZN(n703) );
  NOR2_X1 U680 ( .A1(n604), .A2(n551), .ZN(n605) );
  XNOR2_X1 U681 ( .A(n605), .B(KEYINPUT36), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n606), .A2(n712), .ZN(n607) );
  XNOR2_X1 U683 ( .A(n607), .B(KEYINPUT111), .ZN(n789) );
  NOR2_X1 U684 ( .A1(KEYINPUT76), .A2(n735), .ZN(n608) );
  NOR2_X1 U685 ( .A1(n789), .A2(n608), .ZN(n640) );
  NAND2_X1 U686 ( .A1(n609), .A2(n731), .ZN(n610) );
  XOR2_X1 U687 ( .A(n610), .B(KEYINPUT30), .Z(n613) );
  INV_X1 U688 ( .A(n611), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(n616) );
  XNOR2_X1 U690 ( .A(KEYINPUT108), .B(n614), .ZN(n615) );
  NOR2_X1 U691 ( .A1(n617), .A2(n551), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n629), .A2(n618), .ZN(n619) );
  XNOR2_X1 U693 ( .A(KEYINPUT109), .B(n619), .ZN(n791) );
  XNOR2_X1 U694 ( .A(KEYINPUT77), .B(n791), .ZN(n628) );
  XNOR2_X1 U695 ( .A(n621), .B(KEYINPUT28), .ZN(n623) );
  NAND2_X1 U696 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U697 ( .A(n624), .B(KEYINPUT110), .ZN(n634) );
  OR2_X1 U698 ( .A1(n634), .A2(n365), .ZN(n641) );
  INV_X1 U699 ( .A(n641), .ZN(n758) );
  NAND2_X1 U700 ( .A1(n735), .A2(KEYINPUT76), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n758), .A2(n625), .ZN(n626) );
  NAND2_X1 U702 ( .A1(KEYINPUT47), .A2(n626), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n639) );
  XNOR2_X1 U704 ( .A(n551), .B(KEYINPUT38), .ZN(n732) );
  NAND2_X1 U705 ( .A1(n629), .A2(n732), .ZN(n631) );
  XOR2_X1 U706 ( .A(KEYINPUT81), .B(KEYINPUT39), .Z(n630) );
  XNOR2_X1 U707 ( .A(n631), .B(n630), .ZN(n649) );
  NAND2_X1 U708 ( .A1(n649), .A2(n757), .ZN(n632) );
  XNOR2_X1 U709 ( .A(KEYINPUT40), .B(n632), .ZN(n792) );
  INV_X1 U710 ( .A(KEYINPUT42), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n732), .A2(n731), .ZN(n736) );
  NOR2_X1 U712 ( .A1(n734), .A2(n736), .ZN(n633) );
  XNOR2_X1 U713 ( .A(n633), .B(KEYINPUT41), .ZN(n711) );
  NOR2_X1 U714 ( .A1(n634), .A2(n711), .ZN(n635) );
  XNOR2_X1 U715 ( .A(n636), .B(n635), .ZN(n795) );
  NAND2_X1 U716 ( .A1(n792), .A2(n795), .ZN(n638) );
  INV_X1 U717 ( .A(KEYINPUT76), .ZN(n643) );
  NOR2_X1 U718 ( .A1(n641), .A2(n735), .ZN(n642) );
  NOR2_X1 U719 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U720 ( .A1(KEYINPUT47), .A2(n644), .ZN(n645) );
  INV_X1 U721 ( .A(n660), .ZN(n653) );
  NAND2_X1 U722 ( .A1(n761), .A2(n649), .ZN(n650) );
  XNOR2_X1 U723 ( .A(KEYINPUT112), .B(n650), .ZN(n793) );
  AND2_X1 U724 ( .A1(n793), .A2(n658), .ZN(n651) );
  INV_X1 U725 ( .A(KEYINPUT2), .ZN(n704) );
  AND2_X1 U726 ( .A1(n651), .A2(KEYINPUT79), .ZN(n652) );
  NAND2_X1 U727 ( .A1(n653), .A2(n652), .ZN(n655) );
  NAND2_X1 U728 ( .A1(n655), .A2(n654), .ZN(n661) );
  NAND2_X1 U729 ( .A1(KEYINPUT2), .A2(n793), .ZN(n656) );
  XOR2_X1 U730 ( .A(n656), .B(KEYINPUT74), .Z(n657) );
  AND2_X1 U731 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U732 ( .A1(n694), .A2(G478), .ZN(n663) );
  XOR2_X1 U733 ( .A(n664), .B(n663), .Z(n667) );
  INV_X1 U734 ( .A(G952), .ZN(n665) );
  INV_X1 U735 ( .A(n698), .ZN(n666) );
  NOR2_X1 U736 ( .A1(n667), .A2(n666), .ZN(G63) );
  NAND2_X1 U737 ( .A1(n694), .A2(G475), .ZN(n670) );
  XOR2_X1 U738 ( .A(n668), .B(KEYINPUT59), .Z(n669) );
  XNOR2_X1 U739 ( .A(n670), .B(n669), .ZN(n671) );
  NAND2_X1 U740 ( .A1(n671), .A2(n698), .ZN(n673) );
  INV_X1 U741 ( .A(KEYINPUT60), .ZN(n672) );
  XNOR2_X1 U742 ( .A(n673), .B(n672), .ZN(G60) );
  NAND2_X1 U743 ( .A1(n694), .A2(G210), .ZN(n679) );
  BUF_X1 U744 ( .A(n674), .Z(n675) );
  XNOR2_X1 U745 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n676) );
  XOR2_X1 U746 ( .A(n676), .B(KEYINPUT85), .Z(n677) );
  XNOR2_X1 U747 ( .A(n675), .B(n677), .ZN(n678) );
  XNOR2_X1 U748 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U749 ( .A1(n680), .A2(n698), .ZN(n682) );
  XOR2_X1 U750 ( .A(KEYINPUT122), .B(KEYINPUT56), .Z(n681) );
  XNOR2_X1 U751 ( .A(n682), .B(n681), .ZN(G51) );
  NAND2_X1 U752 ( .A1(n694), .A2(G217), .ZN(n684) );
  XNOR2_X1 U753 ( .A(n684), .B(n683), .ZN(n685) );
  NAND2_X1 U754 ( .A1(n685), .A2(n698), .ZN(n687) );
  INV_X1 U755 ( .A(KEYINPUT124), .ZN(n686) );
  XNOR2_X1 U756 ( .A(n687), .B(n686), .ZN(G66) );
  NAND2_X1 U757 ( .A1(n694), .A2(G469), .ZN(n691) );
  XNOR2_X1 U758 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n688) );
  XNOR2_X1 U759 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U760 ( .A(n691), .B(n690), .ZN(n692) );
  NAND2_X1 U761 ( .A1(n692), .A2(n698), .ZN(n693) );
  XNOR2_X1 U762 ( .A(n693), .B(KEYINPUT123), .ZN(G54) );
  NAND2_X1 U763 ( .A1(n694), .A2(G472), .ZN(n697) );
  XOR2_X1 U764 ( .A(KEYINPUT62), .B(n695), .Z(n696) );
  XNOR2_X1 U765 ( .A(n697), .B(n696), .ZN(n699) );
  NAND2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U767 ( .A(n700), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U768 ( .A(n701), .B(G119), .ZN(G21) );
  XNOR2_X1 U769 ( .A(n702), .B(G122), .ZN(G24) );
  NAND2_X1 U770 ( .A1(n781), .A2(n704), .ZN(n707) );
  NAND2_X1 U771 ( .A1(n703), .A2(n704), .ZN(n705) );
  XNOR2_X1 U772 ( .A(n705), .B(KEYINPUT78), .ZN(n706) );
  NAND2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U774 ( .A(n708), .B(KEYINPUT75), .ZN(n710) );
  NAND2_X1 U775 ( .A1(n710), .A2(n709), .ZN(n752) );
  INV_X1 U776 ( .A(n712), .ZN(n717) );
  INV_X1 U777 ( .A(n715), .ZN(n713) );
  NAND2_X1 U778 ( .A1(n717), .A2(n713), .ZN(n714) );
  NAND2_X1 U779 ( .A1(n714), .A2(KEYINPUT50), .ZN(n719) );
  NOR2_X1 U780 ( .A1(n715), .A2(KEYINPUT50), .ZN(n716) );
  NAND2_X1 U781 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U782 ( .A1(n719), .A2(n718), .ZN(n726) );
  NOR2_X1 U783 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U784 ( .A(n722), .B(KEYINPUT49), .ZN(n724) );
  INV_X1 U785 ( .A(n609), .ZN(n723) );
  AND2_X1 U786 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U787 ( .A1(n726), .A2(n725), .ZN(n728) );
  AND2_X1 U788 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U789 ( .A(KEYINPUT51), .B(n729), .Z(n730) );
  NOR2_X1 U790 ( .A1(n711), .A2(n730), .ZN(n740) );
  NOR2_X1 U791 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U792 ( .A1(n734), .A2(n733), .ZN(n738) );
  NOR2_X1 U793 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U794 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U795 ( .A1(n740), .A2(n363), .ZN(n741) );
  XNOR2_X1 U796 ( .A(n741), .B(KEYINPUT52), .ZN(n742) );
  XNOR2_X1 U797 ( .A(KEYINPUT118), .B(n742), .ZN(n743) );
  NOR2_X1 U798 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U799 ( .A(KEYINPUT119), .B(n745), .Z(n748) );
  NOR2_X1 U800 ( .A1(n711), .A2(n746), .ZN(n747) );
  NOR2_X1 U801 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U802 ( .A(n749), .B(KEYINPUT120), .Z(n750) );
  NOR2_X1 U803 ( .A1(n750), .A2(G953), .ZN(n751) );
  NAND2_X1 U804 ( .A1(n752), .A2(n751), .ZN(n754) );
  XNOR2_X1 U805 ( .A(KEYINPUT121), .B(KEYINPUT53), .ZN(n753) );
  XNOR2_X1 U806 ( .A(n754), .B(n753), .ZN(G75) );
  XOR2_X1 U807 ( .A(G128), .B(KEYINPUT29), .Z(n756) );
  NAND2_X1 U808 ( .A1(n758), .A2(n761), .ZN(n755) );
  XNOR2_X1 U809 ( .A(n756), .B(n755), .ZN(G30) );
  XOR2_X1 U810 ( .A(G146), .B(KEYINPUT115), .Z(n760) );
  NAND2_X1 U811 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U812 ( .A(n760), .B(n759), .ZN(G48) );
  NAND2_X1 U813 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U814 ( .A(n763), .B(KEYINPUT116), .ZN(n764) );
  XNOR2_X1 U815 ( .A(G116), .B(n764), .ZN(G18) );
  NAND2_X1 U816 ( .A1(n766), .A2(n782), .ZN(n770) );
  NAND2_X1 U817 ( .A1(G953), .A2(G224), .ZN(n767) );
  XNOR2_X1 U818 ( .A(KEYINPUT61), .B(n767), .ZN(n768) );
  NAND2_X1 U819 ( .A1(n768), .A2(G898), .ZN(n769) );
  NAND2_X1 U820 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U821 ( .A(n771), .B(KEYINPUT125), .ZN(n777) );
  XNOR2_X1 U822 ( .A(n772), .B(G101), .ZN(n774) );
  NOR2_X1 U823 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U824 ( .A(n775), .B(KEYINPUT126), .Z(n776) );
  XNOR2_X1 U825 ( .A(n777), .B(n776), .ZN(G69) );
  XOR2_X1 U826 ( .A(n779), .B(n778), .Z(n784) );
  XOR2_X1 U827 ( .A(KEYINPUT127), .B(n784), .Z(n780) );
  XNOR2_X1 U828 ( .A(n781), .B(n780), .ZN(n783) );
  NAND2_X1 U829 ( .A1(n783), .A2(n782), .ZN(n788) );
  XNOR2_X1 U830 ( .A(n784), .B(G227), .ZN(n785) );
  NAND2_X1 U831 ( .A1(n785), .A2(G900), .ZN(n786) );
  NAND2_X1 U832 ( .A1(n786), .A2(G953), .ZN(n787) );
  NAND2_X1 U833 ( .A1(n788), .A2(n787), .ZN(G72) );
  XNOR2_X1 U834 ( .A(G125), .B(n789), .ZN(n790) );
  XNOR2_X1 U835 ( .A(n790), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U836 ( .A(G143), .B(n791), .Z(G45) );
  XNOR2_X1 U837 ( .A(G131), .B(n792), .ZN(G33) );
  XOR2_X1 U838 ( .A(G134), .B(n793), .Z(n794) );
  XNOR2_X1 U839 ( .A(KEYINPUT117), .B(n794), .ZN(G36) );
  XNOR2_X1 U840 ( .A(G137), .B(n795), .ZN(G39) );
endmodule

