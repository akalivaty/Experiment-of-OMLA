//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT64), .B(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G58), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n206), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n209), .B1(new_n213), .B2(new_n218), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G226), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G58), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  XNOR2_X1  g0044(.A(KEYINPUT3), .B(G33), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n245), .A2(G223), .A3(G1698), .ZN(new_n246));
  INV_X1    g0046(.A(G77), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G222), .ZN(new_n250));
  OAI221_X1 g0050(.A(new_n246), .B1(new_n247), .B2(new_n245), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT69), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT67), .A2(G41), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT67), .A2(G41), .ZN(new_n256));
  NOR3_X1   g0056(.A1(new_n255), .A2(new_n256), .A3(G45), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G274), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n254), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  OR2_X1    g0060(.A1(KEYINPUT67), .A2(G41), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT67), .A2(G41), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n259), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(KEYINPUT69), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  AOI21_X1  g0068(.A(G1), .B1(new_n268), .B2(new_n262), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT68), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(KEYINPUT68), .A2(G33), .A3(G41), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n211), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n269), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G226), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n253), .A2(new_n267), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G169), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT72), .B(G179), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n279), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n258), .A2(G13), .A3(G20), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT71), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n258), .A2(KEYINPUT71), .A3(G13), .A4(G20), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(G50), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n211), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G20), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n286), .B(new_n291), .C1(G1), .C2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n288), .B1(G50), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n210), .A2(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT70), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT70), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n210), .A2(new_n297), .A3(G33), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT8), .B(G58), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n296), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(G20), .A2(G33), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n291), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n294), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n281), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT74), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n308), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n305), .A2(KEYINPUT74), .A3(KEYINPUT9), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n305), .A2(KEYINPUT9), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n278), .A2(G200), .ZN(new_n314));
  INV_X1    g0114(.A(G190), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n278), .A2(new_n315), .ZN(new_n316));
  NOR3_X1   g0116(.A1(new_n313), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT10), .ZN(new_n318));
  AND3_X1   g0118(.A1(new_n312), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n318), .B1(new_n312), .B2(new_n317), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n307), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n260), .A2(new_n266), .B1(new_n276), .B2(G238), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT13), .ZN(new_n323));
  INV_X1    g0123(.A(G33), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT3), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G33), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n325), .A2(new_n327), .A3(G232), .A4(G1698), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n325), .A2(new_n327), .A3(G226), .A4(new_n248), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G33), .A2(G97), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n252), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n322), .A2(new_n323), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n323), .B1(new_n322), .B2(new_n332), .ZN(new_n335));
  OAI21_X1  g0135(.A(G169), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT14), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n276), .A2(G238), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n267), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n332), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT13), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n333), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n343), .A2(KEYINPUT14), .A3(G169), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n342), .A2(G179), .A3(new_n333), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT76), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n342), .A2(KEYINPUT76), .A3(G179), .A4(new_n333), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n296), .A2(G77), .A3(new_n298), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n302), .A2(G50), .B1(G20), .B2(new_n215), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n291), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT11), .ZN(new_n355));
  INV_X1    g0155(.A(new_n293), .ZN(new_n356));
  OR3_X1    g0156(.A1(new_n286), .A2(KEYINPUT12), .A3(G68), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT12), .B1(new_n286), .B2(G68), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n356), .A2(G68), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n354), .A2(KEYINPUT11), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT75), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n354), .A2(KEYINPUT11), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT75), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n363), .A2(new_n364), .A3(new_n355), .A4(new_n359), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n351), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G200), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n343), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n342), .A2(new_n315), .A3(new_n333), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n356), .A2(G77), .ZN(new_n375));
  XNOR2_X1  g0175(.A(KEYINPUT15), .B(G87), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n295), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n292), .A2(new_n324), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n247), .A2(new_n210), .B1(new_n299), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n290), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n287), .A2(new_n247), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n375), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G107), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n249), .A2(new_n231), .B1(new_n383), .B2(new_n245), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n245), .A2(G238), .A3(G1698), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n252), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n260), .A2(new_n266), .B1(new_n276), .B2(G244), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G169), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n280), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n386), .A2(new_n391), .A3(new_n387), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n382), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n382), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n388), .A2(G190), .ZN(new_n396));
  AOI21_X1  g0196(.A(G200), .B1(new_n386), .B2(new_n387), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT73), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n394), .A2(KEYINPUT73), .A3(new_n398), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n260), .A2(new_n266), .B1(new_n276), .B2(G232), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n325), .A2(new_n327), .A3(G223), .A4(new_n248), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n325), .A2(new_n327), .A3(G226), .A4(G1698), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G33), .A2(G87), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n252), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n405), .A2(KEYINPUT79), .A3(new_n280), .A4(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT79), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n276), .A2(G232), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n267), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(G169), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n414), .A2(new_n391), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n411), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n286), .A2(new_n299), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n300), .B2(new_n293), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G58), .A2(G68), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(G20), .B1(new_n423), .B2(new_n201), .ZN(new_n424));
  INV_X1    g0224(.A(G159), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT77), .B1(new_n378), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT77), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n302), .A2(new_n427), .A3(G159), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n424), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n292), .A2(KEYINPUT64), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT64), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G20), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT7), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n325), .A2(new_n327), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n215), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n326), .A2(G33), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n324), .A2(KEYINPUT3), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n292), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT7), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n429), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n291), .B1(new_n441), .B2(KEYINPUT16), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT16), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n430), .A2(new_n432), .A3(KEYINPUT7), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT78), .B1(new_n324), .B2(KEYINPUT3), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT78), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(new_n326), .A3(G33), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n447), .A3(new_n325), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n433), .B1(new_n245), .B2(G20), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n215), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n443), .B1(new_n451), .B2(new_n429), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n421), .B1(new_n442), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT18), .B1(new_n418), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n292), .B1(new_n216), .B2(new_n422), .ZN(new_n455));
  NOR4_X1   g0255(.A1(new_n425), .A2(KEYINPUT77), .A3(G20), .A4(G33), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n427), .B1(new_n302), .B2(G159), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n433), .B1(new_n435), .B2(new_n292), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n460));
  OAI21_X1  g0260(.A(G68), .B1(new_n460), .B2(new_n245), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n458), .B(KEYINPUT16), .C1(new_n459), .C2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n452), .A2(new_n290), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n419), .B1(new_n356), .B2(new_n299), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(G169), .B1(new_n405), .B2(new_n410), .ZN(new_n466));
  OAI22_X1  g0266(.A1(new_n466), .A2(new_n412), .B1(new_n391), .B2(new_n414), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT18), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n465), .A2(new_n467), .A3(new_n468), .A4(new_n411), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n264), .A2(KEYINPUT69), .A3(new_n265), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT69), .B1(new_n264), .B2(new_n265), .ZN(new_n471));
  AND3_X1   g0271(.A1(KEYINPUT68), .A2(G33), .A3(G41), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT68), .B1(G33), .B2(G41), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n275), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n269), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI22_X1  g0276(.A1(new_n470), .A2(new_n471), .B1(new_n476), .B2(new_n231), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n409), .A2(new_n252), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n369), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n405), .A2(new_n315), .A3(new_n410), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(new_n463), .A3(new_n464), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT17), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n453), .A2(KEYINPUT17), .A3(new_n481), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n454), .A2(new_n469), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  NOR4_X1   g0286(.A1(new_n321), .A2(new_n374), .A3(new_n404), .A4(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n325), .A2(new_n327), .A3(G244), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n489), .A2(G1698), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n245), .A2(G244), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G283), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n490), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n245), .A2(G250), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n248), .B1(new_n495), .B2(KEYINPUT4), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n252), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(KEYINPUT5), .B1(new_n261), .B2(new_n263), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT5), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n258), .B(G45), .C1(new_n499), .C2(G41), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n474), .B(G257), .C1(new_n498), .C2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n500), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n499), .B1(new_n255), .B2(new_n256), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n474), .A2(new_n502), .A3(new_n503), .A4(G274), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n497), .A2(new_n506), .A3(new_n315), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n488), .A2(new_n489), .B1(G33), .B2(G283), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n489), .B1(new_n245), .B2(G250), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n508), .B(new_n492), .C1(new_n248), .C2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n505), .B1(new_n510), .B2(new_n252), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n507), .B1(new_n511), .B2(G200), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n448), .A2(new_n444), .B1(new_n439), .B2(new_n433), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT81), .B1(new_n513), .B2(new_n383), .ZN(new_n514));
  OR2_X1    g0314(.A1(KEYINPUT80), .A2(G107), .ZN(new_n515));
  NAND2_X1  g0315(.A1(KEYINPUT80), .A2(G107), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(G97), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(new_n383), .A3(KEYINPUT6), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OR2_X1    g0322(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n523), .A2(new_n519), .A3(new_n515), .A4(new_n516), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n430), .A2(new_n432), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n525), .A2(new_n526), .B1(G77), .B2(new_n302), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n449), .A2(new_n450), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT81), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(new_n529), .A3(G107), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n514), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n290), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n287), .A2(G97), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n324), .A2(G1), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n286), .A2(new_n291), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n533), .B1(G97), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n512), .A2(new_n532), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n532), .A2(new_n538), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n497), .A2(new_n506), .A3(new_n280), .ZN(new_n541));
  AOI21_X1  g0341(.A(G169), .B1(new_n497), .B2(new_n506), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(KEYINPUT82), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT82), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n537), .B1(new_n531), .B2(new_n290), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n497), .A2(new_n506), .A3(new_n280), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n511), .B2(G169), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n545), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n539), .B1(new_n544), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(G116), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n289), .A2(new_n211), .B1(G20), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n493), .B1(new_n518), .B2(G33), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n552), .B1(new_n526), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT20), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n552), .B(KEYINPUT20), .C1(new_n526), .C2(new_n553), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n556), .A2(new_n557), .B1(new_n551), .B2(new_n287), .ZN(new_n558));
  AOI211_X1 g0358(.A(new_n534), .B(new_n290), .C1(new_n284), .C2(new_n285), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT84), .B1(new_n559), .B2(G116), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n286), .A2(new_n291), .A3(G116), .A4(new_n535), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT84), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n558), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n474), .B(G270), .C1(new_n498), .C2(new_n500), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n565), .A2(new_n504), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n325), .A2(new_n327), .A3(G264), .A4(G1698), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n325), .A2(new_n327), .A3(G257), .A4(new_n248), .ZN(new_n568));
  INV_X1    g0368(.A(G303), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n567), .B(new_n568), .C1(new_n569), .C2(new_n245), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n252), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n415), .B1(new_n566), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n564), .A2(new_n572), .A3(KEYINPUT21), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT85), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n564), .A2(new_n572), .A3(KEYINPUT85), .A4(KEYINPUT21), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n571), .A2(new_n504), .A3(new_n565), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n369), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(G190), .B2(new_n578), .ZN(new_n580));
  INV_X1    g0380(.A(new_n564), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n564), .A2(new_n572), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT21), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n571), .A2(G179), .A3(new_n504), .A4(new_n565), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n583), .A2(new_n584), .B1(new_n564), .B2(new_n586), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n577), .A2(new_n582), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT88), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n502), .A2(new_n503), .B1(new_n274), .B2(new_n275), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n325), .A2(new_n327), .A3(G250), .A4(new_n248), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n325), .A2(new_n327), .A3(G257), .A4(G1698), .ZN(new_n592));
  INV_X1    g0392(.A(G294), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n591), .B(new_n592), .C1(new_n324), .C2(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n590), .A2(G264), .B1(new_n594), .B2(new_n252), .ZN(new_n595));
  AOI21_X1  g0395(.A(G169), .B1(new_n595), .B2(new_n504), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n252), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n474), .B(G264), .C1(new_n498), .C2(new_n500), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n598), .A3(new_n504), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(G179), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n589), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n415), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n602), .B(KEYINPUT88), .C1(G179), .C2(new_n599), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT86), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT25), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n286), .B2(G107), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n284), .A2(new_n383), .A3(new_n285), .A4(new_n605), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n604), .A2(KEYINPUT25), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT87), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n536), .A2(new_n383), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n610), .B1(new_n607), .B2(new_n608), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT87), .B1(new_n617), .B2(new_n614), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(KEYINPUT23), .A2(G107), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n621));
  NOR2_X1   g0421(.A1(KEYINPUT23), .A2(G107), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  OAI221_X1 g0423(.A(new_n620), .B1(G20), .B2(new_n621), .C1(new_n210), .C2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n210), .A2(new_n245), .A3(G87), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT22), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT22), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n210), .A2(new_n245), .A3(new_n627), .A4(G87), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n624), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n291), .B1(new_n629), .B2(KEYINPUT24), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(KEYINPUT24), .B2(new_n629), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n601), .A2(new_n603), .B1(new_n619), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n599), .A2(new_n369), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(G190), .B2(new_n599), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n619), .A2(new_n634), .A3(new_n631), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n325), .A2(new_n327), .A3(G238), .A4(new_n248), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n325), .A2(new_n327), .A3(G244), .A4(G1698), .ZN(new_n637));
  NAND2_X1  g0437(.A1(G33), .A2(G116), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n252), .ZN(new_n640));
  OAI21_X1  g0440(.A(G250), .B1(new_n262), .B2(G1), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n262), .B2(new_n259), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n474), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n640), .A2(G190), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n369), .B1(new_n640), .B2(new_n643), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n430), .A2(new_n432), .A3(G33), .A4(G97), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT19), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(G87), .A2(G97), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n383), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n330), .A2(new_n648), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n651), .B1(new_n526), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n210), .A2(new_n245), .A3(G68), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n649), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n290), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n287), .A2(new_n376), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n559), .A2(G87), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n646), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n640), .A2(new_n280), .A3(new_n643), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT83), .ZN(new_n662));
  INV_X1    g0462(.A(new_n376), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n559), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n656), .A2(new_n657), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT83), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n640), .A2(new_n666), .A3(new_n280), .A4(new_n643), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n640), .A2(new_n643), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n415), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n662), .A2(new_n665), .A3(new_n667), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n660), .A2(new_n670), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n632), .A2(new_n635), .A3(new_n671), .ZN(new_n672));
  AND4_X1   g0472(.A1(new_n487), .A2(new_n550), .A3(new_n588), .A4(new_n672), .ZN(G372));
  INV_X1    g0473(.A(KEYINPUT90), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n338), .A2(new_n344), .B1(new_n348), .B2(new_n349), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n362), .A2(new_n365), .B1(new_n370), .B2(new_n371), .ZN(new_n676));
  OAI22_X1  g0476(.A1(new_n675), .A2(new_n366), .B1(new_n676), .B2(new_n394), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n453), .A2(KEYINPUT17), .A3(new_n481), .ZN(new_n678));
  AOI21_X1  g0478(.A(KEYINPUT17), .B1(new_n453), .B2(new_n481), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n454), .A2(new_n469), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n674), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n319), .A2(new_n320), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n682), .B1(new_n677), .B2(new_n680), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n684), .B1(new_n685), .B2(KEYINPUT90), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n683), .A2(new_n686), .B1(new_n306), .B2(new_n281), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n613), .B1(new_n612), .B2(new_n615), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n617), .A2(KEYINPUT87), .A3(new_n614), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n626), .A2(new_n628), .ZN(new_n690));
  INV_X1    g0490(.A(new_n624), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT24), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n290), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n629), .A2(KEYINPUT24), .ZN(new_n695));
  OAI22_X1  g0495(.A1(new_n688), .A2(new_n689), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n596), .A2(new_n600), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n577), .A2(new_n698), .A3(new_n587), .ZN(new_n699));
  INV_X1    g0499(.A(new_n635), .ZN(new_n700));
  AOI22_X1  g0500(.A1(new_n655), .A2(new_n290), .B1(new_n287), .B2(new_n376), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n701), .A2(new_n664), .B1(new_n415), .B2(new_n668), .ZN(new_n702));
  AOI22_X1  g0502(.A1(new_n661), .A2(new_n702), .B1(new_n646), .B2(new_n659), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n550), .A2(new_n699), .A3(new_n700), .A4(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n544), .A2(new_n549), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT26), .B1(new_n705), .B2(new_n671), .ZN(new_n706));
  OAI21_X1  g0506(.A(KEYINPUT89), .B1(new_n541), .B2(new_n542), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n497), .A2(new_n506), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n415), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT89), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(new_n710), .A3(new_n547), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT26), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n712), .A2(new_n713), .A3(new_n540), .A4(new_n703), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n702), .A2(new_n661), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n704), .A2(new_n706), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n487), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n687), .A2(new_n718), .ZN(G369));
  NAND3_X1  g0519(.A1(new_n210), .A2(new_n258), .A3(G13), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(KEYINPUT27), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(KEYINPUT27), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(G213), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G343), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n619), .B2(new_n631), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n726), .A2(new_n632), .A3(new_n635), .ZN(new_n727));
  INV_X1    g0527(.A(new_n725), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n727), .B1(new_n632), .B2(new_n728), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n577), .A2(new_n587), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(new_n728), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n728), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n727), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n581), .A2(new_n725), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n588), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n736), .B1(new_n730), .B2(new_n735), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G330), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n698), .A2(new_n728), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(new_n732), .B2(new_n727), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n740), .A2(new_n742), .ZN(G399));
  INV_X1    g0543(.A(new_n207), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n261), .A2(new_n263), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n650), .A2(new_n383), .A3(new_n551), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n747), .A2(G1), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n218), .B2(new_n747), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT28), .ZN(new_n752));
  INV_X1    g0552(.A(G330), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT93), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n597), .A2(new_n640), .A3(new_n598), .A4(new_n643), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n586), .A2(new_n756), .A3(new_n511), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT30), .ZN(new_n758));
  AND3_X1   g0558(.A1(new_n578), .A2(new_n280), .A3(new_n668), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n504), .A2(new_n595), .B1(new_n497), .B2(new_n506), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n757), .A2(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n708), .A2(new_n755), .A3(new_n585), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(KEYINPUT30), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n725), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n754), .B1(new_n764), .B2(KEYINPUT31), .ZN(new_n765));
  XNOR2_X1  g0565(.A(KEYINPUT91), .B(KEYINPUT31), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n725), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n391), .B1(new_n566), .B2(new_n571), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n768), .A2(new_n708), .A3(new_n599), .A4(new_n668), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(new_n762), .B2(KEYINPUT30), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT92), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n763), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n761), .A2(KEYINPUT92), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n767), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n757), .A2(new_n758), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n728), .B1(new_n770), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT31), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n776), .A2(KEYINPUT93), .A3(new_n777), .ZN(new_n778));
  AND3_X1   g0578(.A1(new_n765), .A2(new_n774), .A3(new_n778), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n672), .A2(new_n588), .A3(new_n550), .A4(new_n725), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n753), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n717), .A2(new_n725), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT29), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT89), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n710), .B1(new_n709), .B2(new_n547), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n703), .B(new_n540), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(KEYINPUT26), .ZN(new_n788));
  INV_X1    g0588(.A(new_n671), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n544), .A2(new_n789), .A3(new_n549), .A4(new_n713), .ZN(new_n790));
  AND3_X1   g0590(.A1(new_n788), .A2(new_n715), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n601), .A2(new_n603), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(new_n696), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n793), .A2(new_n577), .A3(new_n587), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n794), .A2(new_n550), .A3(new_n700), .A4(new_n703), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n728), .B1(new_n791), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(KEYINPUT29), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n781), .B1(new_n784), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n752), .B1(new_n798), .B2(G1), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT94), .ZN(G364));
  INV_X1    g0600(.A(new_n738), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n737), .A2(G330), .ZN(new_n802));
  INV_X1    g0602(.A(G13), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n526), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G45), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n805), .A2(new_n747), .A3(G1), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT95), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n801), .A2(new_n802), .A3(new_n811), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT96), .Z(new_n813));
  AOI21_X1  g0613(.A(new_n211), .B1(G20), .B2(new_n415), .ZN(new_n814));
  OR3_X1    g0614(.A1(new_n210), .A2(KEYINPUT98), .A3(G190), .ZN(new_n815));
  OAI21_X1  g0615(.A(KEYINPUT98), .B1(new_n210), .B2(G190), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n369), .A2(G179), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n819), .A2(KEYINPUT99), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(KEYINPUT99), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(G179), .A2(G200), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n815), .A2(new_n816), .A3(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n823), .A2(G283), .B1(G329), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT100), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n315), .A2(new_n369), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n391), .A2(new_n526), .A3(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(G326), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n315), .A2(G200), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n391), .A2(new_n526), .A3(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(G322), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n315), .A2(G179), .A3(G200), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n210), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(G294), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n817), .A2(G20), .A3(G190), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n245), .B1(new_n842), .B2(G303), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n832), .A2(new_n836), .A3(new_n840), .A4(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(G311), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n391), .A2(new_n315), .A3(new_n526), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(G200), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n846), .A2(new_n369), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  XOR2_X1   g0650(.A(KEYINPUT33), .B(G317), .Z(new_n851));
  OAI22_X1  g0651(.A1(new_n845), .A2(new_n848), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n828), .A2(new_n844), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n822), .A2(new_n383), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n826), .A2(G159), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT32), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n838), .A2(new_n518), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n435), .B(new_n857), .C1(G87), .C2(new_n842), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n858), .B1(new_n202), .B2(new_n830), .C1(new_n214), .C2(new_n834), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n215), .A2(new_n850), .B1(new_n848), .B2(new_n247), .ZN(new_n860));
  NOR4_X1   g0660(.A1(new_n854), .A2(new_n856), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n814), .B1(new_n853), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n245), .A2(new_n207), .ZN(new_n863));
  INV_X1    g0663(.A(G355), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n863), .A2(new_n864), .B1(G116), .B2(new_n207), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n218), .A2(new_n262), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n240), .B2(new_n262), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n744), .A2(new_n245), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n865), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(G13), .A2(G33), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n871), .A2(G20), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n872), .A2(new_n814), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n811), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT97), .ZN(new_n876));
  INV_X1    g0676(.A(new_n872), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n862), .B(new_n876), .C1(new_n737), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n813), .A2(new_n878), .ZN(G396));
  OAI211_X1 g0679(.A(new_n394), .B(new_n398), .C1(new_n395), .C2(new_n725), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT102), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n394), .B2(new_n725), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n395), .B1(new_n389), .B2(new_n392), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(KEYINPUT102), .A3(new_n728), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n880), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n782), .B(new_n886), .ZN(new_n887));
  OR2_X1    g0687(.A1(new_n887), .A2(new_n781), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(KEYINPUT103), .A3(new_n781), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n888), .A2(new_n810), .A3(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n887), .A2(new_n781), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n891), .A2(KEYINPUT103), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n885), .A2(new_n870), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n814), .A2(new_n870), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT101), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n811), .B1(G77), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(G283), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n551), .A2(new_n848), .B1(new_n850), .B2(new_n897), .ZN(new_n898));
  AOI211_X1 g0698(.A(new_n245), .B(new_n857), .C1(G107), .C2(new_n842), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n593), .B2(new_n834), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n898), .B(new_n900), .C1(G303), .C2(new_n831), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n823), .A2(G87), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n901), .B(new_n902), .C1(new_n845), .C2(new_n825), .ZN(new_n903));
  AOI22_X1  g0703(.A1(G137), .A2(new_n831), .B1(new_n835), .B2(G143), .ZN(new_n904));
  INV_X1    g0704(.A(G150), .ZN(new_n905));
  OAI221_X1 g0705(.A(new_n904), .B1(new_n850), .B2(new_n905), .C1(new_n425), .C2(new_n848), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT34), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n838), .A2(new_n214), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n245), .B1(new_n841), .B2(new_n202), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n909), .B(new_n910), .C1(new_n826), .C2(G132), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n907), .A2(new_n906), .B1(new_n822), .B2(new_n215), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n903), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n896), .B1(new_n914), .B2(new_n814), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n890), .A2(new_n892), .B1(new_n893), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(G384));
  NOR2_X1   g0717(.A1(new_n804), .A2(new_n258), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n367), .B(new_n728), .C1(new_n351), .C2(new_n676), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n362), .A2(new_n365), .A3(new_n728), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n373), .B(new_n920), .C1(new_n675), .C2(new_n366), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n885), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  AOI211_X1 g0722(.A(new_n777), .B(new_n725), .C1(new_n761), .C2(new_n763), .ZN(new_n923));
  INV_X1    g0723(.A(new_n766), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n757), .A2(new_n758), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n763), .A2(new_n925), .A3(new_n769), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n924), .B1(new_n926), .B2(new_n728), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n780), .A2(new_n928), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n922), .A2(new_n929), .A3(KEYINPUT40), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n465), .A2(new_n467), .A3(new_n411), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n465), .A2(new_n724), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n931), .A2(new_n482), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT37), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT37), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n931), .A2(new_n932), .A3(new_n935), .A4(new_n482), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(KEYINPUT104), .B1(new_n678), .B2(new_n679), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT104), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n484), .A2(new_n939), .A3(new_n485), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n682), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n937), .B1(new_n941), .B2(new_n932), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT38), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n462), .A2(new_n290), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n436), .A2(new_n440), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT16), .B1(new_n946), .B2(new_n458), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n464), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n724), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n486), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n947), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n421), .B1(new_n952), .B2(new_n442), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n482), .B(new_n949), .C1(new_n418), .C2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT37), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n936), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n951), .A2(new_n956), .A3(KEYINPUT38), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n944), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n930), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n922), .A2(new_n929), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n951), .A2(new_n956), .A3(KEYINPUT38), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT38), .B1(new_n951), .B2(new_n956), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n960), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n959), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n487), .A2(new_n929), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n966), .B(new_n967), .Z(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(G330), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT107), .Z(new_n970));
  NAND3_X1  g0770(.A1(new_n717), .A2(new_n725), .A3(new_n886), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n394), .A2(new_n728), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n964), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n919), .A2(new_n921), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n454), .A2(new_n469), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n978), .A2(new_n724), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT39), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n951), .A2(new_n956), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n943), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n981), .B1(new_n983), .B2(new_n957), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n962), .B1(new_n943), .B2(new_n942), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n984), .B1(new_n981), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n368), .A2(new_n728), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n977), .B(new_n980), .C1(new_n986), .C2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT105), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n678), .A2(new_n679), .A3(KEYINPUT104), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n939), .B1(new_n484), .B2(new_n485), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n978), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n932), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n993), .A2(new_n994), .B1(new_n936), .B2(new_n934), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n981), .B(new_n957), .C1(new_n995), .C2(KEYINPUT38), .ZN(new_n996));
  OAI21_X1  g0796(.A(KEYINPUT39), .B1(new_n962), .B2(new_n963), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n979), .B1(new_n998), .B2(new_n987), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT105), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n999), .A2(new_n1000), .A3(new_n977), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n990), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n784), .A2(new_n797), .A3(new_n487), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n687), .A2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1002), .B(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n918), .B1(new_n970), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n970), .B2(new_n1005), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n422), .A2(G77), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n218), .A2(new_n1008), .B1(G50), .B2(new_n215), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1009), .A2(G1), .A3(new_n803), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n525), .A2(KEYINPUT35), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n525), .A2(KEYINPUT35), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1011), .A2(G116), .A3(new_n212), .A4(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT36), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1007), .A2(new_n1010), .A3(new_n1014), .ZN(G367));
  NOR2_X1   g0815(.A1(new_n725), .A2(new_n659), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n703), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n715), .B2(new_n1016), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1018), .A2(KEYINPUT43), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n550), .B1(new_n546), .B2(new_n725), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n712), .A2(new_n540), .A3(new_n728), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  OR3_X1    g0824(.A1(new_n1024), .A2(KEYINPUT42), .A3(new_n733), .ZN(new_n1025));
  OAI21_X1  g0825(.A(KEYINPUT42), .B1(new_n1024), .B2(new_n733), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n1023), .A2(new_n632), .B1(new_n549), .B2(new_n544), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1025), .B(new_n1026), .C1(new_n728), .C2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1018), .A2(KEYINPUT43), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1020), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n740), .A2(new_n1024), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1028), .A2(new_n1020), .A3(new_n1029), .ZN(new_n1033));
  AND3_X1   g0833(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1032), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  XOR2_X1   g0836(.A(KEYINPUT108), .B(KEYINPUT41), .Z(new_n1037));
  XNOR2_X1  g0837(.A(new_n746), .B(new_n1037), .ZN(new_n1038));
  OR3_X1    g0838(.A1(new_n734), .A2(KEYINPUT109), .A3(new_n738), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n734), .A2(new_n738), .ZN(new_n1040));
  OAI21_X1  g0840(.A(KEYINPUT109), .B1(new_n734), .B2(new_n738), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n742), .A2(new_n1023), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT44), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n742), .A2(new_n1023), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT45), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n739), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1048), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1050), .A2(new_n740), .A3(new_n1045), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1043), .A2(new_n1049), .A3(new_n798), .A4(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1038), .B1(new_n1052), .B2(new_n798), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n805), .A2(G1), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1036), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n897), .A2(new_n848), .B1(new_n850), .B2(new_n593), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n842), .A2(G116), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT46), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n245), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n1058), .B2(new_n1057), .C1(new_n383), .C2(new_n838), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n569), .A2(new_n834), .B1(new_n830), .B2(new_n845), .ZN(new_n1061));
  INV_X1    g0861(.A(G317), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n518), .A2(new_n818), .B1(new_n825), .B2(new_n1062), .ZN(new_n1063));
  NOR4_X1   g0863(.A1(new_n1056), .A2(new_n1060), .A3(new_n1061), .A4(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n839), .A2(G68), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n905), .B2(new_n834), .ZN(new_n1066));
  INV_X1    g0866(.A(G143), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n1066), .A2(KEYINPUT110), .B1(new_n1067), .B2(new_n830), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(KEYINPUT110), .B2(new_n1066), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT111), .Z(new_n1070));
  INV_X1    g0870(.A(G137), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n247), .A2(new_n818), .B1(new_n825), .B2(new_n1071), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n245), .B1(new_n214), .B2(new_n841), .C1(new_n848), .C2(new_n202), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(G159), .C2(new_n849), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1064), .B1(new_n1070), .B2(new_n1074), .ZN(new_n1075));
  XOR2_X1   g0875(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n1076));
  OR2_X1    g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1077), .A2(new_n814), .A3(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n873), .B1(new_n207), .B2(new_n376), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n235), .B2(new_n868), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n810), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1079), .B(new_n1082), .C1(new_n877), .C2(new_n1018), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1055), .A2(new_n1083), .ZN(G387));
  NAND3_X1  g0884(.A1(new_n1043), .A2(KEYINPUT113), .A3(new_n1054), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT113), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1054), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1086), .B1(new_n1042), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n729), .A2(new_n872), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n863), .A2(new_n749), .B1(G107), .B2(new_n207), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n232), .A2(G45), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n299), .A2(G50), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT50), .ZN(new_n1093));
  AOI211_X1 g0893(.A(G45), .B(new_n748), .C1(G68), .C2(G77), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n744), .B(new_n245), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1090), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n811), .B1(new_n1096), .B2(new_n874), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n215), .A2(new_n848), .B1(new_n850), .B2(new_n299), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n838), .A2(new_n376), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n435), .B(new_n1099), .C1(G77), .C2(new_n842), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n202), .B2(new_n834), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1098), .B(new_n1101), .C1(G159), .C2(new_n831), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1102), .B1(new_n518), .B2(new_n822), .C1(new_n905), .C2(new_n825), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G317), .A2(new_n835), .B1(new_n831), .B2(G322), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1104), .B1(new_n850), .B2(new_n845), .C1(new_n569), .C2(new_n848), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT48), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n839), .A2(G283), .B1(G294), .B2(new_n842), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT49), .Z(new_n1111));
  INV_X1    g0911(.A(G326), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n435), .B1(new_n818), .B2(new_n551), .C1(new_n1112), .C2(new_n825), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1103), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1097), .B1(new_n1114), .B2(new_n814), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1085), .A2(new_n1088), .B1(new_n1089), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n747), .B1(new_n1043), .B2(new_n798), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT114), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n1117), .A2(new_n1118), .B1(new_n798), .B2(new_n1043), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1116), .B1(new_n1120), .B2(new_n1121), .ZN(G393));
  NAND2_X1  g0922(.A1(new_n1043), .A2(new_n798), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1125), .A2(new_n746), .A3(new_n1052), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT118), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1125), .A2(new_n1052), .A3(KEYINPUT118), .A4(new_n746), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1124), .A2(new_n1087), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1024), .A2(new_n872), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n873), .B1(new_n518), .B2(new_n207), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n243), .B2(new_n868), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n245), .B1(new_n247), .B2(new_n838), .C1(new_n850), .C2(new_n202), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(new_n300), .B2(new_n847), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n905), .A2(new_n830), .B1(new_n834), .B2(new_n425), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1136), .B(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n902), .A2(new_n1135), .A3(new_n1138), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n825), .A2(new_n1067), .B1(new_n215), .B2(new_n841), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT116), .Z(new_n1141));
  OAI221_X1 g0941(.A(new_n435), .B1(new_n897), .B2(new_n841), .C1(new_n838), .C2(new_n551), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n850), .A2(new_n569), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n1142), .B(new_n1143), .C1(G294), .C2(new_n847), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n845), .A2(new_n834), .B1(new_n830), .B2(new_n1062), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT52), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n826), .A2(G322), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1144), .B(new_n1147), .C1(new_n1146), .C2(new_n1145), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n1139), .A2(new_n1141), .B1(new_n1148), .B2(new_n854), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1149), .A2(KEYINPUT117), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1150), .A2(new_n814), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1149), .A2(KEYINPUT117), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n810), .B(new_n1133), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1130), .B1(new_n1131), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1128), .A2(new_n1129), .A3(new_n1154), .ZN(G390));
  OAI21_X1  g0955(.A(new_n811), .B1(new_n300), .B2(new_n895), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT119), .Z(new_n1157));
  NAND2_X1  g0957(.A1(new_n842), .A2(G150), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT53), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n435), .B(new_n1159), .C1(G159), .C2(new_n839), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G128), .A2(new_n831), .B1(new_n835), .B2(G132), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(G125), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1162), .B1(new_n202), .B2(new_n818), .C1(new_n1163), .C2(new_n825), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT54), .B(G143), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(G137), .A2(new_n849), .B1(new_n847), .B2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT120), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n822), .A2(new_n215), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n245), .B1(new_n842), .B2(G87), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT121), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G97), .B2(new_n847), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n849), .A2(G107), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n826), .A2(G294), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n830), .A2(new_n897), .B1(new_n247), .B2(new_n838), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G116), .B2(new_n835), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .A4(new_n1176), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n1164), .A2(new_n1168), .B1(new_n1169), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1157), .B1(new_n1178), .B2(new_n814), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n998), .B2(new_n871), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n987), .B1(new_n944), .B2(new_n957), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n972), .B1(new_n796), .B2(new_n886), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n976), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n987), .B1(new_n974), .B2(new_n976), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1184), .B1(new_n1185), .B2(new_n998), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n929), .A2(G330), .A3(new_n886), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1187), .A2(new_n1183), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n781), .A2(new_n922), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1184), .B(new_n1190), .C1(new_n1185), .C2(new_n998), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1180), .B1(new_n1192), .B2(new_n1087), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n487), .A2(G330), .A3(new_n929), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n687), .A2(new_n1003), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n976), .B1(new_n781), .B2(new_n886), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n974), .B1(new_n1196), .B2(new_n1188), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1187), .A2(new_n1183), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1190), .A2(new_n1182), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1195), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n747), .B1(new_n1201), .B2(new_n1192), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1200), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1193), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(G378));
  INV_X1    g1005(.A(new_n1191), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1188), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1183), .B1(new_n971), .B2(new_n973), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n997), .B(new_n996), .C1(new_n1208), .C2(new_n987), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1207), .B1(new_n1209), .B2(new_n1184), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1206), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1195), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n959), .A2(new_n965), .A3(G330), .ZN(new_n1214));
  XOR2_X1   g1014(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1215));
  NOR2_X1   g1015(.A1(new_n305), .A2(new_n723), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n321), .A2(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n321), .A2(new_n1216), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1215), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n321), .A2(new_n1216), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n321), .A2(new_n1216), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1215), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1219), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1214), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1219), .A2(new_n1223), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1226), .A2(new_n959), .A3(new_n965), .A4(G330), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n998), .A2(new_n987), .ZN(new_n1229));
  AND4_X1   g1029(.A1(new_n1000), .A2(new_n1229), .A3(new_n977), .A4(new_n980), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1000), .B1(new_n999), .B2(new_n977), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1228), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n990), .A2(new_n1001), .A3(new_n1225), .A4(new_n1227), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(KEYINPUT57), .B1(new_n1213), .B2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1195), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1203), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT57), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1237), .A2(new_n1238), .A3(new_n1233), .A4(new_n1232), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n747), .B1(new_n1235), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1224), .A2(new_n870), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n811), .B1(G50), .B2(new_n895), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n819), .A2(G58), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n245), .B(new_n745), .C1(new_n842), .C2(G77), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1243), .B(new_n1244), .C1(new_n897), .C2(new_n825), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT122), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1065), .B1(new_n383), .B2(new_n834), .C1(new_n551), .C2(new_n830), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n518), .A2(new_n850), .B1(new_n848), .B2(new_n376), .ZN(new_n1248));
  OR3_X1    g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT58), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n745), .A2(new_n245), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(G33), .A2(G41), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1253), .A2(G50), .A3(new_n1254), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n839), .A2(G150), .B1(new_n842), .B2(new_n1166), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n1163), .B2(new_n830), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n849), .A2(G132), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n848), .B2(new_n1071), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n1257), .B(new_n1259), .C1(G128), .C2(new_n835), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT59), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  XOR2_X1   g1062(.A(KEYINPUT123), .B(G124), .Z(new_n1263));
  OAI221_X1 g1063(.A(new_n1254), .B1(new_n818), .B2(new_n425), .C1(new_n825), .C2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1255), .B1(new_n1262), .B2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1251), .A2(new_n1252), .A3(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1242), .B1(new_n1267), .B2(new_n814), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1241), .A2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n1234), .B2(new_n1087), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1240), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(G375));
  NOR2_X1   g1072(.A1(new_n1200), .A2(new_n1038), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n1236), .B2(new_n1212), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1183), .A2(new_n870), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n811), .B1(G68), .B2(new_n895), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n834), .A2(new_n1071), .ZN(new_n1277));
  OAI221_X1 g1077(.A(new_n245), .B1(new_n425), .B2(new_n841), .C1(new_n838), .C2(new_n202), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1277), .B(new_n1278), .C1(G132), .C2(new_n831), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(G150), .A2(new_n847), .B1(new_n849), .B2(new_n1166), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n826), .A2(G128), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1279), .A2(new_n1243), .A3(new_n1280), .A4(new_n1281), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n822), .A2(new_n247), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n435), .B1(new_n841), .B2(new_n518), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n1284), .B(new_n1099), .C1(G283), .C2(new_n835), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(G107), .A2(new_n847), .B1(new_n849), .B2(G116), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n826), .A2(G303), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n831), .A2(G294), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .A4(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1282), .B1(new_n1283), .B2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1276), .B1(new_n1290), .B2(new_n814), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(new_n1212), .A2(new_n1054), .B1(new_n1275), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1274), .A2(new_n1292), .ZN(G381));
  NAND2_X1  g1093(.A1(new_n1271), .A2(new_n1204), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1154), .A2(new_n1129), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1295), .A2(new_n1055), .A3(new_n1083), .A4(new_n1128), .ZN(new_n1296));
  INV_X1    g1096(.A(G396), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1297), .B(new_n1116), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1298));
  OR3_X1    g1098(.A1(new_n1298), .A2(G384), .A3(G381), .ZN(new_n1299));
  OR3_X1    g1099(.A1(new_n1294), .A2(new_n1296), .A3(new_n1299), .ZN(G407));
  OAI211_X1 g1100(.A(G407), .B(G213), .C1(G343), .C2(new_n1294), .ZN(G409));
  NAND2_X1  g1101(.A1(G387), .A2(G390), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1296), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(G393), .A2(G396), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n1298), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1298), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(new_n1296), .A3(new_n1302), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  OR3_X1    g1108(.A1(new_n1212), .A2(new_n1236), .A3(KEYINPUT60), .ZN(new_n1309));
  OAI21_X1  g1109(.A(KEYINPUT60), .B1(new_n1212), .B2(new_n1236), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1200), .A2(new_n747), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1292), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n916), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1292), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1316), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(G384), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1315), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(G213), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1321), .A2(G343), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  NOR3_X1   g1123(.A1(new_n1240), .A2(new_n1204), .A3(new_n1270), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1270), .ZN(new_n1325));
  OR3_X1    g1125(.A1(new_n1213), .A2(new_n1234), .A3(new_n1038), .ZN(new_n1326));
  AOI21_X1  g1126(.A(G378), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1320), .B(new_n1323), .C1(new_n1324), .C2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT125), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1328), .A2(new_n1329), .A3(KEYINPUT62), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1323), .B1(new_n1324), .B2(new_n1327), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1317), .A2(G384), .ZN(new_n1332));
  AOI211_X1 g1132(.A(new_n1316), .B(new_n916), .C1(new_n1311), .C2(new_n1312), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1322), .A2(G2897), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  NOR3_X1   g1135(.A1(new_n1332), .A2(new_n1333), .A3(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1334), .B1(new_n1315), .B2(new_n1318), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(KEYINPUT61), .B1(new_n1331), .B2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1330), .A2(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(KEYINPUT62), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1308), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT124), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1235), .A2(new_n1239), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1344), .A2(new_n746), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1345), .A2(G378), .A3(new_n1325), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1327), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1322), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1319), .A2(new_n1335), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1315), .A2(new_n1318), .A3(new_n1334), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1343), .B1(new_n1348), .B2(new_n1351), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1331), .A2(new_n1338), .A3(KEYINPUT124), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT63), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1348), .A2(new_n1355), .A3(new_n1320), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1328), .A2(KEYINPUT63), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1356), .A2(new_n1357), .ZN(new_n1358));
  NOR2_X1   g1158(.A1(new_n1308), .A2(KEYINPUT61), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1354), .A2(new_n1358), .A3(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1342), .A2(new_n1360), .ZN(G405));
  OAI21_X1  g1161(.A(G378), .B1(new_n1240), .B2(new_n1270), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1319), .B1(new_n1294), .B2(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1363), .ZN(new_n1364));
  AND3_X1   g1164(.A1(new_n1306), .A2(new_n1296), .A3(new_n1302), .ZN(new_n1365));
  AOI21_X1  g1165(.A(new_n1306), .B1(new_n1296), .B2(new_n1302), .ZN(new_n1366));
  NOR2_X1   g1166(.A1(new_n1365), .A2(new_n1366), .ZN(new_n1367));
  INV_X1    g1167(.A(KEYINPUT126), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n1294), .A2(new_n1319), .A3(new_n1362), .ZN(new_n1369));
  NAND4_X1  g1169(.A1(new_n1364), .A2(new_n1367), .A3(new_n1368), .A4(new_n1369), .ZN(new_n1370));
  AND3_X1   g1170(.A1(new_n1294), .A2(new_n1319), .A3(new_n1362), .ZN(new_n1371));
  OAI21_X1  g1171(.A(new_n1308), .B1(new_n1371), .B2(new_n1363), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1370), .A2(new_n1372), .ZN(new_n1373));
  NOR2_X1   g1173(.A1(new_n1371), .A2(new_n1363), .ZN(new_n1374));
  AOI21_X1  g1174(.A(new_n1368), .B1(new_n1374), .B2(new_n1367), .ZN(new_n1375));
  NOR2_X1   g1175(.A1(new_n1373), .A2(new_n1375), .ZN(G402));
endmodule


