

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(G651), .A2(n624), .ZN(n646) );
  XNOR2_X2 U556 ( .A(KEYINPUT15), .B(n571), .ZN(n924) );
  NOR2_X1 U557 ( .A1(n779), .A2(n778), .ZN(n788) );
  OR2_X1 U558 ( .A1(n723), .A2(n728), .ZN(n724) );
  XNOR2_X1 U559 ( .A(n771), .B(n770), .ZN(n779) );
  XNOR2_X1 U560 ( .A(KEYINPUT27), .B(KEYINPUT98), .ZN(n732) );
  XNOR2_X1 U561 ( .A(n733), .B(n732), .ZN(n736) );
  AND2_X1 U562 ( .A1(n713), .A2(n712), .ZN(n734) );
  INV_X1 U563 ( .A(KEYINPUT31), .ZN(n757) );
  INV_X1 U564 ( .A(KEYINPUT32), .ZN(n770) );
  NAND2_X1 U565 ( .A1(n712), .A2(n713), .ZN(n761) );
  INV_X1 U566 ( .A(KEYINPUT17), .ZN(n522) );
  NOR2_X1 U567 ( .A1(G2104), .A2(n529), .ZN(n890) );
  NOR2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  XNOR2_X1 U569 ( .A(n523), .B(n522), .ZN(n543) );
  NAND2_X1 U570 ( .A1(n543), .A2(G137), .ZN(n525) );
  AND2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n891) );
  NAND2_X1 U572 ( .A1(G113), .A2(n891), .ZN(n524) );
  NAND2_X1 U573 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U574 ( .A(n526), .B(KEYINPUT65), .ZN(n528) );
  INV_X1 U575 ( .A(G2105), .ZN(n529) );
  NAND2_X1 U576 ( .A1(G125), .A2(n890), .ZN(n527) );
  NAND2_X1 U577 ( .A1(n528), .A2(n527), .ZN(n532) );
  AND2_X1 U578 ( .A1(n529), .A2(G2104), .ZN(n886) );
  NAND2_X1 U579 ( .A1(G101), .A2(n886), .ZN(n530) );
  XNOR2_X1 U580 ( .A(KEYINPUT23), .B(n530), .ZN(n531) );
  NOR2_X1 U581 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U582 ( .A(n533), .B(KEYINPUT64), .ZN(n698) );
  BUF_X1 U583 ( .A(n698), .Z(G160) );
  XOR2_X1 U584 ( .A(G543), .B(KEYINPUT0), .Z(n624) );
  NAND2_X1 U585 ( .A1(G52), .A2(n646), .ZN(n536) );
  INV_X1 U586 ( .A(G651), .ZN(n537) );
  NOR2_X1 U587 ( .A1(G543), .A2(n537), .ZN(n534) );
  XOR2_X2 U588 ( .A(KEYINPUT1), .B(n534), .Z(n644) );
  NAND2_X1 U589 ( .A1(G64), .A2(n644), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n542) );
  NOR2_X1 U591 ( .A1(G651), .A2(G543), .ZN(n647) );
  NAND2_X1 U592 ( .A1(G90), .A2(n647), .ZN(n539) );
  NOR2_X1 U593 ( .A1(n624), .A2(n537), .ZN(n650) );
  NAND2_X1 U594 ( .A1(G77), .A2(n650), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U596 ( .A(KEYINPUT9), .B(n540), .Z(n541) );
  NOR2_X1 U597 ( .A1(n542), .A2(n541), .ZN(G171) );
  AND2_X1 U598 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U599 ( .A(G57), .ZN(G237) );
  INV_X1 U600 ( .A(G82), .ZN(G220) );
  BUF_X1 U601 ( .A(n543), .Z(n885) );
  NAND2_X1 U602 ( .A1(G138), .A2(n885), .ZN(n545) );
  NAND2_X1 U603 ( .A1(G102), .A2(n886), .ZN(n544) );
  NAND2_X1 U604 ( .A1(n545), .A2(n544), .ZN(n549) );
  NAND2_X1 U605 ( .A1(G126), .A2(n890), .ZN(n547) );
  NAND2_X1 U606 ( .A1(G114), .A2(n891), .ZN(n546) );
  NAND2_X1 U607 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U608 ( .A1(n549), .A2(n548), .ZN(G164) );
  NAND2_X1 U609 ( .A1(G7), .A2(G661), .ZN(n550) );
  XNOR2_X1 U610 ( .A(n550), .B(KEYINPUT10), .ZN(n551) );
  XNOR2_X1 U611 ( .A(KEYINPUT68), .B(n551), .ZN(G223) );
  INV_X1 U612 ( .A(G223), .ZN(n828) );
  NAND2_X1 U613 ( .A1(n828), .A2(G567), .ZN(n552) );
  XOR2_X1 U614 ( .A(KEYINPUT11), .B(n552), .Z(G234) );
  XNOR2_X1 U615 ( .A(KEYINPUT13), .B(KEYINPUT69), .ZN(n557) );
  NAND2_X1 U616 ( .A1(n647), .A2(G81), .ZN(n553) );
  XNOR2_X1 U617 ( .A(n553), .B(KEYINPUT12), .ZN(n555) );
  NAND2_X1 U618 ( .A1(G68), .A2(n650), .ZN(n554) );
  NAND2_X1 U619 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U620 ( .A(n557), .B(n556), .ZN(n560) );
  NAND2_X1 U621 ( .A1(n644), .A2(G56), .ZN(n558) );
  XOR2_X1 U622 ( .A(KEYINPUT14), .B(n558), .Z(n559) );
  NOR2_X1 U623 ( .A1(n560), .A2(n559), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n646), .A2(G43), .ZN(n561) );
  NAND2_X1 U625 ( .A1(n562), .A2(n561), .ZN(n929) );
  INV_X1 U626 ( .A(G860), .ZN(n598) );
  OR2_X1 U627 ( .A1(n929), .A2(n598), .ZN(G153) );
  INV_X1 U628 ( .A(G171), .ZN(G301) );
  INV_X1 U629 ( .A(G868), .ZN(n601) );
  NOR2_X1 U630 ( .A1(G301), .A2(n601), .ZN(n573) );
  NAND2_X1 U631 ( .A1(G92), .A2(n647), .ZN(n564) );
  NAND2_X1 U632 ( .A1(G79), .A2(n650), .ZN(n563) );
  NAND2_X1 U633 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U634 ( .A1(G54), .A2(n646), .ZN(n566) );
  NAND2_X1 U635 ( .A1(G66), .A2(n644), .ZN(n565) );
  NAND2_X1 U636 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U637 ( .A1(n568), .A2(n567), .ZN(n570) );
  XNOR2_X1 U638 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n569) );
  XNOR2_X1 U639 ( .A(n570), .B(n569), .ZN(n571) );
  INV_X1 U640 ( .A(n924), .ZN(n902) );
  NOR2_X1 U641 ( .A1(n902), .A2(G868), .ZN(n572) );
  NOR2_X1 U642 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U643 ( .A(KEYINPUT72), .B(n574), .ZN(G284) );
  XOR2_X1 U644 ( .A(KEYINPUT5), .B(KEYINPUT73), .Z(n575) );
  XNOR2_X1 U645 ( .A(KEYINPUT74), .B(n575), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n647), .A2(G89), .ZN(n576) );
  XNOR2_X1 U647 ( .A(n576), .B(KEYINPUT4), .ZN(n578) );
  NAND2_X1 U648 ( .A1(G76), .A2(n650), .ZN(n577) );
  NAND2_X1 U649 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U650 ( .A(n580), .B(n579), .ZN(n587) );
  XNOR2_X1 U651 ( .A(KEYINPUT76), .B(KEYINPUT6), .ZN(n585) );
  NAND2_X1 U652 ( .A1(G51), .A2(n646), .ZN(n582) );
  NAND2_X1 U653 ( .A1(G63), .A2(n644), .ZN(n581) );
  NAND2_X1 U654 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U655 ( .A(n583), .B(KEYINPUT75), .ZN(n584) );
  XNOR2_X1 U656 ( .A(n585), .B(n584), .ZN(n586) );
  NAND2_X1 U657 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U658 ( .A(n588), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U659 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U660 ( .A1(G53), .A2(n646), .ZN(n590) );
  NAND2_X1 U661 ( .A1(G65), .A2(n644), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U663 ( .A1(G91), .A2(n647), .ZN(n592) );
  NAND2_X1 U664 ( .A1(G78), .A2(n650), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n932) );
  INV_X1 U667 ( .A(n932), .ZN(G299) );
  NOR2_X1 U668 ( .A1(G286), .A2(n601), .ZN(n595) );
  XOR2_X1 U669 ( .A(KEYINPUT77), .B(n595), .Z(n597) );
  NOR2_X1 U670 ( .A1(G868), .A2(G299), .ZN(n596) );
  NOR2_X1 U671 ( .A1(n597), .A2(n596), .ZN(G297) );
  NAND2_X1 U672 ( .A1(n598), .A2(G559), .ZN(n599) );
  NAND2_X1 U673 ( .A1(n599), .A2(n924), .ZN(n600) );
  XNOR2_X1 U674 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U675 ( .A1(n902), .A2(n601), .ZN(n602) );
  XOR2_X1 U676 ( .A(KEYINPUT78), .B(n602), .Z(n603) );
  NOR2_X1 U677 ( .A1(G559), .A2(n603), .ZN(n605) );
  NOR2_X1 U678 ( .A1(G868), .A2(n929), .ZN(n604) );
  NOR2_X1 U679 ( .A1(n605), .A2(n604), .ZN(G282) );
  NAND2_X1 U680 ( .A1(G123), .A2(n890), .ZN(n606) );
  XNOR2_X1 U681 ( .A(n606), .B(KEYINPUT18), .ZN(n609) );
  NAND2_X1 U682 ( .A1(G111), .A2(n891), .ZN(n607) );
  XOR2_X1 U683 ( .A(KEYINPUT79), .B(n607), .Z(n608) );
  NAND2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U685 ( .A1(G135), .A2(n885), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G99), .A2(n886), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U688 ( .A1(n613), .A2(n612), .ZN(n980) );
  XOR2_X1 U689 ( .A(G2096), .B(n980), .Z(n614) );
  NOR2_X1 U690 ( .A1(G2100), .A2(n614), .ZN(n615) );
  XOR2_X1 U691 ( .A(KEYINPUT80), .B(n615), .Z(G156) );
  NAND2_X1 U692 ( .A1(G85), .A2(n647), .ZN(n617) );
  NAND2_X1 U693 ( .A1(G72), .A2(n650), .ZN(n616) );
  NAND2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U695 ( .A1(G47), .A2(n646), .ZN(n618) );
  XOR2_X1 U696 ( .A(KEYINPUT66), .B(n618), .Z(n619) );
  NOR2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n644), .A2(G60), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n622), .A2(n621), .ZN(G290) );
  NAND2_X1 U700 ( .A1(G49), .A2(n646), .ZN(n623) );
  XNOR2_X1 U701 ( .A(n623), .B(KEYINPUT84), .ZN(n629) );
  NAND2_X1 U702 ( .A1(G87), .A2(n624), .ZN(n626) );
  NAND2_X1 U703 ( .A1(G74), .A2(G651), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U705 ( .A1(n644), .A2(n627), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(G288) );
  NAND2_X1 U707 ( .A1(G86), .A2(n647), .ZN(n631) );
  NAND2_X1 U708 ( .A1(G61), .A2(n644), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n650), .A2(G73), .ZN(n632) );
  XOR2_X1 U711 ( .A(KEYINPUT2), .B(n632), .Z(n633) );
  NOR2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n646), .A2(G48), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n636), .A2(n635), .ZN(G305) );
  NAND2_X1 U715 ( .A1(G50), .A2(n646), .ZN(n638) );
  NAND2_X1 U716 ( .A1(G62), .A2(n644), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U718 ( .A(KEYINPUT85), .B(n639), .ZN(n643) );
  NAND2_X1 U719 ( .A1(G88), .A2(n647), .ZN(n641) );
  NAND2_X1 U720 ( .A1(G75), .A2(n650), .ZN(n640) );
  AND2_X1 U721 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U722 ( .A1(n643), .A2(n642), .ZN(G303) );
  INV_X1 U723 ( .A(G303), .ZN(G166) );
  NAND2_X1 U724 ( .A1(G67), .A2(n644), .ZN(n645) );
  XNOR2_X1 U725 ( .A(n645), .B(KEYINPUT82), .ZN(n655) );
  NAND2_X1 U726 ( .A1(G55), .A2(n646), .ZN(n649) );
  NAND2_X1 U727 ( .A1(G93), .A2(n647), .ZN(n648) );
  NAND2_X1 U728 ( .A1(n649), .A2(n648), .ZN(n653) );
  NAND2_X1 U729 ( .A1(G80), .A2(n650), .ZN(n651) );
  XNOR2_X1 U730 ( .A(KEYINPUT81), .B(n651), .ZN(n652) );
  NOR2_X1 U731 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U732 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U733 ( .A(KEYINPUT83), .B(n656), .ZN(n835) );
  NOR2_X1 U734 ( .A1(G868), .A2(n835), .ZN(n657) );
  XNOR2_X1 U735 ( .A(n657), .B(KEYINPUT87), .ZN(n667) );
  XNOR2_X1 U736 ( .A(n835), .B(G290), .ZN(n658) );
  XNOR2_X1 U737 ( .A(n658), .B(G288), .ZN(n662) );
  XNOR2_X1 U738 ( .A(G305), .B(KEYINPUT19), .ZN(n660) );
  XNOR2_X1 U739 ( .A(n932), .B(G166), .ZN(n659) );
  XNOR2_X1 U740 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U741 ( .A(n662), .B(n661), .ZN(n903) );
  XNOR2_X1 U742 ( .A(KEYINPUT86), .B(n903), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n924), .A2(G559), .ZN(n663) );
  XNOR2_X1 U744 ( .A(n663), .B(n929), .ZN(n834) );
  XNOR2_X1 U745 ( .A(n664), .B(n834), .ZN(n665) );
  NAND2_X1 U746 ( .A1(G868), .A2(n665), .ZN(n666) );
  NAND2_X1 U747 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U748 ( .A1(G2084), .A2(G2078), .ZN(n668) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n670), .ZN(n671) );
  NAND2_X1 U752 ( .A1(n671), .A2(G2072), .ZN(n672) );
  XNOR2_X1 U753 ( .A(KEYINPUT88), .B(n672), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U755 ( .A(KEYINPUT67), .B(G132), .ZN(G219) );
  NOR2_X1 U756 ( .A1(G220), .A2(G219), .ZN(n673) );
  XOR2_X1 U757 ( .A(KEYINPUT22), .B(n673), .Z(n674) );
  NOR2_X1 U758 ( .A1(G218), .A2(n674), .ZN(n675) );
  NAND2_X1 U759 ( .A1(G96), .A2(n675), .ZN(n832) );
  NAND2_X1 U760 ( .A1(n832), .A2(G2106), .ZN(n679) );
  NAND2_X1 U761 ( .A1(G69), .A2(G120), .ZN(n676) );
  NOR2_X1 U762 ( .A1(G237), .A2(n676), .ZN(n677) );
  NAND2_X1 U763 ( .A1(G108), .A2(n677), .ZN(n833) );
  NAND2_X1 U764 ( .A1(n833), .A2(G567), .ZN(n678) );
  NAND2_X1 U765 ( .A1(n679), .A2(n678), .ZN(n837) );
  NAND2_X1 U766 ( .A1(G661), .A2(G483), .ZN(n680) );
  XOR2_X1 U767 ( .A(KEYINPUT89), .B(n680), .Z(n681) );
  NOR2_X1 U768 ( .A1(n837), .A2(n681), .ZN(n831) );
  NAND2_X1 U769 ( .A1(n831), .A2(G36), .ZN(G176) );
  NAND2_X1 U770 ( .A1(G105), .A2(n886), .ZN(n682) );
  XNOR2_X1 U771 ( .A(n682), .B(KEYINPUT38), .ZN(n683) );
  XNOR2_X1 U772 ( .A(n683), .B(KEYINPUT92), .ZN(n685) );
  NAND2_X1 U773 ( .A1(G117), .A2(n891), .ZN(n684) );
  NAND2_X1 U774 ( .A1(n685), .A2(n684), .ZN(n688) );
  NAND2_X1 U775 ( .A1(G141), .A2(n885), .ZN(n686) );
  XNOR2_X1 U776 ( .A(KEYINPUT93), .B(n686), .ZN(n687) );
  NOR2_X1 U777 ( .A1(n688), .A2(n687), .ZN(n691) );
  NAND2_X1 U778 ( .A1(G129), .A2(n890), .ZN(n689) );
  XOR2_X1 U779 ( .A(KEYINPUT91), .B(n689), .Z(n690) );
  NAND2_X1 U780 ( .A1(n691), .A2(n690), .ZN(n874) );
  AND2_X1 U781 ( .A1(n874), .A2(G1996), .ZN(n983) );
  NAND2_X1 U782 ( .A1(G131), .A2(n885), .ZN(n693) );
  NAND2_X1 U783 ( .A1(G95), .A2(n886), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n693), .A2(n692), .ZN(n697) );
  NAND2_X1 U785 ( .A1(G119), .A2(n890), .ZN(n695) );
  NAND2_X1 U786 ( .A1(G107), .A2(n891), .ZN(n694) );
  NAND2_X1 U787 ( .A1(n695), .A2(n694), .ZN(n696) );
  OR2_X1 U788 ( .A1(n697), .A2(n696), .ZN(n878) );
  AND2_X1 U789 ( .A1(n878), .A2(G1991), .ZN(n981) );
  OR2_X1 U790 ( .A1(n983), .A2(n981), .ZN(n699) );
  NOR2_X1 U791 ( .A1(G164), .A2(G1384), .ZN(n713) );
  NAND2_X1 U792 ( .A1(n698), .A2(G40), .ZN(n711) );
  NOR2_X1 U793 ( .A1(n713), .A2(n711), .ZN(n823) );
  NAND2_X1 U794 ( .A1(n699), .A2(n823), .ZN(n813) );
  XNOR2_X1 U795 ( .A(KEYINPUT37), .B(G2067), .ZN(n821) );
  NAND2_X1 U796 ( .A1(G140), .A2(n885), .ZN(n701) );
  NAND2_X1 U797 ( .A1(G104), .A2(n886), .ZN(n700) );
  NAND2_X1 U798 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U799 ( .A(KEYINPUT34), .B(n702), .ZN(n708) );
  NAND2_X1 U800 ( .A1(G128), .A2(n890), .ZN(n704) );
  NAND2_X1 U801 ( .A1(G116), .A2(n891), .ZN(n703) );
  NAND2_X1 U802 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U803 ( .A(KEYINPUT35), .B(n705), .Z(n706) );
  XNOR2_X1 U804 ( .A(KEYINPUT90), .B(n706), .ZN(n707) );
  NOR2_X1 U805 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U806 ( .A(KEYINPUT36), .B(n709), .ZN(n897) );
  NOR2_X1 U807 ( .A1(n821), .A2(n897), .ZN(n987) );
  NAND2_X1 U808 ( .A1(n823), .A2(n987), .ZN(n819) );
  NAND2_X1 U809 ( .A1(n813), .A2(n819), .ZN(n710) );
  XNOR2_X1 U810 ( .A(n710), .B(KEYINPUT94), .ZN(n809) );
  INV_X1 U811 ( .A(n711), .ZN(n712) );
  XNOR2_X1 U812 ( .A(KEYINPUT97), .B(G1961), .ZN(n1006) );
  NAND2_X1 U813 ( .A1(n761), .A2(n1006), .ZN(n715) );
  XNOR2_X1 U814 ( .A(G2078), .B(KEYINPUT25), .ZN(n957) );
  NAND2_X1 U815 ( .A1(n734), .A2(n957), .ZN(n714) );
  NAND2_X1 U816 ( .A1(n715), .A2(n714), .ZN(n754) );
  NAND2_X1 U817 ( .A1(n754), .A2(G171), .ZN(n747) );
  NAND2_X1 U818 ( .A1(G1348), .A2(n761), .ZN(n717) );
  NAND2_X1 U819 ( .A1(G2067), .A2(n734), .ZN(n716) );
  NAND2_X1 U820 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U821 ( .A(KEYINPUT99), .B(n718), .Z(n725) );
  INV_X1 U822 ( .A(n929), .ZN(n720) );
  NAND2_X1 U823 ( .A1(n761), .A2(G1341), .ZN(n719) );
  NAND2_X1 U824 ( .A1(n720), .A2(n719), .ZN(n727) );
  INV_X1 U825 ( .A(n727), .ZN(n721) );
  NAND2_X1 U826 ( .A1(n924), .A2(n721), .ZN(n723) );
  AND2_X1 U827 ( .A1(n734), .A2(G1996), .ZN(n722) );
  XNOR2_X1 U828 ( .A(n722), .B(KEYINPUT26), .ZN(n728) );
  NAND2_X1 U829 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U830 ( .A(n726), .B(KEYINPUT100), .ZN(n731) );
  NOR2_X1 U831 ( .A1(n728), .A2(n727), .ZN(n729) );
  OR2_X1 U832 ( .A1(n729), .A2(n924), .ZN(n730) );
  NAND2_X1 U833 ( .A1(n731), .A2(n730), .ZN(n738) );
  NAND2_X1 U834 ( .A1(G2072), .A2(n734), .ZN(n733) );
  INV_X1 U835 ( .A(G1956), .ZN(n1007) );
  NOR2_X1 U836 ( .A1(n734), .A2(n1007), .ZN(n735) );
  NOR2_X1 U837 ( .A1(n736), .A2(n735), .ZN(n739) );
  NAND2_X1 U838 ( .A1(n932), .A2(n739), .ZN(n737) );
  NAND2_X1 U839 ( .A1(n738), .A2(n737), .ZN(n743) );
  NOR2_X1 U840 ( .A1(n739), .A2(n932), .ZN(n741) );
  INV_X1 U841 ( .A(KEYINPUT28), .ZN(n740) );
  XNOR2_X1 U842 ( .A(n741), .B(n740), .ZN(n742) );
  NAND2_X1 U843 ( .A1(n743), .A2(n742), .ZN(n745) );
  XNOR2_X1 U844 ( .A(KEYINPUT29), .B(KEYINPUT101), .ZN(n744) );
  XNOR2_X1 U845 ( .A(n745), .B(n744), .ZN(n746) );
  NAND2_X1 U846 ( .A1(n747), .A2(n746), .ZN(n760) );
  NAND2_X1 U847 ( .A1(n761), .A2(G8), .ZN(n748) );
  XNOR2_X1 U848 ( .A(n748), .B(KEYINPUT95), .ZN(n791) );
  INV_X1 U849 ( .A(G1966), .ZN(n749) );
  AND2_X1 U850 ( .A1(n791), .A2(n749), .ZN(n777) );
  INV_X1 U851 ( .A(G8), .ZN(n750) );
  NOR2_X1 U852 ( .A1(G2084), .A2(n761), .ZN(n773) );
  OR2_X1 U853 ( .A1(n750), .A2(n773), .ZN(n751) );
  OR2_X1 U854 ( .A1(n777), .A2(n751), .ZN(n752) );
  XNOR2_X1 U855 ( .A(n752), .B(KEYINPUT30), .ZN(n753) );
  NOR2_X1 U856 ( .A1(n753), .A2(G168), .ZN(n756) );
  NOR2_X1 U857 ( .A1(G171), .A2(n754), .ZN(n755) );
  NOR2_X1 U858 ( .A1(n756), .A2(n755), .ZN(n758) );
  XNOR2_X1 U859 ( .A(n758), .B(n757), .ZN(n759) );
  NAND2_X1 U860 ( .A1(n760), .A2(n759), .ZN(n772) );
  NAND2_X1 U861 ( .A1(n772), .A2(G286), .ZN(n767) );
  INV_X1 U862 ( .A(n791), .ZN(n797) );
  NOR2_X1 U863 ( .A1(G1971), .A2(n797), .ZN(n763) );
  NOR2_X1 U864 ( .A1(G2090), .A2(n761), .ZN(n762) );
  NOR2_X1 U865 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U866 ( .A(KEYINPUT103), .B(n764), .Z(n765) );
  NAND2_X1 U867 ( .A1(n765), .A2(G303), .ZN(n766) );
  NAND2_X1 U868 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U869 ( .A(n768), .B(KEYINPUT104), .ZN(n769) );
  NAND2_X1 U870 ( .A1(n769), .A2(G8), .ZN(n771) );
  XNOR2_X1 U871 ( .A(n772), .B(KEYINPUT102), .ZN(n775) );
  NAND2_X1 U872 ( .A1(n773), .A2(G8), .ZN(n774) );
  NAND2_X1 U873 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U874 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U875 ( .A1(G166), .A2(G8), .ZN(n780) );
  NOR2_X1 U876 ( .A1(G2090), .A2(n780), .ZN(n781) );
  NOR2_X1 U877 ( .A1(n788), .A2(n781), .ZN(n782) );
  NOR2_X1 U878 ( .A1(n782), .A2(n791), .ZN(n787) );
  NOR2_X1 U879 ( .A1(G1981), .A2(G305), .ZN(n783) );
  XNOR2_X1 U880 ( .A(n783), .B(KEYINPUT96), .ZN(n784) );
  XNOR2_X1 U881 ( .A(n784), .B(KEYINPUT24), .ZN(n785) );
  AND2_X1 U882 ( .A1(n785), .A2(n791), .ZN(n786) );
  NOR2_X1 U883 ( .A1(n787), .A2(n786), .ZN(n806) );
  INV_X1 U884 ( .A(n788), .ZN(n796) );
  NOR2_X1 U885 ( .A1(G1976), .A2(G288), .ZN(n790) );
  NOR2_X1 U886 ( .A1(G1971), .A2(G303), .ZN(n789) );
  NOR2_X1 U887 ( .A1(n790), .A2(n789), .ZN(n933) );
  AND2_X1 U888 ( .A1(n790), .A2(KEYINPUT33), .ZN(n792) );
  AND2_X1 U889 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U890 ( .A(G1981), .B(G305), .ZN(n942) );
  NOR2_X1 U891 ( .A1(n793), .A2(n942), .ZN(n799) );
  AND2_X1 U892 ( .A1(n799), .A2(KEYINPUT33), .ZN(n802) );
  INV_X1 U893 ( .A(n802), .ZN(n794) );
  AND2_X1 U894 ( .A1(n933), .A2(n794), .ZN(n795) );
  NAND2_X1 U895 ( .A1(n796), .A2(n795), .ZN(n804) );
  NAND2_X1 U896 ( .A1(G1976), .A2(G288), .ZN(n937) );
  INV_X1 U897 ( .A(n937), .ZN(n798) );
  NOR2_X1 U898 ( .A1(n798), .A2(n797), .ZN(n800) );
  AND2_X1 U899 ( .A1(n800), .A2(n799), .ZN(n801) );
  OR2_X1 U900 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n805) );
  AND2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U903 ( .A(n807), .B(KEYINPUT105), .Z(n808) );
  NOR2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n811) );
  XNOR2_X1 U905 ( .A(G1986), .B(G290), .ZN(n936) );
  NAND2_X1 U906 ( .A1(n936), .A2(n823), .ZN(n810) );
  NAND2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n826) );
  NOR2_X1 U908 ( .A1(n874), .A2(G1996), .ZN(n812) );
  XNOR2_X1 U909 ( .A(n812), .B(KEYINPUT106), .ZN(n991) );
  INV_X1 U910 ( .A(n813), .ZN(n816) );
  NOR2_X1 U911 ( .A1(G1991), .A2(n878), .ZN(n982) );
  NOR2_X1 U912 ( .A1(G1986), .A2(G290), .ZN(n814) );
  NOR2_X1 U913 ( .A1(n982), .A2(n814), .ZN(n815) );
  NOR2_X1 U914 ( .A1(n816), .A2(n815), .ZN(n817) );
  NOR2_X1 U915 ( .A1(n991), .A2(n817), .ZN(n818) );
  XNOR2_X1 U916 ( .A(KEYINPUT39), .B(n818), .ZN(n820) );
  NAND2_X1 U917 ( .A1(n820), .A2(n819), .ZN(n822) );
  NAND2_X1 U918 ( .A1(n821), .A2(n897), .ZN(n993) );
  NAND2_X1 U919 ( .A1(n822), .A2(n993), .ZN(n824) );
  NAND2_X1 U920 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U922 ( .A(n827), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n828), .ZN(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U925 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U927 ( .A1(n831), .A2(n830), .ZN(G188) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  INV_X1 U931 ( .A(G69), .ZN(G235) );
  NOR2_X1 U932 ( .A1(n833), .A2(n832), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  NOR2_X1 U934 ( .A1(n834), .A2(G860), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n836), .B(n835), .ZN(G145) );
  INV_X1 U936 ( .A(n837), .ZN(G319) );
  XOR2_X1 U937 ( .A(G2100), .B(G2096), .Z(n839) );
  XNOR2_X1 U938 ( .A(KEYINPUT42), .B(G2678), .ZN(n838) );
  XNOR2_X1 U939 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U940 ( .A(KEYINPUT43), .B(G2090), .Z(n841) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2072), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U943 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U944 ( .A(G2084), .B(G2078), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(G227) );
  XOR2_X1 U946 ( .A(KEYINPUT41), .B(G1976), .Z(n847) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1971), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U949 ( .A(n848), .B(KEYINPUT109), .Z(n850) );
  XNOR2_X1 U950 ( .A(G1996), .B(G1991), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U952 ( .A(G1981), .B(G1961), .Z(n852) );
  XNOR2_X1 U953 ( .A(G1966), .B(G1956), .ZN(n851) );
  XNOR2_X1 U954 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U955 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U956 ( .A(KEYINPUT108), .B(G2474), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(G229) );
  NAND2_X1 U958 ( .A1(G124), .A2(n890), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n857), .B(KEYINPUT44), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n858), .B(KEYINPUT110), .ZN(n860) );
  NAND2_X1 U961 ( .A1(G100), .A2(n886), .ZN(n859) );
  NAND2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n864) );
  NAND2_X1 U963 ( .A1(G136), .A2(n885), .ZN(n862) );
  NAND2_X1 U964 ( .A1(G112), .A2(n891), .ZN(n861) );
  NAND2_X1 U965 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U966 ( .A1(n864), .A2(n863), .ZN(G162) );
  NAND2_X1 U967 ( .A1(G130), .A2(n890), .ZN(n866) );
  NAND2_X1 U968 ( .A1(G118), .A2(n891), .ZN(n865) );
  NAND2_X1 U969 ( .A1(n866), .A2(n865), .ZN(n873) );
  XNOR2_X1 U970 ( .A(KEYINPUT45), .B(KEYINPUT112), .ZN(n871) );
  NAND2_X1 U971 ( .A1(n885), .A2(G142), .ZN(n869) );
  NAND2_X1 U972 ( .A1(n886), .A2(G106), .ZN(n867) );
  XOR2_X1 U973 ( .A(KEYINPUT111), .B(n867), .Z(n868) );
  NAND2_X1 U974 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U975 ( .A(n871), .B(n870), .Z(n872) );
  NOR2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n884) );
  XOR2_X1 U977 ( .A(n874), .B(n980), .Z(n882) );
  XOR2_X1 U978 ( .A(KEYINPUT114), .B(KEYINPUT48), .Z(n876) );
  XNOR2_X1 U979 ( .A(KEYINPUT115), .B(KEYINPUT46), .ZN(n875) );
  XNOR2_X1 U980 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U981 ( .A(n877), .B(G162), .Z(n880) );
  XOR2_X1 U982 ( .A(G164), .B(n878), .Z(n879) );
  XNOR2_X1 U983 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U984 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n884), .B(n883), .ZN(n899) );
  NAND2_X1 U986 ( .A1(G139), .A2(n885), .ZN(n888) );
  NAND2_X1 U987 ( .A1(G103), .A2(n886), .ZN(n887) );
  NAND2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U989 ( .A(KEYINPUT113), .B(n889), .Z(n896) );
  NAND2_X1 U990 ( .A1(G127), .A2(n890), .ZN(n893) );
  NAND2_X1 U991 ( .A1(G115), .A2(n891), .ZN(n892) );
  NAND2_X1 U992 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U993 ( .A(KEYINPUT47), .B(n894), .Z(n895) );
  NOR2_X1 U994 ( .A1(n896), .A2(n895), .ZN(n975) );
  XNOR2_X1 U995 ( .A(n897), .B(n975), .ZN(n898) );
  XNOR2_X1 U996 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U997 ( .A(n900), .B(G160), .Z(n901) );
  NOR2_X1 U998 ( .A1(G37), .A2(n901), .ZN(G395) );
  XNOR2_X1 U999 ( .A(G286), .B(n929), .ZN(n906) );
  XNOR2_X1 U1000 ( .A(n902), .B(G171), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n907), .ZN(G397) );
  XOR2_X1 U1004 ( .A(KEYINPUT107), .B(G2446), .Z(n909) );
  XNOR2_X1 U1005 ( .A(G2435), .B(G2438), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n916) );
  XOR2_X1 U1007 ( .A(G2451), .B(G2430), .Z(n911) );
  XNOR2_X1 U1008 ( .A(G2454), .B(G2427), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1010 ( .A(n912), .B(G2443), .Z(n914) );
  XNOR2_X1 U1011 ( .A(G1341), .B(G1348), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(n914), .B(n913), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(n916), .B(n915), .ZN(n917) );
  NAND2_X1 U1014 ( .A1(n917), .A2(G14), .ZN(n923) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n923), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(G227), .A2(G229), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(KEYINPUT49), .B(n918), .ZN(n919) );
  NOR2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n922) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n921) );
  NAND2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(G108), .ZN(G238) );
  INV_X1 U1023 ( .A(n923), .ZN(G401) );
  XOR2_X1 U1024 ( .A(G16), .B(KEYINPUT56), .Z(n949) );
  XNOR2_X1 U1025 ( .A(n924), .B(G1348), .ZN(n927) );
  XNOR2_X1 U1026 ( .A(G1961), .B(KEYINPUT121), .ZN(n925) );
  XNOR2_X1 U1027 ( .A(n925), .B(G301), .ZN(n926) );
  NAND2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1029 ( .A(n928), .B(KEYINPUT122), .ZN(n947) );
  NAND2_X1 U1030 ( .A1(G1971), .A2(G303), .ZN(n931) );
  XOR2_X1 U1031 ( .A(G1341), .B(n929), .Z(n930) );
  NAND2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n940) );
  XNOR2_X1 U1033 ( .A(n932), .B(G1956), .ZN(n934) );
  NAND2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n938) );
  NAND2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n945) );
  XOR2_X1 U1038 ( .A(G168), .B(G1966), .Z(n941) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1040 ( .A(KEYINPUT57), .B(n943), .Z(n944) );
  NAND2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n974) );
  XNOR2_X1 U1044 ( .A(G1996), .B(G32), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(G33), .B(G2072), .ZN(n950) );
  NOR2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n956) );
  XOR2_X1 U1047 ( .A(G25), .B(G1991), .Z(n952) );
  NAND2_X1 U1048 ( .A1(n952), .A2(G28), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(G26), .B(G2067), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n959) );
  XOR2_X1 U1052 ( .A(G27), .B(n957), .Z(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1054 ( .A(KEYINPUT53), .B(n960), .Z(n964) );
  XNOR2_X1 U1055 ( .A(KEYINPUT54), .B(G34), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(n961), .B(KEYINPUT119), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(G2084), .B(n962), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(KEYINPUT118), .B(G2090), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(G35), .B(n965), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1062 ( .A(KEYINPUT55), .B(n968), .ZN(n970) );
  INV_X1 U1063 ( .A(G29), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n971), .A2(G11), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(KEYINPUT120), .B(n972), .ZN(n973) );
  NOR2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n1005) );
  XNOR2_X1 U1068 ( .A(G2072), .B(n975), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(n976), .B(KEYINPUT117), .ZN(n978) );
  XOR2_X1 U1070 ( .A(G2078), .B(G164), .Z(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1072 ( .A(KEYINPUT50), .B(n979), .Z(n999) );
  XNOR2_X1 U1073 ( .A(G2084), .B(G160), .ZN(n989) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n985) );
  NOR2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n996) );
  XOR2_X1 U1079 ( .A(G2090), .B(G162), .Z(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1081 ( .A(KEYINPUT51), .B(n992), .Z(n994) );
  NAND2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1084 ( .A(KEYINPUT116), .B(n997), .Z(n998) );
  NOR2_X1 U1085 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1086 ( .A(KEYINPUT52), .B(n1000), .ZN(n1002) );
  INV_X1 U1087 ( .A(KEYINPUT55), .ZN(n1001) );
  NAND2_X1 U1088 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1089 ( .A1(n1003), .A2(G29), .ZN(n1004) );
  NAND2_X1 U1090 ( .A1(n1005), .A2(n1004), .ZN(n1034) );
  XNOR2_X1 U1091 ( .A(G5), .B(n1006), .ZN(n1020) );
  XNOR2_X1 U1092 ( .A(G20), .B(n1007), .ZN(n1012) );
  XNOR2_X1 U1093 ( .A(G1341), .B(G19), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(G1981), .B(G6), .ZN(n1008) );
  NOR2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1096 ( .A(KEYINPUT123), .B(n1010), .Z(n1011) );
  NAND2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1015) );
  XOR2_X1 U1098 ( .A(KEYINPUT59), .B(G1348), .Z(n1013) );
  XNOR2_X1 U1099 ( .A(G4), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1101 ( .A(KEYINPUT60), .B(n1016), .Z(n1018) );
  XNOR2_X1 U1102 ( .A(G1966), .B(G21), .ZN(n1017) );
  NOR2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1105 ( .A(KEYINPUT124), .B(n1021), .ZN(n1030) );
  XNOR2_X1 U1106 ( .A(G1986), .B(G24), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(G22), .B(G1971), .ZN(n1022) );
  NOR2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1026) );
  XNOR2_X1 U1109 ( .A(G1976), .B(KEYINPUT125), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(n1024), .B(G23), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1112 ( .A(KEYINPUT58), .B(n1027), .Z(n1028) );
  XOR2_X1 U1113 ( .A(KEYINPUT126), .B(n1028), .Z(n1029) );
  NOR2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1115 ( .A(KEYINPUT61), .B(n1031), .Z(n1032) );
  NOR2_X1 U1116 ( .A1(G16), .A2(n1032), .ZN(n1033) );
  NOR2_X1 U1117 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1118 ( .A(n1035), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

