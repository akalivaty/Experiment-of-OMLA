//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n548, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n610, new_n612,
    new_n613, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1139, new_n1140;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XNOR2_X1  g016(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n463), .A3(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n461), .A2(new_n463), .A3(G137), .ZN(new_n467));
  NAND2_X1  g042(.A1(G101), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(G160));
  OAI21_X1  g045(.A(G2104), .B1(new_n459), .B2(G112), .ZN(new_n471));
  INV_X1    g046(.A(G100), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n471), .B1(new_n472), .B2(new_n459), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n473), .B(KEYINPUT65), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n461), .A2(new_n463), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(new_n459), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n475), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n474), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(new_n459), .B2(G114), .ZN(new_n483));
  NOR2_X1   g058(.A1(G102), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OR2_X1    g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n486), .A2(new_n488), .A3(KEYINPUT66), .A4(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g065(.A(KEYINPUT3), .B(G2104), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT67), .B(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n491), .A2(new_n492), .A3(G138), .A4(new_n459), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n459), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n491), .A2(G126), .A3(G2105), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n490), .A2(new_n493), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n485), .A2(new_n489), .B1(new_n494), .B2(new_n496), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n502), .A2(KEYINPUT68), .A3(new_n498), .A4(new_n493), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  XNOR2_X1  g080(.A(KEYINPUT5), .B(G543), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G50), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n514), .B(new_n516), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n511), .A2(new_n512), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n509), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n526), .B2(new_n519), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT69), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n527), .B(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n530));
  INV_X1    g105(.A(new_n511), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G51), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  AOI22_X1  g109(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n508), .ZN(new_n536));
  INV_X1    g111(.A(G52), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n511), .A2(new_n537), .B1(new_n519), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  AOI22_X1  g115(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n508), .ZN(new_n542));
  INV_X1    g117(.A(G43), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT70), .B(G81), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n511), .A2(new_n543), .B1(new_n519), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(G188));
  NAND3_X1  g127(.A1(new_n531), .A2(KEYINPUT71), .A3(G53), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT71), .ZN(new_n554));
  INV_X1    g129(.A(G53), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n511), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n553), .A2(KEYINPUT9), .A3(new_n556), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(new_n508), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n519), .A2(KEYINPUT72), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n506), .A2(new_n510), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G91), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n557), .A2(new_n558), .A3(new_n560), .A4(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  NAND2_X1  g142(.A1(new_n564), .A2(G87), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n531), .A2(G49), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  NAND3_X1  g146(.A1(new_n510), .A2(G48), .A3(G543), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(new_n564), .B2(G86), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n506), .B2(G61), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT73), .B1(new_n577), .B2(new_n508), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n514), .A2(new_n516), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n575), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT73), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n581), .A2(new_n582), .A3(G651), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n574), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G305));
  NAND2_X1  g161(.A1(new_n531), .A2(G47), .ZN(new_n587));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OAI221_X1 g164(.A(new_n587), .B1(new_n588), .B2(new_n519), .C1(new_n508), .C2(new_n589), .ZN(G290));
  INV_X1    g165(.A(G868), .ZN(new_n591));
  NOR2_X1   g166(.A1(G171), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n564), .A2(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n579), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(G54), .A2(new_n531), .B1(new_n599), .B2(G651), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n593), .B1(new_n602), .B2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(KEYINPUT74), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(KEYINPUT74), .B2(new_n592), .ZN(G284));
  OAI21_X1  g180(.A(new_n604), .B1(KEYINPUT74), .B2(new_n592), .ZN(G321));
  NAND2_X1  g181(.A1(G299), .A2(new_n591), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G168), .B2(new_n591), .ZN(G280));
  XOR2_X1   g183(.A(G280), .B(KEYINPUT75), .Z(G297));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n602), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n602), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n546), .ZN(G323));
  XOR2_X1   g189(.A(G323), .B(KEYINPUT76), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g191(.A1(new_n459), .A2(G111), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT77), .Z(new_n618));
  OAI211_X1 g193(.A(new_n618), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n619));
  AOI22_X1  g194(.A1(G123), .A2(new_n476), .B1(new_n478), .B2(G135), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND3_X1  g197(.A1(new_n459), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2100), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n622), .A2(new_n626), .ZN(G156));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2435), .ZN(new_n629));
  XOR2_X1   g204(.A(G2427), .B(G2438), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(KEYINPUT14), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2451), .B(G2454), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n632), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2443), .B(G2446), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT79), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(G14), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n638), .B2(new_n639), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n641), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(G401));
  XOR2_X1   g222(.A(G2072), .B(G2078), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT17), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XOR2_X1   g225(.A(G2067), .B(G2678), .Z(new_n651));
  NAND3_X1  g226(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT80), .ZN(new_n653));
  INV_X1    g228(.A(new_n650), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n648), .A2(new_n651), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n654), .B(new_n655), .C1(new_n649), .C2(new_n651), .ZN(new_n656));
  NOR3_X1   g231(.A1(new_n654), .A2(new_n648), .A3(new_n651), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT18), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n653), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2096), .B(G2100), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(G227));
  XNOR2_X1  g238(.A(G1961), .B(G1966), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT83), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT84), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n665), .A2(new_n666), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n673), .A2(new_n670), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT20), .Z(new_n675));
  NAND3_X1  g250(.A1(new_n668), .A2(new_n673), .A3(new_n670), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n672), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1991), .B(G1996), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT22), .B(G1981), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G229));
  INV_X1    g259(.A(KEYINPUT36), .ZN(new_n685));
  MUX2_X1   g260(.A(G24), .B(G290), .S(G16), .Z(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(G1986), .Z(new_n687));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G25), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n476), .A2(G119), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n478), .A2(G131), .ZN(new_n691));
  OR2_X1    g266(.A1(G95), .A2(G2105), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n692), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n690), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n689), .B1(new_n695), .B2(new_n688), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT35), .B(G1991), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n687), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G6), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(new_n585), .B2(new_n701), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT32), .B(G1981), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n701), .A2(G22), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G166), .B2(new_n701), .ZN(new_n707));
  INV_X1    g282(.A(G1971), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT85), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G16), .B2(G23), .ZN(new_n711));
  OR3_X1    g286(.A1(new_n710), .A2(G16), .A3(G23), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n711), .B(new_n712), .C1(G288), .C2(new_n701), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT33), .B(G1976), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  AND3_X1   g290(.A1(new_n705), .A2(new_n709), .A3(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n716), .A2(KEYINPUT34), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(KEYINPUT34), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n700), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT86), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n685), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n720), .B2(new_n719), .ZN(new_n722));
  OR3_X1    g297(.A1(new_n719), .A2(new_n720), .A3(KEYINPUT36), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n688), .A2(G35), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G162), .B2(new_n688), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT29), .Z(new_n727));
  INV_X1    g302(.A(KEYINPUT92), .ZN(new_n728));
  INV_X1    g303(.A(G2090), .ZN(new_n729));
  OR3_X1    g304(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n728), .B1(new_n727), .B2(new_n729), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n730), .A2(new_n731), .B1(new_n729), .B2(new_n727), .ZN(new_n732));
  AOI22_X1  g307(.A1(G129), .A2(new_n476), .B1(new_n478), .B2(G141), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n734));
  NAND3_X1  g309(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT26), .Z(new_n736));
  AND3_X1   g311(.A1(new_n733), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G29), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G29), .B2(G32), .ZN(new_n739));
  MUX2_X1   g314(.A(new_n738), .B(new_n739), .S(KEYINPUT91), .Z(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT27), .B(G1996), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT25), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n478), .A2(G139), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n491), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n744), .B(new_n745), .C1(new_n459), .C2(new_n746), .ZN(new_n747));
  MUX2_X1   g322(.A(G33), .B(new_n747), .S(G29), .Z(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(G2072), .Z(new_n749));
  NOR2_X1   g324(.A1(G5), .A2(G16), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G171), .B2(G16), .ZN(new_n751));
  NOR2_X1   g326(.A1(G16), .A2(G19), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n546), .B2(G16), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT88), .B(G1341), .Z(new_n754));
  AOI22_X1  g329(.A1(G1961), .A2(new_n751), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n749), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(G28), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(G28), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n758), .A2(new_n759), .A3(new_n688), .ZN(new_n760));
  OAI221_X1 g335(.A(new_n760), .B1(new_n753), .B2(new_n754), .C1(G1961), .C2(new_n751), .ZN(new_n761));
  NOR3_X1   g336(.A1(new_n742), .A2(new_n756), .A3(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT24), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(G34), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(G34), .ZN(new_n765));
  AOI21_X1  g340(.A(G29), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G160), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(G29), .ZN(new_n768));
  INV_X1    g343(.A(G2084), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT90), .Z(new_n771));
  NAND3_X1  g346(.A1(new_n732), .A2(new_n762), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(G27), .A2(G29), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G164), .B2(G29), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(G2078), .Z(new_n775));
  NAND2_X1  g350(.A1(G168), .A2(G16), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G16), .B2(G21), .ZN(new_n777));
  INV_X1    g352(.A(G1966), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n602), .A2(G16), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G4), .B2(G16), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT87), .B(G1348), .Z(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n775), .B1(new_n777), .B2(new_n778), .C1(new_n780), .C2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n772), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n768), .A2(new_n769), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n619), .A2(G29), .A3(new_n620), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT31), .B(G11), .ZN(new_n787));
  AND3_X1   g362(.A1(new_n701), .A2(KEYINPUT23), .A3(G20), .ZN(new_n788));
  AOI21_X1  g363(.A(KEYINPUT23), .B1(new_n701), .B2(G20), .ZN(new_n789));
  AOI211_X1 g364(.A(new_n788), .B(new_n789), .C1(G299), .C2(G16), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT93), .B(G1956), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT94), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n780), .B2(new_n782), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n777), .A2(new_n778), .B1(new_n790), .B2(new_n792), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n688), .A2(G26), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n476), .A2(G128), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n478), .A2(G140), .ZN(new_n798));
  OR2_X1    g373(.A1(G104), .A2(G2105), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n799), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n796), .B1(new_n802), .B2(new_n688), .ZN(new_n803));
  MUX2_X1   g378(.A(new_n796), .B(new_n803), .S(KEYINPUT28), .Z(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT89), .B(G2067), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  AND4_X1   g381(.A1(new_n787), .A2(new_n794), .A3(new_n795), .A4(new_n806), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n784), .A2(new_n785), .A3(new_n786), .A4(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT95), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n724), .B1(new_n810), .B2(new_n811), .ZN(G311));
  AND2_X1   g387(.A1(new_n808), .A2(new_n809), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n808), .A2(new_n809), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n723), .B(new_n722), .C1(new_n813), .C2(new_n814), .ZN(G150));
  INV_X1    g390(.A(G55), .ZN(new_n816));
  INV_X1    g391(.A(G93), .ZN(new_n817));
  OAI22_X1  g392(.A1(new_n511), .A2(new_n816), .B1(new_n519), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(G80), .A2(G543), .ZN(new_n819));
  INV_X1    g394(.A(G67), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n579), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n818), .B1(G651), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT97), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G860), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT37), .Z(new_n825));
  NOR2_X1   g400(.A1(new_n601), .A2(new_n610), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n823), .A2(new_n546), .ZN(new_n829));
  INV_X1    g404(.A(new_n546), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n830), .A2(new_n822), .ZN(new_n831));
  OAI21_X1  g406(.A(KEYINPUT96), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n831), .A2(KEYINPUT96), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n828), .B(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n825), .B1(new_n835), .B2(G860), .ZN(G145));
  AND2_X1   g411(.A1(new_n478), .A2(G142), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(KEYINPUT99), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n476), .A2(G130), .ZN(new_n839));
  OR2_X1    g414(.A1(G106), .A2(G2105), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n840), .B(G2104), .C1(G118), .C2(new_n459), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n837), .A2(KEYINPUT99), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n838), .A2(new_n839), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n801), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n624), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n621), .B(new_n767), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n480), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n845), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT98), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n499), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n502), .A2(KEYINPUT98), .A3(new_n498), .A4(new_n493), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n747), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n737), .B(new_n695), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n848), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(G37), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n848), .A2(new_n855), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g435(.A(new_n823), .ZN(new_n861));
  OAI21_X1  g436(.A(KEYINPUT101), .B1(new_n861), .B2(G868), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n834), .B(new_n612), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n601), .B(G299), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT41), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n864), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(new_n868), .B2(new_n863), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT100), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  XNOR2_X1  g447(.A(G288), .B(G303), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(G290), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n585), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT42), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n869), .A2(new_n870), .A3(new_n876), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n871), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n862), .B1(new_n880), .B2(new_n591), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n869), .A2(new_n870), .A3(new_n876), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n876), .B1(new_n869), .B2(new_n870), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g459(.A(KEYINPUT101), .B(G868), .C1(new_n884), .C2(new_n871), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n881), .A2(new_n885), .ZN(G295));
  NAND2_X1  g461(.A1(new_n881), .A2(new_n885), .ZN(G331));
  XNOR2_X1  g462(.A(G286), .B(G301), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n834), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n832), .A2(new_n833), .A3(new_n888), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n892), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT103), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n895), .A3(new_n865), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n888), .B1(new_n832), .B2(new_n833), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n868), .ZN(new_n899));
  INV_X1    g474(.A(new_n875), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n857), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n900), .B1(new_n896), .B2(new_n899), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT43), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n864), .B1(new_n893), .B2(new_n895), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n866), .A2(new_n898), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n875), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(new_n857), .A3(new_n901), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n904), .B1(KEYINPUT43), .B2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(KEYINPUT102), .B(KEYINPUT44), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OR3_X1    g486(.A1(new_n902), .A2(KEYINPUT43), .A3(new_n903), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(KEYINPUT43), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(KEYINPUT44), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n914), .ZN(G397));
  AOI21_X1  g490(.A(G1384), .B1(new_n850), .B2(new_n851), .ZN(new_n916));
  XOR2_X1   g491(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(G40), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n466), .A2(new_n469), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n921), .A2(G1996), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n737), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n923), .B(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n921), .ZN(new_n926));
  INV_X1    g501(.A(G2067), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n801), .B(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(G1996), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n928), .B1(new_n929), .B2(new_n737), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n925), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  XOR2_X1   g508(.A(new_n694), .B(new_n697), .Z(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n921), .B1(KEYINPUT106), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(KEYINPUT106), .B2(new_n935), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(G290), .B(G1986), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n938), .B1(new_n926), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G1384), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n499), .A2(G160), .A3(G40), .A4(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(G160), .A2(KEYINPUT45), .A3(G40), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n942), .A2(KEYINPUT110), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT110), .B1(new_n942), .B2(new_n943), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n501), .A2(new_n503), .A3(new_n941), .A4(new_n917), .ZN(new_n947));
  AOI21_X1  g522(.A(G1966), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT50), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n499), .A2(new_n949), .A3(new_n941), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n920), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n501), .A2(new_n941), .A3(new_n503), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n951), .B1(KEYINPUT50), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n769), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(G8), .B1(new_n948), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(G286), .A2(G8), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT120), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n957), .B(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT51), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT121), .ZN(new_n962));
  OR2_X1    g537(.A1(new_n961), .A2(KEYINPUT121), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n956), .A2(new_n960), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n959), .B1(new_n948), .B2(new_n955), .ZN(new_n965));
  INV_X1    g540(.A(G8), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n499), .A2(new_n941), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n967), .B(new_n920), .C1(new_n968), .C2(KEYINPUT45), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n942), .A2(KEYINPUT110), .A3(new_n943), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n969), .A2(new_n947), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n778), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n966), .B1(new_n972), .B2(new_n954), .ZN(new_n973));
  OAI211_X1 g548(.A(KEYINPUT121), .B(new_n961), .C1(new_n973), .C2(new_n959), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n964), .A2(new_n965), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT62), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n977));
  INV_X1    g552(.A(new_n917), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n952), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n852), .A2(KEYINPUT45), .A3(new_n941), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n980), .A3(new_n920), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n977), .B1(new_n981), .B2(G2078), .ZN(new_n982));
  OR2_X1    g557(.A1(new_n953), .A2(G1961), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n977), .A2(G2078), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n982), .B(new_n983), .C1(new_n971), .C2(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n985), .A2(G171), .ZN(new_n986));
  NAND2_X1  g561(.A1(G303), .A2(G8), .ZN(new_n987));
  XOR2_X1   g562(.A(new_n987), .B(KEYINPUT55), .Z(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n981), .A2(new_n708), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n504), .A2(new_n991), .A3(new_n949), .A4(new_n941), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT109), .B1(new_n952), .B2(KEYINPUT50), .ZN(new_n993));
  NAND2_X1  g568(.A1(G160), .A2(G40), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n499), .A2(new_n941), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n994), .B1(new_n995), .B2(KEYINPUT50), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n992), .A2(new_n729), .A3(new_n993), .A4(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n990), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n989), .B1(new_n998), .B2(new_n966), .ZN(new_n999));
  INV_X1    g574(.A(G1976), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n942), .B(G8), .C1(G288), .C2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT52), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n1004));
  INV_X1    g579(.A(G288), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1004), .B1(new_n1005), .B2(G1976), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(new_n1001), .ZN(new_n1007));
  INV_X1    g582(.A(G1981), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n574), .A2(new_n584), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G86), .ZN(new_n1010));
  OAI22_X1  g585(.A1(new_n577), .A2(new_n508), .B1(new_n1010), .B2(new_n519), .ZN(new_n1011));
  OAI21_X1  g586(.A(G1981), .B1(new_n1011), .B2(new_n573), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT49), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n942), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1016), .A2(new_n966), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1009), .A2(new_n1012), .A3(KEYINPUT49), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT108), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT108), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1015), .A2(new_n1021), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1022));
  AOI211_X1 g597(.A(new_n1003), .B(new_n1007), .C1(new_n1020), .C2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n952), .A2(KEYINPUT50), .ZN(new_n1024));
  INV_X1    g599(.A(new_n951), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(new_n729), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT107), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n953), .A2(KEYINPUT107), .A3(new_n729), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n990), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1030), .A2(G8), .A3(new_n988), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n999), .A2(new_n1023), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT62), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n964), .A2(new_n974), .A3(new_n965), .A4(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n976), .A2(new_n986), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1019), .A2(KEYINPUT108), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1022), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1005), .A2(new_n1000), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1009), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1030), .A2(G8), .A3(new_n988), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1040), .A2(new_n1017), .B1(new_n1041), .B2(new_n1023), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1035), .A2(new_n1042), .ZN(new_n1043));
  OAI22_X1  g618(.A1(new_n953), .A2(new_n781), .B1(G2067), .B2(new_n942), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT115), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n1046));
  OAI221_X1 g621(.A(new_n1046), .B1(G2067), .B2(new_n942), .C1(new_n953), .C2(new_n781), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n1047), .A3(new_n602), .ZN(new_n1048));
  XOR2_X1   g623(.A(new_n1048), .B(KEYINPUT116), .Z(new_n1049));
  NAND2_X1  g624(.A1(G299), .A2(KEYINPUT113), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1050), .B(KEYINPUT57), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n981), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT114), .B(G2072), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1054), .B(KEYINPUT56), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n992), .A2(new_n996), .A3(new_n993), .ZN(new_n1057));
  INV_X1    g632(.A(G1956), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1056), .A2(new_n1059), .A3(KEYINPUT117), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT117), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1052), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT118), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1064), .B(new_n1052), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1049), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1056), .A2(new_n1059), .A3(new_n1051), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1067), .A2(KEYINPUT61), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT60), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT60), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1045), .A2(new_n1047), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1070), .A2(new_n602), .A3(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1069), .A2(KEYINPUT60), .A3(new_n601), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1051), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(KEYINPUT61), .B2(new_n1067), .ZN(new_n1076));
  AND4_X1   g651(.A1(new_n1068), .A2(new_n1073), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1053), .A2(new_n929), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT119), .B(G1341), .Z(new_n1079));
  XNOR2_X1  g654(.A(new_n1079), .B(KEYINPUT58), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n942), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n830), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  XOR2_X1   g657(.A(new_n1082), .B(KEYINPUT59), .Z(new_n1083));
  AOI22_X1  g658(.A1(new_n1066), .A2(new_n1067), .B1(new_n1077), .B2(new_n1083), .ZN(new_n1084));
  XOR2_X1   g659(.A(G171), .B(KEYINPUT54), .Z(new_n1085));
  NAND2_X1  g660(.A1(new_n985), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n975), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1007), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1002), .B(new_n1088), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1041), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n918), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n994), .B1(new_n916), .B2(KEYINPUT45), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT122), .B(G2078), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1091), .A2(new_n1092), .A3(KEYINPUT53), .A4(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1085), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n982), .A2(new_n1094), .A3(new_n983), .A4(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1090), .A2(new_n999), .A3(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT123), .B1(new_n1087), .B2(new_n1097), .ZN(new_n1098));
  AND4_X1   g673(.A1(new_n1031), .A2(new_n999), .A3(new_n1023), .A4(new_n1096), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1099), .A2(new_n1100), .A3(new_n975), .A4(new_n1086), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1043), .B1(new_n1084), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT111), .ZN(new_n1104));
  AOI211_X1 g679(.A(new_n966), .B(G286), .C1(new_n972), .C2(new_n954), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1090), .A2(new_n1104), .A3(new_n999), .A4(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT63), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n999), .A2(new_n1023), .A3(new_n1031), .A4(new_n1105), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT111), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1106), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT112), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT112), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1106), .A2(new_n1109), .A3(new_n1112), .A4(new_n1107), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1030), .A2(G8), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1107), .B1(new_n1114), .B2(new_n989), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1090), .A2(new_n1105), .A3(new_n1115), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1111), .A2(new_n1113), .A3(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n940), .B1(new_n1103), .B2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n694), .A2(new_n697), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  OAI22_X1  g695(.A1(new_n932), .A2(new_n1120), .B1(G2067), .B2(new_n801), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(new_n926), .A3(new_n1124), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n921), .A2(G1986), .A3(G290), .ZN(new_n1126));
  XOR2_X1   g701(.A(new_n1126), .B(KEYINPUT48), .Z(new_n1127));
  NAND3_X1  g702(.A1(new_n933), .A2(new_n937), .A3(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n922), .A2(KEYINPUT46), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n922), .A2(KEYINPUT46), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n921), .B1(new_n737), .B2(new_n928), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1132), .B(KEYINPUT126), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1133), .B(new_n1134), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1125), .A2(new_n1128), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1118), .A2(new_n1136), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g712(.A(G227), .ZN(new_n1139));
  AND3_X1   g713(.A1(new_n859), .A2(new_n646), .A3(new_n1139), .ZN(new_n1140));
  NAND4_X1  g714(.A1(new_n909), .A2(G319), .A3(new_n683), .A4(new_n1140), .ZN(G225));
  INV_X1    g715(.A(G225), .ZN(G308));
endmodule


