//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT68), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n463), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  XOR2_X1   g049(.A(new_n474), .B(KEYINPUT69), .Z(new_n475));
  OAI21_X1  g050(.A(G2105), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n477), .B1(new_n464), .B2(G2104), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n466), .A2(KEYINPUT70), .A3(KEYINPUT3), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n478), .A2(new_n470), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT71), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n480), .A2(new_n481), .A3(G137), .A4(new_n482), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n478), .A2(new_n479), .A3(new_n482), .A4(new_n470), .ZN(new_n484));
  INV_X1    g059(.A(G137), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT71), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n466), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G101), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n476), .A2(new_n487), .A3(new_n489), .ZN(G160));
  OAI21_X1  g065(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G112), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n484), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G136), .ZN(new_n495));
  XNOR2_X1  g070(.A(new_n495), .B(KEYINPUT72), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n478), .A2(new_n479), .A3(G2105), .A4(new_n470), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  AOI211_X1 g073(.A(new_n493), .B(new_n496), .C1(G124), .C2(new_n498), .ZN(G162));
  INV_X1    g074(.A(G126), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n482), .A2(G114), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  OAI22_X1  g077(.A1(new_n497), .A2(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n479), .A2(new_n470), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n505));
  INV_X1    g080(.A(G138), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(G2105), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n504), .A2(new_n505), .A3(new_n478), .A4(new_n507), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n478), .A2(new_n479), .A3(new_n507), .A4(new_n470), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT73), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n508), .A2(KEYINPUT4), .A3(new_n510), .ZN(new_n511));
  NOR3_X1   g086(.A1(new_n506), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n512));
  INV_X1    g087(.A(new_n472), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n471), .B1(new_n469), .B2(new_n470), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n503), .B1(new_n511), .B2(new_n515), .ZN(G164));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT5), .B(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n517), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n526), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n521), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n518), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n517), .A2(G89), .ZN(new_n533));
  NAND2_X1  g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n531), .A2(new_n535), .ZN(G168));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n519), .A2(new_n537), .B1(new_n521), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n525), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n539), .A2(new_n541), .ZN(G171));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n532), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n525), .B1(new_n545), .B2(KEYINPUT74), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n546), .B1(KEYINPUT74), .B2(new_n545), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n517), .A2(new_n518), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n517), .A2(G543), .ZN(new_n549));
  AOI22_X1  g124(.A1(G81), .A2(new_n548), .B1(new_n549), .B2(G43), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT75), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND3_X1  g132(.A1(new_n517), .A2(G53), .A3(G543), .ZN(new_n558));
  XOR2_X1   g133(.A(new_n558), .B(KEYINPUT9), .Z(new_n559));
  AOI22_X1  g134(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G91), .ZN(new_n561));
  OAI22_X1  g136(.A1(new_n560), .A2(new_n525), .B1(new_n519), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(G299));
  INV_X1    g139(.A(G171), .ZN(G301));
  INV_X1    g140(.A(G168), .ZN(G286));
  INV_X1    g141(.A(G166), .ZN(G303));
  NAND3_X1  g142(.A1(new_n517), .A2(G49), .A3(G543), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT76), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n518), .A2(G74), .ZN(new_n570));
  AOI22_X1  g145(.A1(G651), .A2(new_n570), .B1(new_n548), .B2(G87), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(G288));
  INV_X1    g147(.A(G86), .ZN(new_n573));
  INV_X1    g148(.A(G48), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n519), .A2(new_n573), .B1(new_n521), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n518), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(new_n525), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n575), .A2(new_n577), .ZN(G305));
  INV_X1    g153(.A(G85), .ZN(new_n579));
  INV_X1    g154(.A(G47), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n519), .A2(new_n579), .B1(new_n521), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n525), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n549), .A2(G54), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n518), .A2(G66), .ZN(new_n588));
  NAND2_X1  g163(.A1(G79), .A2(G543), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n588), .A2(KEYINPUT77), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G651), .ZN(new_n591));
  AOI21_X1  g166(.A(KEYINPUT77), .B1(new_n588), .B2(new_n589), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n587), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT78), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n548), .A2(G92), .ZN(new_n595));
  XOR2_X1   g170(.A(new_n595), .B(KEYINPUT10), .Z(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n586), .B1(new_n598), .B2(G868), .ZN(G321));
  XOR2_X1   g174(.A(G321), .B(KEYINPUT79), .Z(G284));
  NAND2_X1  g175(.A1(G286), .A2(G868), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(new_n563), .B2(G868), .ZN(G297));
  OAI21_X1  g177(.A(new_n601), .B1(new_n563), .B2(G868), .ZN(G280));
  NOR2_X1   g178(.A1(new_n597), .A2(G559), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n604), .B1(G860), .B2(new_n598), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT80), .ZN(G148));
  NAND2_X1  g181(.A1(new_n547), .A2(new_n550), .ZN(new_n607));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(new_n604), .B2(new_n608), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n468), .A2(new_n472), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(new_n488), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT12), .Z(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(G2100), .Z(new_n616));
  AND2_X1   g191(.A1(new_n498), .A2(G123), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT81), .Z(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT82), .ZN(new_n620));
  INV_X1    g195(.A(G111), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n619), .A2(new_n620), .B1(new_n621), .B2(G2105), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n620), .B2(new_n619), .ZN(new_n623));
  INV_X1    g198(.A(G135), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(new_n484), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n618), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2096), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n616), .A2(new_n627), .ZN(G156));
  INV_X1    g203(.A(KEYINPUT86), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT84), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2427), .B(G2430), .Z(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT85), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2451), .B(G2454), .Z(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n639), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n629), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n639), .B(new_n642), .ZN(new_n647));
  INV_X1    g222(.A(new_n645), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(KEYINPUT86), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(G14), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n644), .B2(new_n645), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(KEYINPUT87), .B(KEYINPUT18), .Z(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT17), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  INV_X1    g237(.A(new_n655), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n662), .B1(new_n658), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2096), .B(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(new_n671), .A3(KEYINPUT88), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT88), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n669), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n670), .A2(new_n671), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(new_n673), .ZN(new_n679));
  MUX2_X1   g254(.A(new_n679), .B(new_n678), .S(new_n669), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(G1981), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT89), .B(KEYINPUT90), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n683), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  INV_X1    g263(.A(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n687), .A2(new_n690), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(G229));
  NOR2_X1   g268(.A1(G16), .A2(G23), .ZN(new_n694));
  AND3_X1   g269(.A1(new_n569), .A2(new_n571), .A3(KEYINPUT92), .ZN(new_n695));
  AOI21_X1  g270(.A(KEYINPUT92), .B1(new_n569), .B2(new_n571), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n694), .B1(new_n697), .B2(G16), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT33), .B(G1976), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G22), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G166), .B2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(G1971), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(G6), .A2(G16), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n575), .A2(new_n577), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(G16), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT32), .B(G1981), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n700), .A2(new_n705), .A3(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n698), .A2(new_n699), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(KEYINPUT34), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(KEYINPUT34), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n584), .A2(G16), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G16), .B2(G24), .ZN(new_n718));
  OAI21_X1  g293(.A(KEYINPUT93), .B1(new_n718), .B2(new_n689), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n689), .B2(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G25), .ZN(new_n722));
  INV_X1    g297(.A(G119), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n482), .A2(G107), .ZN(new_n724));
  OAI21_X1  g299(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n725));
  OAI22_X1  g300(.A1(new_n497), .A2(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n494), .B2(G131), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n722), .B1(new_n727), .B2(new_n721), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT35), .B(G1991), .Z(new_n729));
  XOR2_X1   g304(.A(new_n728), .B(new_n729), .Z(new_n730));
  OAI21_X1  g305(.A(new_n720), .B1(KEYINPUT91), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(KEYINPUT91), .B2(new_n730), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n715), .A2(new_n716), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT36), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n551), .A2(new_n701), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n701), .B2(G19), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(G1341), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n482), .A2(G103), .A3(G2104), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT25), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n494), .B2(G139), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n612), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(new_n482), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(new_n721), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n721), .B2(G33), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n749), .A2(G2072), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(G2072), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n740), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n721), .A2(G35), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G162), .B2(new_n721), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT29), .B(G2090), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G28), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(KEYINPUT30), .ZN(new_n758));
  AOI21_X1  g333(.A(G29), .B1(new_n757), .B2(KEYINPUT30), .ZN(new_n759));
  OR2_X1    g334(.A1(KEYINPUT31), .A2(G11), .ZN(new_n760));
  NAND2_X1  g335(.A1(KEYINPUT31), .A2(G11), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G171), .A2(new_n701), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G5), .B2(new_n701), .ZN(new_n764));
  INV_X1    g339(.A(G1961), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n626), .A2(G29), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n701), .A2(G20), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT23), .Z(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G299), .B2(G16), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT99), .B(G1956), .Z(new_n771));
  OAI21_X1  g346(.A(new_n767), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI211_X1 g347(.A(new_n766), .B(new_n772), .C1(new_n770), .C2(new_n771), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n764), .A2(new_n765), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n701), .A2(G21), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G168), .B2(new_n701), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1966), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n774), .B(new_n777), .C1(new_n739), .C2(G1341), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n752), .A2(new_n756), .A3(new_n773), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n701), .A2(G4), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n598), .B2(new_n701), .ZN(new_n781));
  INV_X1    g356(.A(G1348), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n721), .A2(G26), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT28), .ZN(new_n785));
  INV_X1    g360(.A(G128), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n482), .A2(G116), .ZN(new_n787));
  OAI21_X1  g362(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n788));
  OAI22_X1  g363(.A1(new_n497), .A2(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n494), .B2(G140), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(new_n721), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT94), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n791), .A2(new_n792), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n785), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G2067), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n721), .A2(G32), .ZN(new_n799));
  NAND3_X1  g374(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT26), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n802), .A2(new_n803), .B1(G105), .B2(new_n488), .ZN(new_n804));
  INV_X1    g379(.A(G129), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n497), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n494), .A2(G141), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n799), .B1(new_n808), .B2(new_n721), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT27), .B(G1996), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT97), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n809), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(G34), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(KEYINPUT24), .ZN(new_n814));
  AOI21_X1  g389(.A(G29), .B1(new_n813), .B2(KEYINPUT24), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(KEYINPUT95), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(KEYINPUT95), .B2(new_n815), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT96), .Z(new_n818));
  NAND3_X1  g393(.A1(new_n476), .A2(new_n487), .A3(new_n489), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(new_n721), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G2084), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n783), .A2(new_n798), .A3(new_n812), .A4(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(G27), .A2(G29), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(G164), .B2(G29), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT98), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G2078), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n779), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n735), .A2(new_n736), .A3(new_n827), .ZN(G150));
  INV_X1    g403(.A(G150), .ZN(G311));
  NAND2_X1  g404(.A1(new_n598), .A2(G559), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT38), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT100), .B(G55), .Z(new_n832));
  AOI22_X1  g407(.A1(G93), .A2(new_n548), .B1(new_n549), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n833), .A2(KEYINPUT101), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n833), .A2(KEYINPUT101), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(new_n525), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n836), .A2(new_n551), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n834), .B2(new_n835), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(new_n607), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n831), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT39), .ZN(new_n844));
  AOI21_X1  g419(.A(G860), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n844), .B2(new_n843), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n840), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT37), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(G145));
  INV_X1    g424(.A(G37), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT103), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT4), .ZN(new_n852));
  AND4_X1   g427(.A1(new_n478), .A2(new_n479), .A3(new_n507), .A4(new_n470), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n852), .B1(new_n853), .B2(new_n505), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n854), .A2(new_n510), .B1(new_n612), .B2(new_n512), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n851), .B1(new_n855), .B2(new_n503), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n509), .A2(KEYINPUT73), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT4), .B1(new_n509), .B2(KEYINPUT73), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n515), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n503), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(KEYINPUT103), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n862), .A2(new_n808), .ZN(new_n863));
  AOI211_X1 g438(.A(new_n851), .B(new_n503), .C1(new_n511), .C2(new_n515), .ZN(new_n864));
  AOI21_X1  g439(.A(KEYINPUT103), .B1(new_n859), .B2(new_n860), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n808), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n746), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n862), .A2(new_n808), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n866), .A2(new_n867), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n871), .A3(new_n745), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n790), .B(KEYINPUT104), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n869), .A2(new_n874), .A3(new_n872), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n498), .A2(G130), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n482), .A2(G118), .ZN(new_n880));
  OAI21_X1  g455(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(G142), .B2(new_n494), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n614), .B(new_n883), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n727), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n878), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT105), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n884), .B(new_n727), .Z(new_n888));
  NAND3_X1  g463(.A1(new_n888), .A2(new_n877), .A3(new_n876), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(G160), .B(KEYINPUT102), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(G162), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n626), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n878), .A2(KEYINPUT105), .A3(new_n885), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n890), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n886), .A2(new_n893), .A3(new_n889), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n897), .A2(KEYINPUT106), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(KEYINPUT106), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n850), .B(new_n896), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g476(.A(KEYINPUT110), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n840), .A2(new_n608), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n842), .A2(KEYINPUT107), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n842), .A2(KEYINPUT107), .ZN(new_n906));
  OAI22_X1  g481(.A1(new_n905), .A2(new_n906), .B1(G559), .B2(new_n597), .ZN(new_n907));
  INV_X1    g482(.A(new_n906), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(new_n604), .A3(new_n904), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n597), .A2(G299), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n594), .A2(new_n563), .A3(new_n596), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT41), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n911), .A2(KEYINPUT41), .A3(new_n912), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n907), .A2(new_n909), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n914), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n584), .ZN(new_n922));
  OAI21_X1  g497(.A(G290), .B1(new_n695), .B2(new_n696), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(G166), .B(new_n707), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT109), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n922), .A2(new_n921), .A3(new_n923), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n925), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n927), .B(new_n929), .C1(new_n931), .C2(new_n924), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n928), .A2(KEYINPUT109), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n920), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n934), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(new_n919), .A3(new_n914), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n902), .B(new_n903), .C1(new_n939), .C2(new_n608), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n608), .B1(new_n936), .B2(new_n938), .ZN(new_n941));
  INV_X1    g516(.A(new_n903), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT110), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(G295));
  OAI21_X1  g519(.A(new_n903), .B1(new_n939), .B2(new_n608), .ZN(G331));
  INV_X1    g520(.A(KEYINPUT112), .ZN(new_n946));
  OR3_X1    g521(.A1(G171), .A2(G168), .A3(KEYINPUT111), .ZN(new_n947));
  AOI21_X1  g522(.A(G286), .B1(KEYINPUT111), .B2(G171), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(KEYINPUT111), .B2(G171), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n839), .A2(new_n841), .A3(new_n947), .A4(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  AOI22_X1  g526(.A1(new_n839), .A2(new_n841), .B1(new_n949), .B2(new_n947), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n946), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n913), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n950), .A2(KEYINPUT112), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n952), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n950), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n958), .A2(new_n916), .A3(new_n917), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n927), .B1(new_n931), .B2(new_n924), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT113), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n958), .A2(new_n913), .ZN(new_n964));
  INV_X1    g539(.A(new_n918), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n953), .A2(new_n955), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(G37), .B1(new_n967), .B2(new_n962), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n962), .B1(new_n956), .B2(new_n959), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n963), .A2(new_n968), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n954), .A2(new_n950), .A3(new_n957), .ZN(new_n975));
  INV_X1    g550(.A(new_n955), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(new_n946), .B2(new_n958), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n975), .B(new_n962), .C1(new_n977), .C2(new_n918), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n850), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n967), .A2(new_n962), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT43), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n973), .A2(new_n974), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n975), .B1(new_n977), .B2(new_n918), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n961), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n968), .A2(new_n972), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n978), .B(new_n850), .C1(new_n969), .C2(new_n970), .ZN(new_n988));
  INV_X1    g563(.A(new_n971), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT43), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n968), .A2(KEYINPUT114), .A3(new_n984), .A4(new_n972), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n987), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n982), .B1(KEYINPUT44), .B2(new_n992), .ZN(G397));
  INV_X1    g568(.A(G1384), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT45), .B1(new_n866), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n476), .A2(new_n487), .A3(G40), .A4(new_n489), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n790), .B(G2067), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n998), .B1(new_n867), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1996), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n1003), .A2(KEYINPUT46), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(KEYINPUT46), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1001), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g581(.A(new_n1006), .B(KEYINPUT47), .Z(new_n1007));
  INV_X1    g582(.A(new_n998), .ZN(new_n1008));
  NOR2_X1   g583(.A1(G290), .A2(G1986), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1011), .A2(KEYINPUT48), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n808), .B(G1996), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n999), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n727), .B(new_n729), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n998), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n1011), .B2(KEYINPUT48), .ZN(new_n1017));
  AND4_X1   g592(.A1(new_n729), .A2(new_n1013), .A3(new_n727), .A4(new_n999), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1018), .B1(new_n797), .B2(new_n790), .ZN(new_n1019));
  OAI22_X1  g594(.A1(new_n1012), .A2(new_n1017), .B1(new_n1008), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1007), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G8), .ZN(new_n1022));
  NOR2_X1   g597(.A1(G166), .A2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g598(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n1024));
  OR2_X1    g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1023), .B1(KEYINPUT117), .B2(KEYINPUT55), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT45), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(G1384), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n864), .A2(new_n865), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(G1384), .B1(new_n859), .B2(new_n860), .ZN(new_n1033));
  OAI211_X1 g608(.A(G40), .B(G160), .C1(new_n1033), .C2(KEYINPUT45), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1028), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n859), .A2(new_n860), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n994), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n997), .B1(new_n1037), .B2(new_n1029), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n856), .A2(new_n861), .A3(new_n1030), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(KEYINPUT116), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1035), .A2(new_n704), .A3(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1036), .A2(new_n1043), .A3(new_n994), .ZN(new_n1044));
  INV_X1    g619(.A(new_n997), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1042), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n1046), .A2(G2090), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1041), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1027), .B1(new_n1048), .B2(G8), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1027), .ZN(new_n1050));
  AOI211_X1 g625(.A(new_n1022), .B(new_n1050), .C1(new_n1041), .C2(new_n1047), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n697), .A2(G1976), .ZN(new_n1052));
  INV_X1    g627(.A(G1976), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(G288), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1045), .A2(new_n1033), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(new_n1056), .A3(G8), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1056), .B1(new_n1055), .B2(G8), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1052), .B(new_n1054), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1037), .A2(new_n997), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT118), .B1(new_n1061), .B2(new_n1022), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n1057), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n707), .B(G1981), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT49), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1064), .B(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1062), .A2(new_n1057), .B1(new_n697), .B2(G1976), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1060), .B(new_n1067), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1049), .A2(new_n1051), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n1072));
  INV_X1    g647(.A(G2084), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1042), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1029), .B1(G164), .B2(G1384), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(G164), .B2(new_n1031), .ZN(new_n1077));
  OAI211_X1 g652(.A(KEYINPUT120), .B(new_n1030), .C1(new_n855), .C2(new_n503), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1075), .A2(new_n1077), .A3(new_n1078), .A4(new_n1045), .ZN(new_n1079));
  INV_X1    g654(.A(G1966), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1073), .A2(new_n1074), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1022), .B1(new_n1081), .B2(G168), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1074), .A2(new_n1073), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(G286), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1072), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1083), .A2(new_n1084), .A3(G168), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(G8), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1089), .A2(KEYINPUT51), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT62), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1046), .A2(new_n765), .ZN(new_n1092));
  INV_X1    g667(.A(G2078), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT53), .ZN(new_n1094));
  AOI21_X1  g669(.A(G2078), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1095));
  OAI221_X1 g670(.A(new_n1092), .B1(new_n1079), .B2(new_n1094), .C1(new_n1095), .C2(KEYINPUT53), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1096), .A2(G171), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1081), .A2(G168), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT51), .B1(new_n1089), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1082), .A2(new_n1072), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1071), .A2(new_n1091), .A3(new_n1097), .A4(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1070), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1066), .ZN(new_n1105));
  NOR2_X1   g680(.A1(G288), .A2(G1976), .ZN(new_n1106));
  XOR2_X1   g681(.A(new_n1106), .B(KEYINPUT119), .Z(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(G1981), .B2(G305), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1104), .A2(new_n1051), .B1(new_n1063), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1085), .A2(G8), .A3(G168), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT63), .B1(new_n1071), .B2(new_n1112), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1069), .A2(new_n1054), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1063), .A2(new_n1052), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT52), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1022), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1114), .B(new_n1116), .C1(new_n1117), .C2(new_n1027), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT63), .ZN(new_n1119));
  NOR4_X1   g694(.A1(new_n1118), .A2(new_n1119), .A3(new_n1051), .A4(new_n1111), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1103), .B(new_n1110), .C1(new_n1113), .C2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT56), .B(G2072), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1038), .A2(new_n1039), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(G1956), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1046), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n563), .B(KEYINPUT57), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1046), .A2(new_n782), .B1(new_n1061), .B2(new_n797), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1129), .B1(new_n597), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1123), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(KEYINPUT121), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1123), .A2(new_n1125), .A3(new_n1127), .A4(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1131), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1129), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1039), .A2(new_n1002), .A3(new_n1045), .A4(new_n1075), .ZN(new_n1141));
  XOR2_X1   g716(.A(KEYINPUT58), .B(G1341), .Z(new_n1142));
  NAND2_X1  g717(.A1(new_n1055), .A2(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1141), .A2(KEYINPUT122), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT122), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n551), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT59), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT59), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1148), .B(new_n551), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1129), .A2(KEYINPUT61), .A3(new_n1132), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1140), .A2(new_n1150), .A3(KEYINPUT123), .A4(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n598), .B1(new_n1130), .B2(KEYINPUT60), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g730(.A(KEYINPUT124), .B(new_n598), .C1(new_n1130), .C2(KEYINPUT60), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1130), .A2(KEYINPUT60), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1157), .B(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1152), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1151), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1161), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT123), .B1(new_n1162), .B2(new_n1140), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1137), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(KEYINPUT54), .B1(new_n1096), .B2(G171), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1092), .B1(new_n1095), .B2(KEYINPUT53), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT53), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1167), .B1(KEYINPUT126), .B2(new_n1093), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1039), .B(new_n1168), .C1(KEYINPUT126), .C2(new_n1093), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n996), .A2(KEYINPUT125), .A3(new_n1045), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1171), .B1(new_n995), .B2(new_n997), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1169), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(G171), .B1(new_n1166), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  OAI211_X1 g751(.A(KEYINPUT127), .B(G171), .C1(new_n1166), .C2(new_n1173), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1165), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  OR3_X1    g753(.A1(new_n1166), .A2(new_n1173), .A3(G171), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1096), .A2(G171), .ZN(new_n1180));
  AOI21_X1  g755(.A(KEYINPUT54), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1071), .A2(new_n1182), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n1178), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1121), .B1(new_n1164), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1010), .A2(KEYINPUT115), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n584), .A2(new_n689), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1186), .B(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1016), .B1(new_n1008), .B2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1021), .B1(new_n1185), .B2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g765(.A1(G227), .A2(new_n461), .ZN(new_n1192));
  NOR3_X1   g766(.A1(new_n691), .A2(new_n692), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g767(.A1(new_n653), .A2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g768(.A(new_n1194), .B1(new_n981), .B2(new_n973), .ZN(new_n1195));
  AND2_X1   g769(.A1(new_n1195), .A2(new_n900), .ZN(G308));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n900), .ZN(G225));
endmodule


