//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1210, new_n1211, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1259, new_n1260, new_n1261;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  AOI22_X1  g0003(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n204));
  INV_X1    g0004(.A(G87), .ZN(new_n205));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  INV_X1    g0007(.A(G264), .ZN(new_n208));
  OAI221_X1 g0008(.A(new_n204), .B1(new_n205), .B2(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  OR2_X1    g0009(.A1(new_n209), .A2(KEYINPUT65), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(KEYINPUT65), .ZN(new_n211));
  INV_X1    g0011(.A(G50), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n212), .A2(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G77), .B2(G244), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n210), .A2(new_n211), .A3(new_n217), .ZN(new_n218));
  AND2_X1   g0018(.A1(G116), .A2(G270), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n203), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT1), .Z(new_n221));
  NOR2_X1   g0021(.A1(new_n203), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n206), .B(new_n223), .C1(new_n224), .C2(new_n208), .ZN(new_n225));
  AND2_X1   g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G20), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT64), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(G50), .B1(G58), .B2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI22_X1  g0031(.A1(new_n225), .A2(KEYINPUT0), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n221), .B(new_n232), .C1(KEYINPUT0), .C2(new_n225), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT66), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G1), .A2(G13), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT16), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT7), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n255), .B1(new_n259), .B2(G20), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  AND2_X1   g0061(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n262));
  NOR2_X1   g0062(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G20), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n264), .A2(KEYINPUT7), .A3(new_n265), .A4(new_n258), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n214), .B1(new_n260), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G58), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(new_n214), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G58), .A2(G68), .ZN(new_n270));
  OAI21_X1  g0070(.A(G20), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT70), .B1(G20), .B2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NOR3_X1   g0073(.A1(KEYINPUT70), .A2(G20), .A3(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G159), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n271), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n254), .B1(new_n267), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT77), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(G33), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(new_n265), .A3(new_n257), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n214), .B1(new_n284), .B2(KEYINPUT7), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n283), .A2(new_n255), .A3(new_n265), .A4(new_n257), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n277), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n253), .B(new_n278), .C1(new_n289), .C2(new_n254), .ZN(new_n290));
  INV_X1    g0090(.A(G223), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n283), .A2(new_n257), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n213), .A2(G1698), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n293), .A2(new_n294), .B1(G33), .B2(G87), .ZN(new_n295));
  AND2_X1   g0095(.A1(G33), .A2(G41), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(new_n252), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT67), .B1(new_n296), .B2(new_n252), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT67), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G41), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n226), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G41), .ZN(new_n305));
  INV_X1    g0105(.A(G45), .ZN(new_n306));
  AOI21_X1  g0106(.A(G1), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(G274), .A3(new_n307), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n307), .A2(KEYINPUT68), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(KEYINPUT68), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n309), .A2(new_n304), .A3(G232), .A4(new_n310), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n299), .A2(G190), .A3(new_n308), .A4(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT8), .B(G58), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n251), .B(new_n252), .C1(G1), .C2(new_n265), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G13), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n317), .A2(G1), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G20), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n313), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT78), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT78), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n316), .A2(new_n323), .A3(new_n320), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT79), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n322), .A2(KEYINPUT79), .A3(new_n324), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n308), .B(new_n311), .C1(new_n295), .C2(new_n298), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G200), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n290), .A2(new_n312), .A3(new_n329), .A4(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT17), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n332), .B(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n290), .A2(new_n329), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n330), .A2(G169), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(new_n330), .ZN(new_n338));
  AND3_X1   g0138(.A1(new_n335), .A2(new_n338), .A3(KEYINPUT18), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT18), .B1(new_n335), .B2(new_n338), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n334), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n265), .B1(new_n270), .B2(new_n212), .ZN(new_n343));
  XOR2_X1   g0143(.A(new_n343), .B(KEYINPUT71), .Z(new_n344));
  INV_X1    g0144(.A(G150), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n261), .A2(G20), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  OAI22_X1  g0147(.A1(new_n275), .A2(new_n345), .B1(new_n347), .B2(new_n313), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n253), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n319), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n212), .ZN(new_n351));
  INV_X1    g0151(.A(new_n315), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G50), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n349), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT9), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n309), .A2(new_n304), .A3(new_n310), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G226), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n308), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT69), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n292), .A2(G222), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n259), .B(new_n362), .C1(new_n291), .C2(new_n292), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(new_n297), .C1(G77), .C2(new_n259), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n358), .A2(KEYINPUT69), .A3(new_n308), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n361), .A2(G190), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n356), .A2(new_n366), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n355), .A2(KEYINPUT9), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n361), .A2(new_n364), .A3(new_n365), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G200), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n367), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT10), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT10), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n367), .A2(new_n373), .A3(new_n368), .A4(new_n370), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n369), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n337), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n377), .B(new_n354), .C1(G169), .C2(new_n376), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n309), .A2(new_n304), .A3(G238), .A4(new_n310), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n379), .A2(new_n308), .ZN(new_n380));
  AND2_X1   g0180(.A1(G232), .A2(G1698), .ZN(new_n381));
  AND2_X1   g0181(.A1(KEYINPUT3), .A2(G33), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n381), .B1(new_n382), .B2(new_n256), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT73), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G33), .A2(G97), .ZN(new_n386));
  OAI211_X1 g0186(.A(G226), .B(new_n292), .C1(new_n382), .C2(new_n256), .ZN(new_n387));
  OAI211_X1 g0187(.A(KEYINPUT73), .B(new_n381), .C1(new_n382), .C2(new_n256), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n385), .A2(new_n386), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n389), .A2(KEYINPUT74), .A3(new_n297), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT74), .B1(new_n389), .B2(new_n297), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n380), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT13), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT13), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n394), .B(new_n380), .C1(new_n390), .C2(new_n391), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G190), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n251), .A2(new_n252), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n273), .A2(new_n274), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n400), .A2(G50), .B1(G20), .B2(new_n214), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n346), .A2(G77), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n399), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n403), .A2(KEYINPUT11), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n318), .A2(G20), .A3(new_n214), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT12), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n403), .A2(KEYINPUT11), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n352), .A2(G68), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n404), .A2(new_n406), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(G200), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(new_n393), .B2(new_n395), .ZN(new_n411));
  OR3_X1    g0211(.A1(new_n398), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  AND4_X1   g0212(.A1(new_n342), .A2(new_n375), .A3(new_n378), .A4(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT76), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT75), .ZN(new_n415));
  INV_X1    g0215(.A(G169), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n393), .B2(new_n395), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n393), .A2(G179), .A3(new_n395), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT14), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n415), .A2(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AND4_X1   g0220(.A1(new_n415), .A2(new_n396), .A3(new_n419), .A4(G169), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n414), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n418), .A2(new_n419), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n396), .A2(new_n415), .A3(G169), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n417), .A2(new_n415), .A3(new_n419), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(KEYINPUT76), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n422), .A2(new_n427), .A3(new_n409), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n357), .A2(G244), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n292), .A2(G232), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n259), .B(new_n430), .C1(new_n215), .C2(new_n292), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n431), .B(new_n297), .C1(G107), .C2(new_n259), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n429), .A2(new_n308), .A3(new_n432), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT72), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n337), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT72), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n433), .B(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n416), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n319), .A2(G77), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n400), .A2(new_n314), .B1(G20), .B2(G77), .ZN(new_n440));
  XOR2_X1   g0240(.A(KEYINPUT15), .B(G87), .Z(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n440), .B1(new_n442), .B2(new_n347), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n439), .B1(new_n443), .B2(new_n253), .ZN(new_n444));
  INV_X1    g0244(.A(G77), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n445), .B2(new_n315), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n435), .A2(new_n438), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n446), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n434), .B2(new_n410), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n437), .A2(new_n397), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n413), .A2(new_n428), .A3(new_n447), .A4(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n207), .B1(new_n260), .B2(new_n266), .ZN(new_n453));
  OAI21_X1  g0253(.A(G77), .B1(new_n273), .B2(new_n274), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT6), .ZN(new_n455));
  INV_X1    g0255(.A(G97), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n455), .A2(new_n456), .A3(G107), .ZN(new_n457));
  XNOR2_X1  g0257(.A(G97), .B(G107), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n457), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n454), .B1(new_n459), .B2(new_n265), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n253), .B1(new_n453), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n350), .A2(new_n456), .ZN(new_n462));
  INV_X1    g0262(.A(G1), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G33), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n253), .B1(KEYINPUT80), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT81), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT80), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n467), .A2(new_n463), .A3(G33), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n465), .A2(new_n466), .A3(new_n319), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n464), .A2(KEYINPUT80), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n399), .A2(new_n319), .A3(new_n470), .A4(new_n468), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT81), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n469), .A2(new_n472), .A3(G97), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n461), .A2(new_n462), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(G1698), .B1(new_n283), .B2(new_n257), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT4), .B1(new_n475), .B2(G244), .ZN(new_n476));
  OAI211_X1 g0276(.A(G250), .B(G1698), .C1(new_n382), .C2(new_n256), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G283), .ZN(new_n478));
  OAI211_X1 g0278(.A(KEYINPUT4), .B(new_n292), .C1(new_n382), .C2(new_n256), .ZN(new_n479));
  INV_X1    g0279(.A(G244), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n477), .B(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n297), .B1(new_n476), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n463), .A2(G45), .ZN(new_n483));
  NOR2_X1   g0283(.A1(KEYINPUT5), .A2(G41), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n304), .A2(G274), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n483), .ZN(new_n489));
  INV_X1    g0289(.A(new_n486), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(new_n484), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n304), .A2(G257), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n482), .A2(new_n397), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(G200), .B1(new_n482), .B2(new_n494), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n474), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT82), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n482), .A2(new_n494), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n416), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n482), .A2(new_n337), .A3(new_n494), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n461), .A2(new_n462), .A3(new_n473), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n474), .B(KEYINPUT82), .C1(new_n495), .C2(new_n496), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n499), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(G238), .A2(G1698), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n292), .A2(G244), .ZN(new_n508));
  AOI211_X1 g0308(.A(new_n507), .B(new_n508), .C1(new_n283), .C2(new_n257), .ZN(new_n509));
  INV_X1    g0309(.A(G116), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n261), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT85), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n283), .A2(new_n257), .ZN(new_n513));
  INV_X1    g0313(.A(new_n507), .ZN(new_n514));
  INV_X1    g0314(.A(new_n508), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT85), .ZN(new_n517));
  INV_X1    g0317(.A(new_n511), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n512), .A2(new_n297), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT83), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n206), .B1(new_n483), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n489), .A2(KEYINPUT83), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n304), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT84), .ZN(new_n525));
  XNOR2_X1  g0325(.A(new_n524), .B(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n489), .A2(KEYINPUT67), .A3(G274), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n520), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G200), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT19), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n530), .A2(new_n265), .A3(G33), .A4(G97), .ZN(new_n531));
  NOR3_X1   g0331(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n265), .B2(new_n386), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n531), .B1(new_n533), .B2(new_n530), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n513), .A2(new_n265), .A3(G68), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n536), .A2(new_n399), .B1(new_n319), .B2(new_n441), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n469), .A2(new_n472), .A3(G87), .ZN(new_n538));
  OR2_X1    g0338(.A1(new_n538), .A2(KEYINPUT87), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(KEYINPUT87), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n520), .A2(new_n526), .A3(G190), .A4(new_n527), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n529), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n528), .A2(new_n416), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n520), .A2(new_n526), .A3(new_n337), .A4(new_n527), .ZN(new_n545));
  XNOR2_X1  g0345(.A(new_n441), .B(KEYINPUT86), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n546), .A2(new_n469), .A3(new_n472), .ZN(new_n547));
  OAI221_X1 g0347(.A(new_n547), .B1(new_n319), .B2(new_n441), .C1(new_n536), .C2(new_n399), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT93), .ZN(new_n551));
  INV_X1    g0351(.A(G294), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n261), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(G250), .A2(G1698), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n283), .B2(new_n257), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n292), .A2(G257), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n553), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n551), .B1(new_n558), .B2(new_n298), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n304), .A2(G264), .A3(new_n491), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n488), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  AOI211_X1 g0362(.A(new_n556), .B(new_n554), .C1(new_n283), .C2(new_n257), .ZN(new_n563));
  OAI211_X1 g0363(.A(KEYINPUT93), .B(new_n297), .C1(new_n563), .C2(new_n553), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n559), .A2(new_n397), .A3(new_n562), .A4(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n558), .A2(new_n298), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n410), .B1(new_n566), .B2(new_n561), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n469), .A2(new_n472), .A3(G107), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n265), .A2(G107), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT25), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n318), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n205), .A2(G20), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n262), .A2(new_n263), .A3(new_n261), .ZN(new_n575));
  OAI211_X1 g0375(.A(KEYINPUT22), .B(new_n574), .C1(new_n575), .C2(new_n256), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n574), .B1(new_n382), .B2(new_n256), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT22), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT23), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n265), .B2(G107), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n577), .A2(new_n578), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n346), .A2(G116), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n576), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT24), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT24), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n576), .A2(new_n582), .A3(new_n586), .A4(new_n583), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n573), .B1(new_n588), .B2(new_n253), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n571), .B1(new_n318), .B2(new_n570), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n568), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  AOI211_X1 g0392(.A(new_n590), .B(new_n573), .C1(new_n588), .C2(new_n253), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n559), .A2(new_n562), .A3(new_n564), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n566), .A2(new_n561), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n594), .A2(G169), .B1(new_n595), .B2(G179), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n592), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n506), .A2(new_n550), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n513), .A2(G264), .A3(G1698), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT89), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n259), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n475), .A2(G257), .B1(G303), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n513), .A2(KEYINPUT89), .A3(G264), .A4(G1698), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n602), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n297), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n304), .A2(G270), .A3(new_n491), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n488), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT88), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT88), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n488), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT90), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n607), .A2(new_n613), .A3(KEYINPUT90), .ZN(new_n617));
  OR3_X1    g0417(.A1(new_n471), .A2(KEYINPUT91), .A3(new_n510), .ZN(new_n618));
  OAI21_X1  g0418(.A(KEYINPUT91), .B1(new_n471), .B2(new_n510), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n478), .B(new_n265), .C1(G33), .C2(new_n456), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n620), .B(new_n253), .C1(new_n265), .C2(G116), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT20), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n618), .A2(new_n619), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n319), .A2(G116), .ZN(new_n626));
  XNOR2_X1  g0426(.A(new_n626), .B(KEYINPUT92), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n416), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n616), .A2(new_n617), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT21), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n614), .A2(new_n337), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n625), .A2(new_n627), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n616), .A2(KEYINPUT21), .A3(new_n617), .A4(new_n628), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n631), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n616), .A2(new_n617), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(G190), .ZN(new_n638));
  INV_X1    g0438(.A(new_n633), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n638), .B(new_n639), .C1(new_n410), .C2(new_n637), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n452), .A2(new_n599), .A3(new_n641), .ZN(G372));
  INV_X1    g0442(.A(new_n378), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n428), .A2(new_n447), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n332), .B(KEYINPUT17), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n645), .A3(new_n412), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n335), .A2(new_n338), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT18), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n335), .A2(new_n338), .A3(KEYINPUT18), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n643), .B1(new_n652), .B2(new_n375), .ZN(new_n653));
  INV_X1    g0453(.A(new_n452), .ZN(new_n654));
  AND4_X1   g0454(.A1(new_n504), .A2(new_n499), .A3(new_n505), .A4(new_n592), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n631), .A2(new_n634), .A3(new_n635), .ZN(new_n656));
  INV_X1    g0456(.A(new_n596), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT94), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n589), .A2(new_n591), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT94), .B1(new_n593), .B2(new_n596), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n543), .B(new_n655), .C1(new_n656), .C2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n549), .ZN(new_n664));
  INV_X1    g0464(.A(new_n504), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n543), .A2(new_n549), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n543), .A2(new_n549), .A3(new_n665), .A4(KEYINPUT26), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n654), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n653), .A2(new_n672), .ZN(G369));
  NOR2_X1   g0473(.A1(new_n317), .A2(G20), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n463), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n639), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n656), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n641), .B2(new_n682), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  INV_X1    g0485(.A(new_n597), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n593), .B2(new_n681), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n593), .A2(new_n596), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n680), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n636), .A2(new_n680), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n686), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n662), .A2(new_n681), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n692), .A2(new_n696), .ZN(G399));
  NOR2_X1   g0497(.A1(new_n223), .A2(G41), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n532), .A2(new_n510), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(G1), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n230), .B2(new_n699), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT29), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT95), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n666), .A2(new_n706), .A3(new_n667), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n706), .B1(new_n666), .B2(new_n667), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n669), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n543), .B(new_n655), .C1(new_n656), .C2(new_n688), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(new_n549), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n705), .B1(new_n711), .B2(new_n681), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n680), .B1(new_n663), .B2(new_n670), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n713), .A2(new_n705), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n598), .A2(new_n636), .A3(new_n640), .A4(new_n681), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n528), .A2(new_n500), .A3(new_n566), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(new_n560), .A3(new_n632), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n717), .A2(new_n632), .A3(KEYINPUT30), .A4(new_n560), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n595), .A2(G179), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(new_n528), .A3(new_n500), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n720), .B(new_n721), .C1(new_n637), .C2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n680), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT31), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n724), .A2(new_n727), .A3(new_n680), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G330), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n715), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT96), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n704), .B1(new_n732), .B2(G1), .ZN(G364));
  XNOR2_X1  g0533(.A(new_n685), .B(KEYINPUT97), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n674), .A2(G45), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n699), .A2(G1), .A3(new_n736), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n735), .B(new_n737), .C1(G330), .C2(new_n684), .ZN(new_n738));
  INV_X1    g0538(.A(new_n737), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n397), .A2(new_n410), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n265), .A2(new_n337), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT100), .Z(new_n743));
  OR2_X1    g0543(.A1(new_n741), .A2(KEYINPUT99), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n741), .A2(KEYINPUT99), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G190), .A2(G200), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n743), .A2(G326), .B1(new_n748), .B2(G311), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n397), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n337), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n749), .B1(new_n552), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT101), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n265), .A2(G179), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n746), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n259), .B1(new_n758), .B2(G329), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n410), .A2(G190), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n741), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g0561(.A(KEYINPUT33), .B(G317), .Z(new_n762));
  NAND2_X1  g0562(.A1(new_n740), .A2(new_n756), .ZN(new_n763));
  XOR2_X1   g0563(.A(new_n763), .B(KEYINPUT102), .Z(new_n764));
  INV_X1    g0564(.A(G303), .ZN(new_n765));
  OAI221_X1 g0565(.A(new_n759), .B1(new_n761), .B2(new_n762), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n744), .A2(new_n750), .A3(new_n745), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n766), .B1(G322), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G283), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n756), .A2(new_n760), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n755), .B(new_n769), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n763), .A2(new_n205), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n758), .A2(G159), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT32), .ZN(new_n775));
  INV_X1    g0575(.A(new_n761), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n775), .B1(G68), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n742), .ZN(new_n778));
  INV_X1    g0578(.A(new_n771), .ZN(new_n779));
  AOI22_X1  g0579(.A1(G50), .A2(new_n778), .B1(new_n779), .B2(G107), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(new_n268), .B2(new_n767), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(G77), .B2(new_n748), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n753), .A2(new_n456), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n603), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n777), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n772), .B1(new_n773), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n252), .B1(G20), .B2(new_n416), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n265), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT98), .ZN(new_n790));
  INV_X1    g0590(.A(new_n787), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n513), .A2(new_n223), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n231), .A2(new_n306), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n794), .B(new_n795), .C1(new_n246), .C2(new_n306), .ZN(new_n796));
  INV_X1    g0596(.A(G355), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n259), .A2(new_n222), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n796), .B1(G116), .B2(new_n222), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n786), .A2(new_n787), .B1(new_n793), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n790), .B(KEYINPUT103), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n739), .B(new_n800), .C1(new_n684), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n738), .A2(new_n802), .ZN(G396));
  OR2_X1    g0603(.A1(new_n447), .A2(new_n680), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n449), .A2(new_n450), .B1(new_n448), .B2(new_n681), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n447), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n713), .B(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n730), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n737), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n768), .A2(G143), .B1(G150), .B2(new_n776), .ZN(new_n811));
  INV_X1    g0611(.A(G137), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n811), .B1(new_n812), .B2(new_n742), .C1(new_n276), .C2(new_n747), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT34), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n513), .B1(new_n212), .B2(new_n764), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n779), .A2(G68), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n752), .A2(G58), .B1(new_n758), .B2(G132), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n776), .A2(KEYINPUT105), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n776), .A2(KEYINPUT105), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n823), .A2(G283), .B1(G294), .B2(new_n768), .ZN(new_n824));
  INV_X1    g0624(.A(G311), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n771), .A2(new_n205), .B1(new_n757), .B2(new_n825), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n826), .B(new_n783), .C1(G303), .C2(new_n778), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n824), .B(new_n827), .C1(new_n510), .C2(new_n747), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n603), .B1(new_n764), .B2(new_n207), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT106), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n815), .A2(new_n819), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n807), .A2(new_n788), .B1(new_n787), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n787), .A2(new_n788), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n739), .B1(G77), .B2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT104), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n810), .A2(new_n837), .ZN(G384));
  INV_X1    g0638(.A(KEYINPUT40), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n428), .A2(new_n412), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n409), .A2(new_n680), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT107), .Z(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n428), .A2(new_n412), .A3(new_n842), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n807), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT38), .ZN(new_n847));
  INV_X1    g0647(.A(new_n678), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n335), .B1(new_n338), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n849), .A2(new_n850), .A3(new_n332), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n289), .A2(new_n254), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n277), .B1(new_n285), .B2(new_n286), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n399), .B1(new_n853), .B2(KEYINPUT16), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n325), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n856), .A2(KEYINPUT109), .A3(new_n848), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT109), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n852), .A2(new_n854), .B1(new_n322), .B2(new_n324), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n858), .B1(new_n859), .B2(new_n678), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n856), .A2(new_n338), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n857), .A2(new_n860), .A3(new_n861), .A4(new_n332), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n851), .B1(KEYINPUT37), .B2(new_n862), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n645), .A2(new_n651), .B1(new_n860), .B2(new_n857), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n847), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n857), .A2(new_n860), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n334), .B2(new_n341), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n862), .A2(KEYINPUT37), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n867), .B(KEYINPUT38), .C1(new_n868), .C2(new_n851), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT110), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n726), .A2(new_n871), .A3(new_n728), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(new_n726), .B2(new_n728), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n846), .B(new_n870), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n807), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n428), .A2(new_n412), .A3(new_n842), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n842), .B1(new_n428), .B2(new_n412), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n726), .A2(new_n728), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT110), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n726), .A2(new_n871), .A3(new_n728), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT111), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n335), .A2(new_n848), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n645), .B2(new_n651), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n850), .B1(new_n849), .B2(new_n332), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n851), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n847), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n869), .A2(new_n883), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n883), .B1(new_n869), .B2(new_n888), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n890), .A2(new_n891), .A3(new_n839), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n839), .A2(new_n874), .B1(new_n882), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n452), .B1(new_n880), .B2(new_n881), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n893), .B(new_n894), .Z(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(G330), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n876), .A2(new_n877), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n447), .A2(new_n680), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n713), .B2(new_n875), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT108), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n713), .A2(new_n875), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n804), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n844), .A2(new_n845), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT108), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n900), .A2(new_n905), .A3(new_n870), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n341), .A2(new_n678), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n865), .A2(new_n869), .A3(KEYINPUT39), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT39), .B1(new_n869), .B2(new_n888), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n428), .A2(new_n680), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n906), .A2(new_n907), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n654), .B1(new_n712), .B2(new_n714), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n653), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n913), .B(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n896), .B(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n463), .B2(new_n674), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT35), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n228), .B1(new_n459), .B2(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n920), .B(G116), .C1(new_n919), .C2(new_n459), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT36), .ZN(new_n922));
  OAI21_X1  g0722(.A(G77), .B1(new_n268), .B2(new_n214), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n923), .A2(new_n230), .B1(G50), .B2(new_n214), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(G1), .A3(new_n317), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n918), .A2(new_n922), .A3(new_n925), .ZN(G367));
  NAND2_X1  g0726(.A1(new_n743), .A2(G143), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n345), .B2(new_n767), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(G77), .B2(new_n779), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n822), .A2(new_n276), .B1(new_n212), .B2(new_n747), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT114), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n259), .B1(new_n763), .B2(new_n268), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n753), .A2(new_n214), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n934), .B(new_n935), .C1(G137), .C2(new_n758), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n929), .A2(new_n932), .A3(new_n933), .A4(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n822), .A2(new_n552), .ZN(new_n938));
  INV_X1    g0738(.A(new_n513), .ZN(new_n939));
  INV_X1    g0739(.A(G317), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n939), .B1(new_n940), .B2(new_n757), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT46), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n763), .B2(new_n510), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n943), .B1(new_n456), .B2(new_n771), .C1(new_n753), .C2(new_n207), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n941), .B(new_n944), .C1(G283), .C2(new_n748), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n764), .A2(new_n942), .A3(new_n510), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(G311), .B2(new_n743), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n945), .B(new_n947), .C1(new_n765), .C2(new_n767), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n937), .B1(new_n938), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT47), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n737), .B1(new_n950), .B2(new_n787), .ZN(new_n951));
  INV_X1    g0751(.A(new_n794), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n793), .B1(new_n222), .B2(new_n442), .C1(new_n241), .C2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n541), .A2(new_n681), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n664), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n550), .B2(new_n954), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n951), .B(new_n953), .C1(new_n801), .C2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n736), .A2(G1), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n693), .A2(new_n690), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n686), .B2(new_n693), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT113), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n960), .B(new_n685), .C1(KEYINPUT97), .C2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n734), .A2(KEYINPUT113), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n962), .B1(new_n963), .B2(new_n960), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n732), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n506), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n474), .B2(new_n681), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n665), .A2(new_n680), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n696), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT44), .Z(new_n973));
  NOR2_X1   g0773(.A1(new_n696), .A2(new_n971), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT45), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n692), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n966), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n732), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n698), .B(KEYINPUT41), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n958), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n694), .A2(new_n968), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT112), .ZN(new_n984));
  OR3_X1    g0784(.A1(new_n983), .A2(new_n984), .A3(KEYINPUT42), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(KEYINPUT42), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n984), .B1(new_n983), .B2(KEYINPUT42), .ZN(new_n987));
  INV_X1    g0787(.A(new_n688), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n504), .B1(new_n968), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n681), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n985), .A2(new_n986), .A3(new_n987), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n692), .A2(new_n970), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n993), .B(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n995), .B(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n957), .B1(new_n982), .B2(new_n997), .ZN(G387));
  OR2_X1    g0798(.A1(new_n732), .A2(new_n964), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n999), .A2(new_n698), .A3(new_n965), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n758), .A2(G326), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n823), .A2(G311), .B1(G317), .B2(new_n768), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n765), .B2(new_n747), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G322), .B2(new_n743), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT48), .Z(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n770), .B2(new_n753), .C1(new_n552), .C2(new_n763), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT49), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n513), .B(new_n1001), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n1007), .B2(new_n1006), .C1(new_n510), .C2(new_n771), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n546), .A2(new_n752), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n763), .A2(new_n445), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n314), .B2(new_n776), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n345), .B2(new_n757), .C1(new_n276), .C2(new_n742), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n513), .B1(new_n456), .B2(new_n771), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n212), .A2(new_n767), .B1(new_n747), .B2(new_n214), .ZN(new_n1016));
  OR4_X1    g0816(.A1(new_n1011), .A2(new_n1014), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n791), .B1(new_n1009), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n690), .A2(new_n801), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n794), .B1(new_n238), .B2(new_n306), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n701), .B2(new_n798), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n214), .A2(new_n445), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n314), .A2(new_n212), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n700), .B1(new_n1023), .B2(KEYINPUT50), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1024), .B(new_n306), .C1(KEYINPUT50), .C2(new_n1023), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1021), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n223), .A2(new_n207), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n792), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n1018), .A2(new_n1019), .A3(new_n1028), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n1029), .A2(new_n739), .B1(new_n958), .B2(new_n964), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1000), .A2(new_n1030), .ZN(G393));
  NAND2_X1  g0831(.A1(new_n978), .A2(new_n958), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n793), .B1(new_n456), .B2(new_n222), .C1(new_n249), .C2(new_n952), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n767), .A2(new_n276), .B1(new_n345), .B2(new_n742), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT51), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n758), .A2(G143), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n823), .A2(G50), .B1(new_n314), .B2(new_n748), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n763), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G68), .A2(new_n1038), .B1(new_n779), .B2(G87), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n752), .A2(G77), .ZN(new_n1040));
  AND3_X1   g0840(.A1(new_n1039), .A2(new_n513), .A3(new_n1040), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1041), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n767), .A2(new_n825), .B1(new_n940), .B2(new_n742), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT115), .Z(new_n1044));
  OR2_X1    g0844(.A1(new_n1044), .A2(KEYINPUT52), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(KEYINPUT52), .ZN(new_n1046));
  INV_X1    g0846(.A(G322), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n603), .B1(new_n757), .B2(new_n1047), .C1(new_n207), .C2(new_n771), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n822), .A2(new_n765), .B1(new_n552), .B2(new_n747), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(G116), .C2(new_n752), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1045), .A2(new_n1046), .A3(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n763), .A2(new_n770), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1042), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n737), .B1(new_n1053), .B2(new_n787), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1033), .B(new_n1054), .C1(new_n970), .C2(new_n790), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1032), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1056), .A2(KEYINPUT116), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT116), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n1032), .B2(new_n1055), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n979), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n698), .B1(new_n966), .B2(new_n978), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n1057), .A2(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(G390));
  NAND2_X1  g0862(.A1(new_n778), .A2(G283), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1063), .A2(new_n1040), .A3(new_n817), .A4(new_n603), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n764), .A2(new_n205), .B1(new_n510), .B2(new_n767), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n822), .A2(new_n207), .B1(new_n456), .B2(new_n747), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1064), .B(new_n1065), .C1(KEYINPUT121), .C2(new_n1066), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(KEYINPUT121), .B2(new_n1066), .C1(new_n552), .C2(new_n757), .ZN(new_n1068));
  XOR2_X1   g0868(.A(KEYINPUT54), .B(G143), .Z(new_n1069));
  AOI22_X1  g0869(.A1(new_n823), .A2(G137), .B1(new_n748), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1071), .A2(KEYINPUT119), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n763), .A2(new_n345), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT53), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n603), .B1(new_n758), .B2(G125), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1074), .B(new_n1075), .C1(new_n276), .C2(new_n753), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n1071), .B2(KEYINPUT119), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n779), .A2(G50), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n768), .A2(G132), .B1(G128), .B2(new_n778), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT120), .Z(new_n1080));
  NAND4_X1  g0880(.A1(new_n1072), .A2(new_n1077), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1068), .A2(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n1082), .A2(new_n791), .B1(new_n314), .B2(new_n834), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n908), .A2(new_n909), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n737), .B(new_n1083), .C1(new_n1084), .C2(new_n788), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n846), .B(G330), .C1(new_n872), .C2(new_n873), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n711), .A2(new_n681), .A3(new_n806), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1087), .A2(new_n804), .B1(new_n845), .B2(new_n844), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n869), .A2(new_n888), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(KEYINPUT111), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n889), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n911), .B(KEYINPUT117), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n1088), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n902), .A2(new_n903), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n911), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n910), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1086), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n806), .A2(new_n804), .A3(G330), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n729), .A2(new_n903), .A3(KEYINPUT118), .A4(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT118), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n726), .A2(new_n728), .A3(new_n1098), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1100), .B1(new_n897), .B2(new_n1101), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1087), .A2(new_n804), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n903), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n890), .A2(new_n891), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1092), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n897), .A2(new_n899), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1084), .B1(new_n1109), .B2(new_n911), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1103), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1097), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1085), .B1(new_n1112), .B2(new_n958), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT122), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n654), .B(G330), .C1(new_n873), .C2(new_n872), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(new_n653), .A3(new_n914), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n897), .A2(new_n1101), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1086), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n902), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1098), .B1(new_n872), .B2(new_n873), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n897), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1104), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1116), .B1(new_n1119), .B2(new_n1124), .ZN(new_n1125));
  OR2_X1    g0925(.A1(new_n1125), .A2(new_n1112), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1112), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n698), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1114), .A2(new_n1128), .ZN(G378));
  XNOR2_X1  g0929(.A(new_n1116), .B(KEYINPUT123), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n874), .A2(new_n839), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n882), .A2(new_n892), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(new_n1133), .A3(G330), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n913), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n906), .A2(new_n907), .A3(new_n912), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1136), .A2(new_n893), .A3(G330), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n375), .A2(new_n378), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT55), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n354), .A2(new_n848), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT56), .Z(new_n1141));
  XNOR2_X1  g0941(.A(new_n1139), .B(new_n1141), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1135), .A2(new_n1137), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1142), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1131), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT57), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n699), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1131), .B(KEYINPUT57), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(KEYINPUT124), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1142), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1135), .A2(new_n1137), .A3(new_n1142), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT124), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1154), .A2(new_n1155), .A3(KEYINPUT57), .A4(new_n1131), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1147), .A2(new_n1149), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1142), .A2(new_n788), .ZN(new_n1158));
  INV_X1    g0958(.A(G128), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n1159), .A2(new_n767), .B1(new_n747), .B2(new_n812), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G125), .A2(new_n778), .B1(new_n776), .B2(G132), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n345), .B2(new_n753), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1160), .B(new_n1162), .C1(new_n1038), .C2(new_n1069), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT59), .ZN(new_n1164));
  AOI21_X1  g0964(.A(G41), .B1(new_n758), .B2(G124), .ZN(new_n1165));
  AOI21_X1  g0965(.A(G33), .B1(new_n779), .B2(G159), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n778), .A2(G116), .B1(new_n758), .B2(G283), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n456), .B2(new_n761), .C1(new_n207), .C2(new_n767), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n546), .B2(new_n748), .ZN(new_n1170));
  NOR4_X1   g0970(.A1(new_n935), .A2(new_n1012), .A3(new_n513), .A4(G41), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(new_n268), .C2(new_n771), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT58), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n212), .B1(new_n575), .B2(G41), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1167), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n737), .B1(new_n1175), .B2(new_n787), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1158), .B(new_n1176), .C1(G50), .C2(new_n834), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n1154), .B2(new_n958), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1157), .A2(new_n1179), .ZN(G375));
  OAI221_X1 g0980(.A(new_n603), .B1(new_n757), .B2(new_n765), .C1(new_n445), .C2(new_n771), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1181), .B(new_n1011), .C1(G294), .C2(new_n778), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n764), .A2(new_n456), .B1(new_n207), .B2(new_n747), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G116), .B2(new_n823), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1182), .B(new_n1184), .C1(new_n770), .C2(new_n767), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n812), .A2(new_n767), .B1(new_n747), .B2(new_n345), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n764), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1186), .B1(G159), .B2(new_n1187), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n771), .A2(new_n268), .B1(new_n757), .B2(new_n1159), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n939), .B(new_n1189), .C1(G50), .C2(new_n752), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n823), .A2(new_n1069), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n778), .A2(G132), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1188), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n1185), .A2(new_n1193), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n1194), .A2(new_n791), .B1(G68), .B2(new_n834), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n737), .B(new_n1195), .C1(new_n897), .C2(new_n788), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1119), .A2(new_n1124), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1196), .B1(new_n1197), .B2(new_n958), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n981), .B(KEYINPUT125), .Z(new_n1199));
  OR2_X1    g0999(.A1(new_n1125), .A2(new_n1199), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1119), .A2(new_n1124), .A3(new_n1116), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1198), .B1(new_n1200), .B2(new_n1201), .ZN(G381));
  OR2_X1    g1002(.A1(G387), .A2(G390), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1203), .A2(G381), .ZN(new_n1204));
  OR2_X1    g1004(.A1(G393), .A2(G396), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1205), .A2(G384), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1128), .A2(new_n1113), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(G375), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1204), .A2(new_n1206), .A3(new_n1208), .ZN(G407));
  INV_X1    g1009(.A(G213), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n1208), .B2(new_n679), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(G407), .A2(new_n1211), .ZN(G409));
  XOR2_X1   g1012(.A(G393), .B(G396), .Z(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT127), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(G387), .A2(G390), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1203), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1215), .B1(new_n1203), .B2(new_n1216), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1214), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1218), .A2(new_n1214), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1157), .A2(G378), .A3(new_n1179), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT126), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1157), .A2(KEYINPUT126), .A3(G378), .A4(new_n1179), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1145), .A2(new_n1199), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1207), .B1(new_n1227), .B2(new_n1179), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1226), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n699), .B1(new_n1201), .B2(KEYINPUT60), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1125), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1231), .B(new_n1232), .C1(KEYINPUT60), .C2(new_n1201), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n1198), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(new_n810), .A3(new_n837), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1233), .A2(G384), .A3(new_n1198), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1210), .A2(G343), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1230), .A2(new_n1238), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(G2897), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1237), .B(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1228), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1243), .B1(new_n1244), .B2(new_n1239), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT62), .B1(new_n1241), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT61), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1244), .A2(new_n1237), .A3(new_n1239), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT62), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1247), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1221), .B1(new_n1246), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT61), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1248), .A2(KEYINPUT63), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT63), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1230), .A2(new_n1240), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1254), .B1(new_n1255), .B2(new_n1243), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1252), .B(new_n1253), .C1(new_n1256), .C2(new_n1248), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1251), .A2(new_n1257), .ZN(G405));
  NAND3_X1  g1058(.A1(G375), .A2(new_n1128), .A3(new_n1113), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1226), .A2(new_n1259), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(new_n1238), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1261), .B(new_n1221), .ZN(G402));
endmodule


