//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959;
  XNOR2_X1  g000(.A(G110), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G107), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT3), .A3(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT78), .B1(new_n192), .B2(G104), .ZN(new_n195));
  OR3_X1    g009(.A1(new_n192), .A2(KEYINPUT78), .A3(G104), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT4), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G101), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT79), .ZN(new_n200));
  XNOR2_X1  g014(.A(new_n199), .B(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(G101), .ZN(new_n202));
  INV_X1    g016(.A(G101), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n194), .A2(new_n203), .A3(new_n196), .A4(new_n195), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(KEYINPUT4), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n201), .A2(new_n205), .ZN(new_n206));
  XOR2_X1   g020(.A(KEYINPUT66), .B(G119), .Z(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G116), .ZN(new_n208));
  INV_X1    g022(.A(G119), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G116), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT2), .B(G113), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n208), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT66), .B(G119), .ZN(new_n215));
  INV_X1    g029(.A(G116), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n212), .B1(new_n217), .B2(new_n210), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n214), .A2(new_n218), .A3(KEYINPUT67), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n220), .B(new_n212), .C1(new_n217), .C2(new_n210), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT84), .B1(new_n206), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n219), .A2(new_n221), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT84), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n225), .A2(new_n201), .A3(new_n226), .A4(new_n205), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n208), .A2(KEYINPUT5), .A3(new_n211), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n228), .B(G113), .C1(KEYINPUT5), .C2(new_n208), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n190), .A2(G107), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n192), .A2(G104), .ZN(new_n231));
  OAI21_X1  g045(.A(G101), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n204), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n229), .A2(new_n214), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n227), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n188), .B1(new_n224), .B2(new_n235), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n223), .A2(new_n187), .A3(new_n234), .A4(new_n227), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(KEYINPUT6), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT6), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n239), .B(new_n188), .C1(new_n224), .C2(new_n235), .ZN(new_n240));
  INV_X1    g054(.A(G146), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G143), .ZN(new_n242));
  INV_X1    g056(.A(G143), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G146), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT64), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(KEYINPUT0), .A3(G128), .ZN(new_n247));
  XOR2_X1   g061(.A(KEYINPUT0), .B(G128), .Z(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT64), .A3(new_n245), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G125), .ZN(new_n251));
  INV_X1    g065(.A(G128), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n243), .A2(G146), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n241), .A2(G143), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G128), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n252), .A2(new_n253), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n252), .A2(KEYINPUT1), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(new_n242), .A3(new_n244), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G125), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n251), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G224), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(G953), .ZN(new_n265));
  XOR2_X1   g079(.A(new_n263), .B(new_n265), .Z(new_n266));
  NAND3_X1  g080(.A1(new_n238), .A2(new_n240), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT86), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT7), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n265), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n268), .B2(new_n269), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n251), .A2(new_n262), .A3(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n272), .B(KEYINPUT87), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n269), .B1(new_n265), .B2(KEYINPUT88), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n263), .B(new_n274), .C1(KEYINPUT88), .C2(new_n265), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  XOR2_X1   g090(.A(new_n187), .B(KEYINPUT8), .Z(new_n277));
  INV_X1    g091(.A(KEYINPUT85), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n234), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n229), .A2(new_n214), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n204), .A2(new_n232), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(new_n278), .A3(new_n281), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n277), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n276), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(G902), .B1(new_n286), .B2(new_n237), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n267), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(G210), .B1(G237), .B2(G902), .ZN(new_n289));
  XOR2_X1   g103(.A(new_n289), .B(KEYINPUT89), .Z(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G214), .B1(G237), .B2(G902), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n267), .A2(new_n287), .A3(new_n290), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G953), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n296), .A2(G952), .ZN(new_n297));
  NAND2_X1  g111(.A1(G234), .A2(G237), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(G902), .A3(G953), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT21), .B(G898), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n295), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G902), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT91), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(new_n261), .A3(G140), .ZN(new_n310));
  INV_X1    g124(.A(G140), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G125), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n261), .A2(G140), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n310), .B1(new_n314), .B2(new_n309), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n315), .A2(new_n241), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n314), .A2(G146), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n308), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n317), .ZN(new_n319));
  OAI211_X1 g133(.A(KEYINPUT91), .B(new_n319), .C1(new_n315), .C2(new_n241), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G237), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(new_n296), .A3(G214), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(new_n243), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n322), .A2(new_n296), .A3(G143), .A4(G214), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(KEYINPUT18), .A2(G131), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n326), .B(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n321), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT16), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n312), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n332), .B1(new_n315), .B2(new_n331), .ZN(new_n333));
  OR2_X1    g147(.A1(new_n333), .A2(G146), .ZN(new_n334));
  INV_X1    g148(.A(G131), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n326), .A2(KEYINPUT92), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT17), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT92), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n324), .A2(new_n325), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(G131), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(G131), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n336), .A2(new_n337), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n333), .A2(G146), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n339), .A2(KEYINPUT17), .A3(G131), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n334), .A2(new_n342), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(G113), .B(G122), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(new_n190), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n330), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n347), .B1(new_n330), .B2(new_n345), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n307), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G475), .ZN(new_n352));
  NOR2_X1   g166(.A1(G475), .A2(G902), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n347), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n336), .A2(new_n341), .A3(new_n340), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n343), .ZN(new_n357));
  OR3_X1    g171(.A1(new_n314), .A2(KEYINPUT93), .A3(KEYINPUT19), .ZN(new_n358));
  OAI211_X1 g172(.A(KEYINPUT19), .B(new_n310), .C1(new_n314), .C2(new_n309), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT93), .B1(new_n314), .B2(KEYINPUT19), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n358), .A2(new_n241), .A3(new_n359), .A4(new_n360), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n361), .A2(KEYINPUT94), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(KEYINPUT94), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n357), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n328), .B1(new_n320), .B2(new_n318), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n355), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI211_X1 g180(.A(KEYINPUT20), .B(new_n354), .C1(new_n366), .C2(new_n348), .ZN(new_n367));
  XOR2_X1   g181(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n368));
  NAND2_X1  g182(.A1(new_n362), .A2(new_n363), .ZN(new_n369));
  INV_X1    g183(.A(new_n357), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n365), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n348), .B1(new_n371), .B2(new_n347), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n368), .B1(new_n372), .B2(new_n353), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n352), .B1(new_n367), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT95), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g190(.A(KEYINPUT95), .B(new_n352), .C1(new_n367), .C2(new_n373), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n243), .A2(G128), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n252), .A2(G143), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G134), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n378), .A2(new_n379), .A3(G134), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT13), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n379), .A2(new_n384), .A3(G134), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n378), .A2(new_n379), .A3(new_n384), .A4(G134), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n216), .A2(G122), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT96), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n388), .B(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n216), .A2(G122), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n390), .A2(G107), .A3(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n388), .B(KEYINPUT96), .ZN(new_n393));
  INV_X1    g207(.A(new_n391), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n192), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n386), .B(new_n387), .C1(new_n392), .C2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n391), .B1(new_n393), .B2(KEYINPUT14), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT14), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n390), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n192), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n393), .A2(new_n192), .A3(new_n394), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n382), .A3(new_n383), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n396), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(KEYINPUT9), .B(G234), .ZN(new_n404));
  INV_X1    g218(.A(G217), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n404), .A2(new_n405), .A3(G953), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT97), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n396), .B(new_n406), .C1(new_n400), .C2(new_n402), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n403), .A2(KEYINPUT97), .A3(new_n407), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n307), .A3(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G478), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(KEYINPUT15), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n413), .B(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n376), .A2(new_n377), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(G221), .B1(new_n404), .B2(G902), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n260), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT10), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n421), .A2(new_n281), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT80), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n259), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n258), .A2(new_n242), .A3(new_n244), .A4(KEYINPUT80), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n425), .A2(new_n257), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT81), .B1(new_n427), .B2(new_n281), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n425), .A2(new_n257), .A3(new_n426), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT81), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n429), .A2(new_n430), .A3(new_n204), .A4(new_n232), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n423), .B1(new_n432), .B2(new_n422), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n199), .A2(new_n200), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n199), .A2(new_n200), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n250), .B(new_n205), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT11), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n438), .B1(new_n381), .B2(G137), .ZN(new_n439));
  INV_X1    g253(.A(G137), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(KEYINPUT11), .A3(G134), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n381), .A2(G137), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(G131), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n437), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(G110), .B(G140), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n296), .A2(G227), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n446), .B(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n430), .B1(new_n233), .B2(new_n429), .ZN(new_n450));
  AND4_X1   g264(.A1(new_n430), .A2(new_n429), .A3(new_n204), .A4(new_n232), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n422), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n443), .B(new_n335), .ZN(new_n453));
  INV_X1    g267(.A(new_n423), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n452), .A2(new_n436), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n445), .A2(new_n449), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n260), .B1(new_n204), .B2(new_n232), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n450), .B2(new_n451), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT82), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT12), .B1(new_n444), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(new_n444), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n457), .B1(new_n428), .B2(new_n431), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n461), .B1(new_n464), .B2(new_n453), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n466), .A2(new_n455), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n456), .B(G469), .C1(new_n467), .C2(new_n449), .ZN(new_n468));
  NAND2_X1  g282(.A1(G469), .A2(G902), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n462), .B1(new_n459), .B2(new_n444), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n464), .A2(new_n453), .A3(new_n461), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n449), .B(new_n455), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT83), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n466), .A2(KEYINPUT83), .A3(new_n449), .A4(new_n455), .ZN(new_n476));
  INV_X1    g290(.A(new_n455), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n453), .B1(new_n433), .B2(new_n436), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n448), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n475), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G469), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n481), .A3(new_n307), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n420), .B1(new_n470), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n306), .A2(new_n418), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT28), .ZN(new_n486));
  OR2_X1    g300(.A1(new_n443), .A2(G131), .ZN(new_n487));
  INV_X1    g301(.A(new_n442), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n381), .A2(G137), .ZN(new_n489));
  OAI21_X1  g303(.A(G131), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n487), .A2(new_n260), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n250), .A2(new_n444), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT68), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n247), .A2(new_n249), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(new_n453), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT68), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n225), .A2(KEYINPUT69), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT69), .B1(new_n219), .B2(new_n221), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n499), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT69), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n222), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n498), .B(new_n495), .C1(new_n505), .C2(new_n501), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n486), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT74), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI211_X1 g323(.A(new_n497), .B(new_n492), .C1(new_n500), .C2(new_n502), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT74), .B1(new_n510), .B2(KEYINPUT28), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n509), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT26), .B(G101), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n322), .A2(new_n296), .A3(G210), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT29), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(G902), .B1(new_n512), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT65), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n250), .A2(new_n444), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT65), .B1(new_n496), .B2(new_n453), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n524), .A3(new_n491), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT30), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n527), .B(new_n225), .C1(new_n499), .C2(new_n526), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n506), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n518), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT73), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n510), .A2(KEYINPUT28), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT71), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n525), .A2(new_n533), .A3(new_n225), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n506), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n533), .B1(new_n525), .B2(new_n225), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT28), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n532), .A2(new_n537), .A3(new_n517), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT73), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n529), .A2(new_n539), .A3(new_n518), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n531), .A2(new_n538), .A3(new_n519), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n521), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n532), .A2(new_n537), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n528), .A2(new_n506), .A3(new_n517), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT31), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n528), .A2(KEYINPUT31), .A3(new_n506), .A4(new_n517), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n543), .A2(new_n518), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(G472), .A2(G902), .ZN(new_n549));
  XOR2_X1   g363(.A(new_n549), .B(KEYINPUT72), .Z(new_n550));
  OAI21_X1  g364(.A(KEYINPUT32), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT32), .ZN(new_n552));
  INV_X1    g366(.A(new_n550), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n546), .A2(new_n547), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n517), .B1(new_n532), .B2(new_n537), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n552), .B(new_n553), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  AOI22_X1  g370(.A1(G472), .A2(new_n542), .B1(new_n551), .B2(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT75), .B(KEYINPUT23), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n558), .B1(new_n207), .B2(G128), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n207), .A2(G128), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT23), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n252), .A2(G119), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n559), .B(new_n560), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n562), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT24), .B(G110), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI22_X1  g380(.A1(new_n563), .A2(G110), .B1(new_n566), .B2(KEYINPUT77), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n566), .A2(KEYINPUT77), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n343), .B(new_n319), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n334), .A2(new_n343), .ZN(new_n570));
  OR2_X1    g384(.A1(new_n564), .A2(new_n565), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n563), .A2(G110), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT22), .B(G137), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n296), .A2(G221), .A3(G234), .ZN(new_n576));
  XOR2_X1   g390(.A(new_n575), .B(new_n576), .Z(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n569), .A2(new_n573), .A3(new_n577), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n307), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT25), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n581), .B(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n405), .B1(G234), .B2(new_n307), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n579), .A2(new_n580), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n584), .A2(G902), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n557), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n485), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G101), .ZN(G3));
  OAI21_X1  g406(.A(G472), .B1(new_n548), .B2(G902), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(new_n589), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n483), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n376), .A2(new_n377), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n408), .A2(KEYINPUT33), .A3(new_n410), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT98), .B(KEYINPUT33), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n411), .A2(new_n412), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT99), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n411), .A2(KEYINPUT99), .A3(new_n412), .A4(new_n602), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n601), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n414), .A2(G902), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n413), .A2(new_n414), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT100), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n413), .A2(KEYINPUT100), .A3(new_n414), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n607), .A2(new_n608), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n600), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n305), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n598), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT34), .B(G104), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  INV_X1    g432(.A(new_n373), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n354), .B1(new_n366), .B2(new_n348), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n368), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n619), .A2(KEYINPUT101), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n373), .A2(new_n623), .B1(G475), .B2(new_n351), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n305), .A2(new_n416), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n598), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT35), .B(G107), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G9));
  NOR2_X1   g443(.A1(new_n578), .A2(KEYINPUT36), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n574), .B(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n631), .A2(new_n587), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n583), .B2(new_n584), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n485), .A2(new_n594), .A3(new_n593), .A4(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT37), .B(G110), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G12));
  NOR2_X1   g451(.A1(new_n557), .A2(new_n633), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n267), .A2(new_n287), .A3(new_n290), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n290), .B1(new_n267), .B2(new_n287), .ZN(new_n640));
  INV_X1    g454(.A(new_n293), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT102), .B(G900), .Z(new_n643));
  OAI21_X1  g457(.A(new_n299), .B1(new_n643), .B2(new_n301), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n622), .A2(new_n416), .A3(new_n624), .A4(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n645), .B(KEYINPUT103), .Z(new_n646));
  NAND4_X1  g460(.A1(new_n638), .A2(new_n642), .A3(new_n483), .A4(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G128), .ZN(G30));
  INV_X1    g462(.A(KEYINPUT38), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n649), .B1(new_n639), .B2(new_n640), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n292), .A2(KEYINPUT38), .A3(new_n294), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n551), .A2(new_n556), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n529), .A2(new_n517), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n503), .A2(new_n506), .A3(new_n518), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n307), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(G472), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n600), .A2(new_n417), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n634), .A2(new_n641), .ZN(new_n660));
  AND4_X1   g474(.A1(new_n652), .A2(new_n658), .A3(new_n659), .A4(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n644), .B(KEYINPUT39), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n483), .A2(KEYINPUT40), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(KEYINPUT40), .B1(new_n483), .B2(new_n663), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n662), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n666), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n668), .A2(KEYINPUT104), .A3(new_n664), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n661), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT105), .B(G143), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G45));
  INV_X1    g486(.A(new_n613), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n599), .A3(new_n644), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n675), .A2(KEYINPUT106), .A3(new_n642), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n677), .B1(new_n674), .B2(new_n295), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n638), .A2(new_n676), .A3(new_n483), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G146), .ZN(G48));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n480), .A2(new_n307), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(G469), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(KEYINPUT107), .A3(new_n482), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n682), .A2(new_n685), .A3(G469), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n681), .B1(new_n687), .B2(new_n419), .ZN(new_n688));
  AOI211_X1 g502(.A(KEYINPUT108), .B(new_n420), .C1(new_n684), .C2(new_n686), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n590), .A3(new_n615), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NAND3_X1  g507(.A1(new_n690), .A2(new_n626), .A3(new_n590), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  NAND2_X1  g509(.A1(new_n482), .A2(KEYINPUT107), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n481), .B1(new_n480), .B2(new_n307), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n686), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n419), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT108), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n687), .A2(new_n681), .A3(new_n419), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n701), .A2(new_n642), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n701), .A2(KEYINPUT109), .A3(new_n642), .A4(new_n702), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n638), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n708), .A2(new_n304), .A3(new_n418), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n209), .ZN(G21));
  NOR2_X1   g525(.A1(new_n512), .A2(new_n517), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n553), .B1(new_n712), .B2(new_n554), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n713), .A2(new_n593), .ZN(new_n714));
  INV_X1    g528(.A(new_n589), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n659), .A2(new_n642), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n716), .A2(new_n717), .A3(new_n304), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n690), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G122), .ZN(G24));
  NAND2_X1  g534(.A1(new_n714), .A2(new_n634), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n674), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(new_n705), .B2(new_n706), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n261), .ZN(G27));
  OAI21_X1  g539(.A(new_n293), .B1(new_n639), .B2(new_n640), .ZN(new_n726));
  NOR4_X1   g540(.A1(new_n557), .A2(new_n589), .A3(new_n484), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n675), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT42), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n727), .A2(KEYINPUT42), .A3(new_n675), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n731), .B1(new_n730), .B2(new_n732), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G131), .ZN(G33));
  NAND2_X1  g550(.A1(new_n727), .A2(new_n646), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G134), .ZN(G36));
  INV_X1    g554(.A(new_n482), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n467), .A2(new_n449), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n742), .A2(new_n456), .A3(new_n743), .A4(KEYINPUT45), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n456), .B1(new_n467), .B2(new_n449), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT112), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n481), .B1(new_n745), .B2(new_n746), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n744), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n469), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT46), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n741), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(KEYINPUT46), .A3(new_n469), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n754), .A2(new_n419), .A3(new_n663), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT43), .B1(new_n599), .B2(new_n613), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n673), .A2(new_n757), .A3(new_n376), .A4(new_n377), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n633), .B1(new_n593), .B2(new_n594), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n760), .A2(new_n756), .A3(new_n758), .A4(KEYINPUT44), .ZN(new_n764));
  INV_X1    g578(.A(new_n726), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT113), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n764), .A2(KEYINPUT113), .A3(new_n765), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n755), .B(new_n763), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G137), .ZN(G39));
  NAND2_X1  g583(.A1(new_n542), .A2(G472), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n653), .ZN(new_n771));
  NOR4_X1   g585(.A1(new_n771), .A2(new_n674), .A3(new_n726), .A4(new_n715), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT47), .B1(new_n754), .B2(new_n419), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT47), .ZN(new_n774));
  AOI211_X1 g588(.A(new_n774), .B(new_n420), .C1(new_n752), .C2(new_n753), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n772), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G140), .ZN(G42));
  NAND3_X1  g591(.A1(new_n715), .A2(new_n293), .A3(new_n419), .ZN(new_n778));
  NOR4_X1   g592(.A1(new_n778), .A2(new_n658), .A3(new_n599), .A4(new_n613), .ZN(new_n779));
  INV_X1    g593(.A(new_n652), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n687), .B(KEYINPUT49), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n719), .A2(new_n691), .A3(new_n694), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n710), .A2(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n735), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT109), .B1(new_n690), .B2(new_n642), .ZN(new_n786));
  INV_X1    g600(.A(new_n706), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n722), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n679), .A2(new_n647), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n658), .A2(new_n483), .A3(new_n633), .A4(new_n644), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n788), .B(new_n790), .C1(new_n717), .C2(new_n791), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n792), .A2(KEYINPUT52), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(KEYINPUT52), .ZN(new_n794));
  INV_X1    g608(.A(new_n377), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT20), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n372), .A2(new_n796), .A3(new_n353), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n797), .B1(new_n368), .B2(new_n620), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT95), .B1(new_n798), .B2(new_n352), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n613), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n598), .A2(new_n305), .A3(new_n418), .A4(new_n800), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n635), .A2(new_n591), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n625), .A2(new_n417), .A3(new_n644), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(KEYINPUT114), .Z(new_n804));
  OAI21_X1  g618(.A(new_n723), .B1(new_n804), .B2(new_n708), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n483), .A3(new_n765), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n802), .A2(new_n806), .A3(new_n739), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n785), .A2(new_n793), .A3(new_n794), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT54), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n808), .A2(new_n809), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n730), .A2(new_n732), .ZN(new_n813));
  AOI211_X1 g627(.A(new_n809), .B(new_n813), .C1(new_n784), .C2(KEYINPUT115), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n794), .A2(new_n807), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n784), .A2(KEYINPUT115), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n814), .A2(new_n815), .A3(new_n793), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n811), .B1(KEYINPUT54), .B2(new_n818), .ZN(new_n819));
  AOI211_X1 g633(.A(new_n775), .B(new_n773), .C1(new_n420), .C2(new_n687), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n759), .A2(new_n300), .ZN(new_n821));
  OR4_X1    g635(.A1(new_n716), .A2(new_n820), .A3(new_n726), .A4(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n688), .A2(new_n689), .A3(new_n726), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n658), .A2(new_n589), .A3(new_n299), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n825), .A2(KEYINPUT117), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(KEYINPUT117), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n826), .A2(new_n600), .A3(new_n613), .A4(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n821), .A2(new_n716), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(new_n641), .A3(new_n780), .A4(new_n690), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT50), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n823), .A2(new_n300), .A3(new_n759), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n721), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n822), .A2(KEYINPUT51), .A3(new_n828), .A4(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n590), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n837), .B(KEYINPUT48), .Z(new_n838));
  NAND3_X1  g652(.A1(new_n826), .A2(new_n614), .A3(new_n827), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n707), .A2(new_n829), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n297), .A2(new_n838), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n822), .A2(KEYINPUT116), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n822), .A2(KEYINPUT116), .ZN(new_n843));
  AND4_X1   g657(.A1(new_n828), .A2(new_n842), .A3(new_n834), .A4(new_n843), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n835), .B(new_n841), .C1(new_n844), .C2(KEYINPUT51), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n819), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(G952), .A2(G953), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n782), .B1(new_n846), .B2(new_n847), .ZN(G75));
  NOR2_X1   g662(.A1(new_n296), .A2(G952), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT56), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n818), .A2(G902), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n851), .B1(new_n852), .B2(new_n291), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n238), .A2(new_n240), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(new_n266), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT55), .Z(new_n856));
  OAI21_X1  g670(.A(new_n850), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n853), .A2(new_n856), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT118), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n853), .A2(new_n860), .A3(new_n856), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n857), .B1(new_n859), .B2(new_n861), .ZN(G51));
  XOR2_X1   g676(.A(new_n818), .B(KEYINPUT54), .Z(new_n863));
  XNOR2_X1  g677(.A(new_n469), .B(KEYINPUT57), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n480), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n852), .A2(new_n749), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n849), .B1(new_n865), .B2(new_n866), .ZN(G54));
  AND4_X1   g681(.A1(KEYINPUT58), .A2(new_n818), .A3(G475), .A4(G902), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n850), .B1(new_n868), .B2(new_n372), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n372), .B2(new_n868), .ZN(G60));
  NAND2_X1  g684(.A1(G478), .A2(G902), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT59), .Z(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n607), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n850), .B1(new_n863), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n607), .B1(new_n819), .B2(new_n873), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(G63));
  NAND2_X1  g691(.A1(G217), .A2(G902), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT60), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n879), .B1(new_n812), .B2(new_n817), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n631), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n881), .B(new_n850), .C1(new_n586), .C2(new_n880), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n882), .A2(new_n883), .A3(KEYINPUT61), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT61), .B1(new_n882), .B2(new_n883), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(G66));
  OAI21_X1  g700(.A(G953), .B1(new_n303), .B2(new_n264), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n784), .A2(new_n802), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n887), .B1(new_n889), .B2(G953), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n854), .B1(G898), .B2(new_n296), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT120), .Z(new_n892));
  XNOR2_X1  g706(.A(new_n890), .B(new_n892), .ZN(G69));
  NAND2_X1  g707(.A1(new_n483), .A2(new_n663), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n557), .A2(new_n589), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n800), .A2(KEYINPUT121), .A3(new_n418), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n800), .A2(new_n418), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n726), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n895), .A2(KEYINPUT122), .A3(new_n896), .A4(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n897), .A2(new_n898), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n902), .A2(new_n896), .A3(new_n765), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n483), .A2(new_n663), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n771), .A2(new_n904), .A3(new_n715), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n901), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n900), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n768), .A2(new_n907), .A3(new_n776), .ZN(new_n908));
  INV_X1    g722(.A(new_n670), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n788), .A2(new_n909), .A3(new_n790), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n908), .B1(new_n910), .B2(KEYINPUT62), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n789), .B1(new_n707), .B2(new_n722), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT62), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n912), .A2(new_n913), .A3(new_n909), .ZN(new_n914));
  AOI21_X1  g728(.A(G953), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n527), .B1(new_n499), .B2(new_n526), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n916), .B(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT123), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n920));
  INV_X1    g734(.A(new_n918), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n913), .B1(new_n912), .B2(new_n909), .ZN(new_n922));
  NOR4_X1   g736(.A1(new_n724), .A2(KEYINPUT62), .A3(new_n670), .A4(new_n789), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n922), .A2(new_n923), .A3(new_n908), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n920), .B(new_n921), .C1(new_n924), .C2(G953), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n921), .B1(G900), .B2(G953), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n755), .A2(new_n590), .A3(new_n642), .A4(new_n659), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n739), .A2(new_n768), .A3(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n928), .A2(new_n735), .A3(new_n776), .A4(new_n912), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n926), .B1(new_n929), .B2(G953), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n919), .A2(new_n925), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n296), .B1(G227), .B2(G900), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT125), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n919), .A2(new_n925), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n919), .A2(new_n925), .A3(KEYINPUT124), .ZN(new_n938));
  INV_X1    g752(.A(new_n932), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n930), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  AND4_X1   g755(.A1(new_n934), .A2(new_n937), .A3(new_n938), .A4(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n940), .B1(new_n935), .B2(new_n936), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n934), .B1(new_n943), .B2(new_n938), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n933), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g761(.A(KEYINPUT126), .B(new_n933), .C1(new_n942), .C2(new_n944), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(G72));
  NAND2_X1  g763(.A1(new_n924), .A2(new_n889), .ZN(new_n950));
  NAND2_X1  g764(.A1(G472), .A2(G902), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT63), .Z(new_n952));
  AOI21_X1  g766(.A(new_n654), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT127), .Z(new_n954));
  NAND3_X1  g768(.A1(new_n531), .A2(new_n544), .A3(new_n540), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n810), .A2(new_n952), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n952), .B1(new_n929), .B2(new_n888), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n529), .A2(new_n517), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n849), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n954), .A2(new_n956), .A3(new_n959), .ZN(G57));
endmodule


