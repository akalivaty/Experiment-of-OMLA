

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702;

  NOR2_X1 U357 ( .A1(n578), .A2(n673), .ZN(n581) );
  XNOR2_X2 U358 ( .A(KEYINPUT68), .B(KEYINPUT3), .ZN(n431) );
  XNOR2_X2 U359 ( .A(n432), .B(n431), .ZN(n443) );
  XNOR2_X2 U360 ( .A(n445), .B(n444), .ZN(n681) );
  AND2_X1 U361 ( .A1(n342), .A2(n341), .ZN(n665) );
  AND2_X2 U362 ( .A1(n572), .A2(n571), .ZN(n669) );
  NAND2_X1 U363 ( .A1(n356), .A2(n354), .ZN(n690) );
  XNOR2_X1 U364 ( .A(n365), .B(n340), .ZN(n364) );
  AND2_X1 U365 ( .A1(n500), .A2(n367), .ZN(n366) );
  XNOR2_X1 U366 ( .A(n392), .B(n461), .ZN(n496) );
  NOR2_X1 U367 ( .A1(n639), .A2(n638), .ZN(n504) );
  XNOR2_X1 U368 ( .A(n376), .B(n447), .ZN(n689) );
  XNOR2_X1 U369 ( .A(n483), .B(n377), .ZN(n376) );
  XOR2_X1 U370 ( .A(G131), .B(KEYINPUT67), .Z(n483) );
  XNOR2_X1 U371 ( .A(G128), .B(KEYINPUT78), .ZN(n402) );
  XOR2_X1 U372 ( .A(G134), .B(G137), .Z(n377) );
  XNOR2_X2 U373 ( .A(G469), .B(n412), .ZN(n528) );
  XNOR2_X1 U374 ( .A(n359), .B(n358), .ZN(n678) );
  INV_X1 U375 ( .A(KEYINPUT45), .ZN(n358) );
  NOR2_X1 U376 ( .A1(n622), .A2(n355), .ZN(n354) );
  XNOR2_X1 U377 ( .A(n343), .B(n565), .ZN(n356) );
  INV_X1 U378 ( .A(n621), .ZN(n355) );
  INV_X1 U379 ( .A(KEYINPUT82), .ZN(n350) );
  NAND2_X1 U380 ( .A1(n364), .A2(n361), .ZN(n383) );
  INV_X1 U381 ( .A(n605), .ZN(n361) );
  XNOR2_X1 U382 ( .A(G116), .B(KEYINPUT91), .ZN(n433) );
  XOR2_X1 U383 ( .A(KEYINPUT5), .B(KEYINPUT90), .Z(n434) );
  INV_X1 U384 ( .A(n430), .ZN(n432) );
  XNOR2_X1 U385 ( .A(G113), .B(G119), .ZN(n430) );
  INV_X1 U386 ( .A(G143), .ZN(n403) );
  XNOR2_X1 U387 ( .A(G107), .B(G104), .ZN(n406) );
  XOR2_X1 U388 ( .A(KEYINPUT86), .B(G110), .Z(n407) );
  XNOR2_X1 U389 ( .A(n689), .B(n448), .ZN(n439) );
  NAND2_X1 U390 ( .A1(n334), .A2(n333), .ZN(n343) );
  XNOR2_X1 U391 ( .A(n537), .B(n536), .ZN(n566) );
  INV_X1 U392 ( .A(KEYINPUT39), .ZN(n536) );
  NOR2_X1 U393 ( .A1(n550), .A2(n535), .ZN(n537) );
  INV_X1 U394 ( .A(n625), .ZN(n535) );
  NAND2_X1 U395 ( .A1(n522), .A2(n624), .ZN(n559) );
  AND2_X1 U396 ( .A1(n374), .A2(n520), .ZN(n521) );
  XNOR2_X1 U397 ( .A(n498), .B(n497), .ZN(n501) );
  XNOR2_X1 U398 ( .A(n391), .B(n390), .ZN(n389) );
  XNOR2_X1 U399 ( .A(n456), .B(KEYINPUT19), .ZN(n394) );
  NOR2_X1 U400 ( .A1(n671), .A2(G902), .ZN(n379) );
  NAND2_X1 U401 ( .A1(n386), .A2(n384), .ZN(n571) );
  NOR2_X1 U402 ( .A1(G952), .A2(n691), .ZN(n673) );
  OR2_X1 U403 ( .A1(n678), .A2(n690), .ZN(n388) );
  NOR2_X1 U404 ( .A1(n662), .A2(G953), .ZN(n353) );
  NOR2_X1 U405 ( .A1(n508), .A2(n495), .ZN(n542) );
  XNOR2_X1 U406 ( .A(KEYINPUT4), .B(G146), .ZN(n686) );
  XNOR2_X1 U407 ( .A(G125), .B(G140), .ZN(n421) );
  XOR2_X1 U408 ( .A(G116), .B(G107), .Z(n464) );
  XNOR2_X1 U409 ( .A(G113), .B(G143), .ZN(n479) );
  XOR2_X1 U410 ( .A(G122), .B(G104), .Z(n484) );
  XNOR2_X1 U411 ( .A(n534), .B(n357), .ZN(n625) );
  XNOR2_X1 U412 ( .A(KEYINPUT38), .B(KEYINPUT71), .ZN(n357) );
  OR2_X1 U413 ( .A1(G237), .A2(G902), .ZN(n455) );
  INV_X1 U414 ( .A(n538), .ZN(n375) );
  INV_X1 U415 ( .A(KEYINPUT100), .ZN(n390) );
  AND2_X1 U416 ( .A1(n635), .A2(n527), .ZN(n378) );
  NAND2_X1 U417 ( .A1(n394), .A2(n393), .ZN(n392) );
  XNOR2_X1 U418 ( .A(n438), .B(n439), .ZN(n582) );
  XNOR2_X1 U419 ( .A(n369), .B(n368), .ZN(n418) );
  XNOR2_X1 U420 ( .A(KEYINPUT87), .B(G119), .ZN(n368) );
  XNOR2_X1 U421 ( .A(n370), .B(G110), .ZN(n369) );
  XNOR2_X1 U422 ( .A(KEYINPUT80), .B(KEYINPUT24), .ZN(n370) );
  XNOR2_X1 U423 ( .A(G128), .B(G137), .ZN(n414) );
  INV_X1 U424 ( .A(KEYINPUT2), .ZN(n387) );
  NOR2_X1 U425 ( .A1(n690), .A2(n453), .ZN(n385) );
  XNOR2_X1 U426 ( .A(n410), .B(n409), .ZN(n411) );
  INV_X1 U427 ( .A(G140), .ZN(n409) );
  XNOR2_X1 U428 ( .A(n408), .B(n397), .ZN(n410) );
  XNOR2_X1 U429 ( .A(n642), .B(n373), .ZN(n520) );
  INV_X1 U430 ( .A(KEYINPUT6), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n472), .B(n395), .ZN(n473) );
  XNOR2_X1 U432 ( .A(n371), .B(n544), .ZN(n698) );
  OR2_X1 U433 ( .A1(n658), .A2(n547), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n372), .B(n338), .ZN(n702) );
  OR2_X1 U435 ( .A1(n562), .A2(n563), .ZN(n344) );
  INV_X1 U436 ( .A(n534), .ZN(n560) );
  XNOR2_X1 U437 ( .A(n553), .B(n552), .ZN(n701) );
  NOR2_X1 U438 ( .A1(n547), .A2(n360), .ZN(n612) );
  NAND2_X1 U439 ( .A1(n367), .A2(n363), .ZN(n362) );
  INV_X1 U440 ( .A(n642), .ZN(n363) );
  XNOR2_X1 U441 ( .A(n382), .B(n381), .ZN(n672) );
  INV_X1 U442 ( .A(n673), .ZN(n341) );
  XNOR2_X1 U443 ( .A(n352), .B(n351), .ZN(G75) );
  XNOR2_X1 U444 ( .A(KEYINPUT53), .B(KEYINPUT117), .ZN(n351) );
  NAND2_X1 U445 ( .A1(n353), .A2(n336), .ZN(n352) );
  XNOR2_X1 U446 ( .A(n364), .B(G119), .ZN(G21) );
  XOR2_X1 U447 ( .A(n546), .B(n545), .Z(n333) );
  AND2_X1 U448 ( .A1(n564), .A2(n344), .ZN(n334) );
  XNOR2_X1 U449 ( .A(G110), .B(KEYINPUT16), .ZN(n335) );
  XOR2_X1 U450 ( .A(n388), .B(KEYINPUT2), .Z(n336) );
  AND2_X1 U451 ( .A1(G953), .A2(G898), .ZN(n337) );
  XOR2_X1 U452 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n338) );
  XNOR2_X1 U453 ( .A(n663), .B(KEYINPUT59), .ZN(n339) );
  XNOR2_X1 U454 ( .A(KEYINPUT64), .B(KEYINPUT32), .ZN(n340) );
  XNOR2_X1 U455 ( .A(G902), .B(KEYINPUT15), .ZN(n453) );
  NAND2_X1 U456 ( .A1(n570), .A2(n569), .ZN(n572) );
  NOR2_X1 U457 ( .A1(n559), .A2(n560), .ZN(n561) );
  XNOR2_X1 U458 ( .A(n664), .B(n339), .ZN(n342) );
  INV_X1 U459 ( .A(n344), .ZN(n619) );
  NOR2_X1 U460 ( .A1(n667), .A2(G902), .ZN(n475) );
  XNOR2_X1 U461 ( .A(n474), .B(n473), .ZN(n667) );
  NOR2_X1 U462 ( .A1(n614), .A2(n375), .ZN(n374) );
  NAND2_X1 U463 ( .A1(n345), .A2(n400), .ZN(n359) );
  XNOR2_X1 U464 ( .A(n347), .B(n346), .ZN(n345) );
  INV_X1 U465 ( .A(KEYINPUT44), .ZN(n346) );
  NAND2_X1 U466 ( .A1(n349), .A2(n348), .ZN(n347) );
  INV_X1 U467 ( .A(n700), .ZN(n348) );
  XNOR2_X1 U468 ( .A(n383), .B(n350), .ZN(n349) );
  INV_X1 U469 ( .A(n394), .ZN(n360) );
  NOR2_X2 U470 ( .A1(n512), .A2(n362), .ZN(n605) );
  NAND2_X1 U471 ( .A1(n501), .A2(n639), .ZN(n512) );
  NAND2_X1 U472 ( .A1(n501), .A2(n366), .ZN(n365) );
  INV_X1 U473 ( .A(n635), .ZN(n367) );
  NAND2_X1 U474 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U475 ( .A1(n702), .A2(n698), .ZN(n546) );
  XNOR2_X1 U476 ( .A(n543), .B(n396), .ZN(n658) );
  NAND2_X1 U477 ( .A1(n566), .A2(n611), .ZN(n372) );
  XNOR2_X2 U478 ( .A(n441), .B(n440), .ZN(n642) );
  NAND2_X1 U479 ( .A1(n380), .A2(n378), .ZN(n529) );
  XNOR2_X2 U480 ( .A(n379), .B(n427), .ZN(n635) );
  INV_X1 U481 ( .A(n528), .ZN(n380) );
  XNOR2_X1 U482 ( .A(n671), .B(n670), .ZN(n381) );
  NAND2_X1 U483 ( .A1(n669), .A2(G217), .ZN(n382) );
  NOR2_X1 U484 ( .A1(n690), .A2(n387), .ZN(n384) );
  NAND2_X1 U485 ( .A1(n386), .A2(n385), .ZN(n570) );
  INV_X1 U486 ( .A(n678), .ZN(n386) );
  NAND2_X1 U487 ( .A1(n496), .A2(n389), .ZN(n498) );
  NAND2_X1 U488 ( .A1(n542), .A2(n634), .ZN(n391) );
  NOR2_X1 U489 ( .A1(n516), .A2(n337), .ZN(n393) );
  XNOR2_X1 U490 ( .A(n452), .B(n451), .ZN(n573) );
  XNOR2_X1 U491 ( .A(n681), .B(n399), .ZN(n452) );
  XOR2_X1 U492 ( .A(n471), .B(n470), .Z(n395) );
  XNOR2_X1 U493 ( .A(KEYINPUT41), .B(KEYINPUT106), .ZN(n396) );
  AND2_X1 U494 ( .A1(G227), .A2(n691), .ZN(n397) );
  AND2_X1 U495 ( .A1(G210), .A2(n455), .ZN(n398) );
  XOR2_X1 U496 ( .A(n446), .B(KEYINPUT17), .Z(n399) );
  XNOR2_X1 U497 ( .A(KEYINPUT101), .B(n515), .ZN(n400) );
  NAND2_X1 U498 ( .A1(n701), .A2(n555), .ZN(n556) );
  INV_X1 U499 ( .A(KEYINPUT48), .ZN(n565) );
  XNOR2_X1 U500 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U501 ( .A(n439), .B(n411), .ZN(n590) );
  INV_X1 U502 ( .A(KEYINPUT63), .ZN(n586) );
  INV_X1 U503 ( .A(KEYINPUT103), .ZN(n552) );
  XNOR2_X1 U504 ( .A(n587), .B(n586), .ZN(n588) );
  INV_X1 U505 ( .A(n453), .ZN(n567) );
  XNOR2_X1 U506 ( .A(KEYINPUT1), .B(KEYINPUT65), .ZN(n413) );
  INV_X1 U507 ( .A(n402), .ZN(n401) );
  NAND2_X1 U508 ( .A1(n401), .A2(G143), .ZN(n405) );
  NAND2_X1 U509 ( .A1(n403), .A2(n402), .ZN(n404) );
  NAND2_X1 U510 ( .A1(n405), .A2(n404), .ZN(n447) );
  XNOR2_X1 U511 ( .A(G101), .B(n686), .ZN(n448) );
  XNOR2_X1 U512 ( .A(n407), .B(n406), .ZN(n408) );
  INV_X2 U513 ( .A(G953), .ZN(n691) );
  NOR2_X1 U514 ( .A1(G902), .A2(n590), .ZN(n412) );
  XNOR2_X1 U515 ( .A(n413), .B(n528), .ZN(n523) );
  INV_X1 U516 ( .A(n523), .ZN(n639) );
  XOR2_X1 U517 ( .A(KEYINPUT88), .B(KEYINPUT23), .Z(n415) );
  XNOR2_X1 U518 ( .A(n415), .B(n414), .ZN(n420) );
  NAND2_X1 U519 ( .A1(G234), .A2(n691), .ZN(n416) );
  XOR2_X1 U520 ( .A(KEYINPUT8), .B(n416), .Z(n469) );
  NAND2_X1 U521 ( .A1(G221), .A2(n469), .ZN(n417) );
  XNOR2_X1 U522 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U523 ( .A(n420), .B(n419), .ZN(n422) );
  XNOR2_X1 U524 ( .A(n421), .B(KEYINPUT10), .ZN(n687) );
  XNOR2_X1 U525 ( .A(G146), .B(n687), .ZN(n488) );
  XNOR2_X1 U526 ( .A(n422), .B(n488), .ZN(n671) );
  XOR2_X1 U527 ( .A(KEYINPUT74), .B(KEYINPUT25), .Z(n425) );
  NAND2_X1 U528 ( .A1(n453), .A2(G234), .ZN(n423) );
  XNOR2_X1 U529 ( .A(n423), .B(KEYINPUT20), .ZN(n428) );
  NAND2_X1 U530 ( .A1(n428), .A2(G217), .ZN(n424) );
  XNOR2_X1 U531 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U532 ( .A(KEYINPUT89), .B(n426), .ZN(n427) );
  NAND2_X1 U533 ( .A1(n428), .A2(G221), .ZN(n429) );
  XOR2_X1 U534 ( .A(KEYINPUT21), .B(n429), .Z(n634) );
  NAND2_X1 U535 ( .A1(n635), .A2(n634), .ZN(n638) );
  XNOR2_X1 U536 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U537 ( .A(n443), .B(n435), .Z(n437) );
  NOR2_X1 U538 ( .A1(G953), .A2(G237), .ZN(n476) );
  NAND2_X1 U539 ( .A1(n476), .A2(G210), .ZN(n436) );
  XNOR2_X1 U540 ( .A(n437), .B(n436), .ZN(n438) );
  NOR2_X1 U541 ( .A1(G902), .A2(n582), .ZN(n441) );
  XNOR2_X1 U542 ( .A(G472), .B(KEYINPUT69), .ZN(n440) );
  AND2_X1 U543 ( .A1(n504), .A2(n520), .ZN(n442) );
  XNOR2_X1 U544 ( .A(KEYINPUT33), .B(n442), .ZN(n657) );
  INV_X1 U545 ( .A(KEYINPUT0), .ZN(n461) );
  XNOR2_X1 U546 ( .A(n443), .B(n335), .ZN(n445) );
  XNOR2_X1 U547 ( .A(n464), .B(n484), .ZN(n444) );
  XNOR2_X1 U548 ( .A(G125), .B(KEYINPUT18), .ZN(n446) );
  XNOR2_X1 U549 ( .A(n448), .B(n447), .ZN(n450) );
  NAND2_X1 U550 ( .A1(G224), .A2(n691), .ZN(n449) );
  NAND2_X1 U551 ( .A1(n573), .A2(n453), .ZN(n454) );
  XNOR2_X2 U552 ( .A(n454), .B(n398), .ZN(n534) );
  NAND2_X1 U553 ( .A1(G214), .A2(n455), .ZN(n624) );
  NAND2_X1 U554 ( .A1(n534), .A2(n624), .ZN(n456) );
  NAND2_X1 U555 ( .A1(G234), .A2(G237), .ZN(n457) );
  XNOR2_X1 U556 ( .A(n457), .B(KEYINPUT14), .ZN(n623) );
  NOR2_X1 U557 ( .A1(G902), .A2(n691), .ZN(n459) );
  NOR2_X1 U558 ( .A1(G953), .A2(G952), .ZN(n458) );
  NOR2_X1 U559 ( .A1(n459), .A2(n458), .ZN(n460) );
  NAND2_X1 U560 ( .A1(n623), .A2(n460), .ZN(n516) );
  INV_X1 U561 ( .A(n496), .ZN(n505) );
  NOR2_X1 U562 ( .A1(n657), .A2(n505), .ZN(n463) );
  XNOR2_X1 U563 ( .A(KEYINPUT34), .B(KEYINPUT76), .ZN(n462) );
  XNOR2_X1 U564 ( .A(n463), .B(n462), .ZN(n493) );
  XNOR2_X1 U565 ( .A(G134), .B(n447), .ZN(n468) );
  XOR2_X1 U566 ( .A(KEYINPUT97), .B(KEYINPUT95), .Z(n466) );
  XNOR2_X1 U567 ( .A(n464), .B(KEYINPUT9), .ZN(n465) );
  XNOR2_X1 U568 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U569 ( .A(n468), .B(n467), .Z(n474) );
  NAND2_X1 U570 ( .A1(G217), .A2(n469), .ZN(n472) );
  XOR2_X1 U571 ( .A(KEYINPUT98), .B(KEYINPUT7), .Z(n471) );
  XNOR2_X1 U572 ( .A(G122), .B(KEYINPUT96), .ZN(n470) );
  XOR2_X1 U573 ( .A(G478), .B(n475), .Z(n508) );
  XNOR2_X1 U574 ( .A(KEYINPUT13), .B(G475), .ZN(n491) );
  XOR2_X1 U575 ( .A(KEYINPUT93), .B(KEYINPUT11), .Z(n478) );
  NAND2_X1 U576 ( .A1(G214), .A2(n476), .ZN(n477) );
  XNOR2_X1 U577 ( .A(n478), .B(n477), .ZN(n482) );
  XOR2_X1 U578 ( .A(KEYINPUT12), .B(KEYINPUT94), .Z(n480) );
  XNOR2_X1 U579 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U580 ( .A(n482), .B(n481), .Z(n487) );
  INV_X1 U581 ( .A(n483), .ZN(n485) );
  XOR2_X1 U582 ( .A(n485), .B(n484), .Z(n486) );
  XNOR2_X1 U583 ( .A(n487), .B(n486), .ZN(n489) );
  XNOR2_X1 U584 ( .A(n489), .B(n488), .ZN(n663) );
  NOR2_X1 U585 ( .A1(G902), .A2(n663), .ZN(n490) );
  XOR2_X1 U586 ( .A(n491), .B(n490), .Z(n509) );
  INV_X1 U587 ( .A(n509), .ZN(n495) );
  NAND2_X1 U588 ( .A1(n508), .A2(n495), .ZN(n549) );
  XNOR2_X1 U589 ( .A(n549), .B(KEYINPUT75), .ZN(n492) );
  NAND2_X1 U590 ( .A1(n493), .A2(n492), .ZN(n494) );
  XNOR2_X1 U591 ( .A(n494), .B(KEYINPUT35), .ZN(n700) );
  XOR2_X1 U592 ( .A(KEYINPUT70), .B(KEYINPUT22), .Z(n497) );
  XOR2_X1 U593 ( .A(n523), .B(KEYINPUT84), .Z(n563) );
  XOR2_X1 U594 ( .A(KEYINPUT77), .B(n520), .Z(n499) );
  NOR2_X1 U595 ( .A1(n563), .A2(n499), .ZN(n500) );
  NOR2_X1 U596 ( .A1(n505), .A2(n638), .ZN(n503) );
  NOR2_X1 U597 ( .A1(n642), .A2(n528), .ZN(n502) );
  NAND2_X1 U598 ( .A1(n503), .A2(n502), .ZN(n602) );
  NAND2_X1 U599 ( .A1(n642), .A2(n504), .ZN(n647) );
  NOR2_X1 U600 ( .A1(n505), .A2(n647), .ZN(n507) );
  XNOR2_X1 U601 ( .A(KEYINPUT92), .B(KEYINPUT31), .ZN(n506) );
  XNOR2_X1 U602 ( .A(n507), .B(n506), .ZN(n617) );
  NAND2_X1 U603 ( .A1(n602), .A2(n617), .ZN(n511) );
  NOR2_X1 U604 ( .A1(n509), .A2(n508), .ZN(n611) );
  NAND2_X1 U605 ( .A1(n509), .A2(n508), .ZN(n616) );
  INV_X1 U606 ( .A(n616), .ZN(n607) );
  NOR2_X1 U607 ( .A1(n611), .A2(n607), .ZN(n510) );
  XOR2_X1 U608 ( .A(KEYINPUT99), .B(n510), .Z(n630) );
  INV_X1 U609 ( .A(n630), .ZN(n548) );
  NAND2_X1 U610 ( .A1(n511), .A2(n548), .ZN(n514) );
  NOR2_X1 U611 ( .A1(n520), .A2(n512), .ZN(n513) );
  NAND2_X1 U612 ( .A1(n635), .A2(n513), .ZN(n598) );
  NAND2_X1 U613 ( .A1(n514), .A2(n598), .ZN(n515) );
  INV_X1 U614 ( .A(n611), .ZN(n614) );
  INV_X1 U615 ( .A(n634), .ZN(n517) );
  NOR2_X1 U616 ( .A1(n517), .A2(n516), .ZN(n519) );
  NAND2_X1 U617 ( .A1(G953), .A2(G900), .ZN(n518) );
  NAND2_X1 U618 ( .A1(n519), .A2(n518), .ZN(n526) );
  NOR2_X1 U619 ( .A1(n635), .A2(n526), .ZN(n538) );
  XNOR2_X1 U620 ( .A(n521), .B(KEYINPUT102), .ZN(n522) );
  NOR2_X1 U621 ( .A1(n523), .A2(n559), .ZN(n524) );
  XNOR2_X1 U622 ( .A(n524), .B(KEYINPUT43), .ZN(n525) );
  NOR2_X1 U623 ( .A1(n534), .A2(n525), .ZN(n622) );
  INV_X1 U624 ( .A(n526), .ZN(n527) );
  XNOR2_X1 U625 ( .A(n529), .B(KEYINPUT73), .ZN(n532) );
  NAND2_X1 U626 ( .A1(n642), .A2(n624), .ZN(n530) );
  XOR2_X1 U627 ( .A(KEYINPUT30), .B(n530), .Z(n531) );
  NAND2_X1 U628 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U629 ( .A(n533), .B(KEYINPUT72), .ZN(n550) );
  XOR2_X1 U630 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n544) );
  AND2_X1 U631 ( .A1(n642), .A2(n538), .ZN(n539) );
  XNOR2_X1 U632 ( .A(KEYINPUT28), .B(n539), .ZN(n541) );
  XOR2_X1 U633 ( .A(n528), .B(KEYINPUT104), .Z(n540) );
  NAND2_X1 U634 ( .A1(n541), .A2(n540), .ZN(n547) );
  INV_X1 U635 ( .A(n542), .ZN(n628) );
  NOR2_X1 U636 ( .A1(n629), .A2(n628), .ZN(n543) );
  XOR2_X1 U637 ( .A(KEYINPUT46), .B(KEYINPUT81), .Z(n545) );
  NAND2_X1 U638 ( .A1(n612), .A2(n548), .ZN(n554) );
  OR2_X1 U639 ( .A1(KEYINPUT47), .A2(n554), .ZN(n558) );
  NOR2_X1 U640 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U641 ( .A1(n534), .A2(n551), .ZN(n553) );
  NAND2_X1 U642 ( .A1(n554), .A2(KEYINPUT47), .ZN(n555) );
  XNOR2_X1 U643 ( .A(n556), .B(KEYINPUT79), .ZN(n557) );
  AND2_X1 U644 ( .A1(n558), .A2(n557), .ZN(n564) );
  XOR2_X1 U645 ( .A(KEYINPUT36), .B(n561), .Z(n562) );
  NAND2_X1 U646 ( .A1(n607), .A2(n566), .ZN(n621) );
  NAND2_X1 U647 ( .A1(n567), .A2(KEYINPUT2), .ZN(n568) );
  XNOR2_X1 U648 ( .A(KEYINPUT66), .B(n568), .ZN(n569) );
  NAND2_X1 U649 ( .A1(n669), .A2(G210), .ZN(n577) );
  XNOR2_X1 U650 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n575) );
  XNOR2_X1 U651 ( .A(n573), .B(KEYINPUT118), .ZN(n574) );
  XNOR2_X1 U652 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U653 ( .A(n577), .B(n576), .ZN(n578) );
  INV_X1 U654 ( .A(KEYINPUT119), .ZN(n579) );
  XNOR2_X1 U655 ( .A(n579), .B(KEYINPUT56), .ZN(n580) );
  XNOR2_X1 U656 ( .A(n581), .B(n580), .ZN(G51) );
  XNOR2_X1 U657 ( .A(n582), .B(KEYINPUT62), .ZN(n584) );
  NAND2_X1 U658 ( .A1(n669), .A2(G472), .ZN(n583) );
  XNOR2_X1 U659 ( .A(n584), .B(n583), .ZN(n585) );
  NOR2_X2 U660 ( .A1(n585), .A2(n673), .ZN(n589) );
  XNOR2_X1 U661 ( .A(KEYINPUT83), .B(KEYINPUT85), .ZN(n587) );
  XNOR2_X1 U662 ( .A(n589), .B(n588), .ZN(G57) );
  XOR2_X1 U663 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n592) );
  XNOR2_X1 U664 ( .A(n590), .B(KEYINPUT120), .ZN(n591) );
  XNOR2_X1 U665 ( .A(n592), .B(n591), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n669), .A2(G469), .ZN(n593) );
  XNOR2_X1 U667 ( .A(n594), .B(n593), .ZN(n595) );
  NOR2_X2 U668 ( .A1(n595), .A2(n673), .ZN(n597) );
  INV_X1 U669 ( .A(KEYINPUT121), .ZN(n596) );
  XNOR2_X1 U670 ( .A(n597), .B(n596), .ZN(G54) );
  XNOR2_X1 U671 ( .A(G101), .B(n598), .ZN(G3) );
  NOR2_X1 U672 ( .A1(n614), .A2(n602), .ZN(n599) );
  XOR2_X1 U673 ( .A(G104), .B(n599), .Z(G6) );
  XOR2_X1 U674 ( .A(KEYINPUT108), .B(KEYINPUT26), .Z(n601) );
  XNOR2_X1 U675 ( .A(G107), .B(KEYINPUT27), .ZN(n600) );
  XNOR2_X1 U676 ( .A(n601), .B(n600), .ZN(n604) );
  NOR2_X1 U677 ( .A1(n616), .A2(n602), .ZN(n603) );
  XOR2_X1 U678 ( .A(n604), .B(n603), .Z(G9) );
  XNOR2_X1 U679 ( .A(G110), .B(n605), .ZN(n606) );
  XNOR2_X1 U680 ( .A(n606), .B(KEYINPUT109), .ZN(G12) );
  XOR2_X1 U681 ( .A(KEYINPUT110), .B(KEYINPUT29), .Z(n609) );
  NAND2_X1 U682 ( .A1(n612), .A2(n607), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n609), .B(n608), .ZN(n610) );
  XNOR2_X1 U684 ( .A(G128), .B(n610), .ZN(G30) );
  NAND2_X1 U685 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U686 ( .A(n613), .B(G146), .ZN(G48) );
  NOR2_X1 U687 ( .A1(n617), .A2(n614), .ZN(n615) );
  XOR2_X1 U688 ( .A(G113), .B(n615), .Z(G15) );
  NOR2_X1 U689 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U690 ( .A(G116), .B(n618), .Z(G18) );
  XNOR2_X1 U691 ( .A(G125), .B(n619), .ZN(n620) );
  XNOR2_X1 U692 ( .A(n620), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U693 ( .A(G134), .B(n621), .ZN(G36) );
  XOR2_X1 U694 ( .A(G140), .B(n622), .Z(G42) );
  NAND2_X1 U695 ( .A1(G952), .A2(n623), .ZN(n655) );
  NOR2_X1 U696 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U697 ( .A(KEYINPUT113), .B(n626), .Z(n627) );
  NOR2_X1 U698 ( .A1(n628), .A2(n627), .ZN(n632) );
  NOR2_X1 U699 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U700 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U701 ( .A1(n657), .A2(n633), .ZN(n651) );
  OR2_X1 U702 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U703 ( .A(n636), .B(KEYINPUT49), .ZN(n637) );
  XNOR2_X1 U704 ( .A(KEYINPUT111), .B(n637), .ZN(n645) );
  XOR2_X1 U705 ( .A(KEYINPUT50), .B(KEYINPUT112), .Z(n641) );
  NAND2_X1 U706 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U707 ( .A(n641), .B(n640), .ZN(n643) );
  NOR2_X1 U708 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U709 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U710 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U711 ( .A(KEYINPUT51), .B(n648), .ZN(n649) );
  NOR2_X1 U712 ( .A1(n658), .A2(n649), .ZN(n650) );
  NOR2_X1 U713 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U714 ( .A(KEYINPUT114), .B(n652), .ZN(n653) );
  XNOR2_X1 U715 ( .A(KEYINPUT52), .B(n653), .ZN(n654) );
  NOR2_X1 U716 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U717 ( .A(KEYINPUT115), .B(n656), .Z(n660) );
  NOR2_X1 U718 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U719 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U720 ( .A(KEYINPUT116), .B(n661), .Z(n662) );
  NAND2_X1 U721 ( .A1(n669), .A2(G475), .ZN(n664) );
  XNOR2_X1 U722 ( .A(n665), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U723 ( .A1(G478), .A2(n669), .ZN(n666) );
  XNOR2_X1 U724 ( .A(n667), .B(n666), .ZN(n668) );
  NOR2_X1 U725 ( .A1(n673), .A2(n668), .ZN(G63) );
  XOR2_X1 U726 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n670) );
  NOR2_X1 U727 ( .A1(n673), .A2(n672), .ZN(G66) );
  NAND2_X1 U728 ( .A1(G224), .A2(G953), .ZN(n674) );
  XNOR2_X1 U729 ( .A(n674), .B(KEYINPUT61), .ZN(n675) );
  XNOR2_X1 U730 ( .A(KEYINPUT124), .B(n675), .ZN(n676) );
  NAND2_X1 U731 ( .A1(n676), .A2(G898), .ZN(n677) );
  XNOR2_X1 U732 ( .A(n677), .B(KEYINPUT125), .ZN(n680) );
  NOR2_X1 U733 ( .A1(n678), .A2(G953), .ZN(n679) );
  NOR2_X1 U734 ( .A1(n680), .A2(n679), .ZN(n685) );
  NOR2_X1 U735 ( .A1(G898), .A2(n691), .ZN(n683) );
  XOR2_X1 U736 ( .A(n681), .B(G101), .Z(n682) );
  NOR2_X1 U737 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U738 ( .A(n685), .B(n684), .Z(G69) );
  XOR2_X1 U739 ( .A(n687), .B(n686), .Z(n688) );
  XNOR2_X1 U740 ( .A(n689), .B(n688), .ZN(n693) );
  XNOR2_X1 U741 ( .A(n693), .B(n690), .ZN(n692) );
  NAND2_X1 U742 ( .A1(n692), .A2(n691), .ZN(n697) );
  XNOR2_X1 U743 ( .A(G227), .B(n693), .ZN(n694) );
  NAND2_X1 U744 ( .A1(n694), .A2(G900), .ZN(n695) );
  NAND2_X1 U745 ( .A1(G953), .A2(n695), .ZN(n696) );
  NAND2_X1 U746 ( .A1(n697), .A2(n696), .ZN(G72) );
  XNOR2_X1 U747 ( .A(G137), .B(n698), .ZN(n699) );
  XNOR2_X1 U748 ( .A(n699), .B(KEYINPUT126), .ZN(G39) );
  XOR2_X1 U749 ( .A(n700), .B(G122), .Z(G24) );
  XNOR2_X1 U750 ( .A(G143), .B(n701), .ZN(G45) );
  XNOR2_X1 U751 ( .A(n702), .B(G131), .ZN(G33) );
endmodule

