//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n797, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  INV_X1    g004(.A(G8gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G64gat), .ZN(new_n208));
  AND2_X1   g007(.A1(new_n208), .A2(G57gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(G57gat), .ZN(new_n210));
  AND2_X1   g009(.A1(G71gat), .A2(G78gat), .ZN(new_n211));
  OAI22_X1  g010(.A1(new_n209), .A2(new_n210), .B1(KEYINPUT9), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G71gat), .B(G78gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT21), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n207), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(new_n217), .B(G183gat), .Z(new_n218));
  AND2_X1   g017(.A1(G231gat), .A2(G233gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT88), .B(KEYINPUT89), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n214), .A2(KEYINPUT21), .ZN(new_n223));
  XNOR2_X1  g022(.A(G127gat), .B(G155gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(G211gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n223), .B(new_n225), .ZN(new_n226));
  XOR2_X1   g025(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n222), .B(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(G29gat), .A2(G36gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT14), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G43gat), .B(G50gat), .ZN(new_n233));
  INV_X1    g032(.A(G29gat), .ZN(new_n234));
  XOR2_X1   g033(.A(KEYINPUT86), .B(G36gat), .Z(new_n235));
  OAI221_X1 g034(.A(new_n232), .B1(KEYINPUT15), .B2(new_n233), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(KEYINPUT15), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n236), .B(new_n237), .Z(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(KEYINPUT17), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT7), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT91), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT92), .ZN(new_n242));
  OAI211_X1 g041(.A(G85gat), .B(G92gat), .C1(new_n240), .C2(KEYINPUT91), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT92), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n241), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(new_n243), .ZN(new_n248));
  NAND2_X1  g047(.A1(G99gat), .A2(G106gat), .ZN(new_n249));
  INV_X1    g048(.A(G85gat), .ZN(new_n250));
  INV_X1    g049(.A(G92gat), .ZN(new_n251));
  AOI22_X1  g050(.A1(KEYINPUT8), .A2(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n245), .A2(new_n248), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G99gat), .B(G106gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT93), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n255), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n257), .A2(new_n245), .A3(new_n248), .A4(new_n252), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n239), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT90), .B(KEYINPUT95), .Z(new_n261));
  NAND3_X1  g060(.A1(new_n238), .A2(new_n258), .A3(new_n256), .ZN(new_n262));
  NAND3_X1  g061(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OR3_X1    g063(.A1(new_n260), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n261), .B1(new_n260), .B2(new_n264), .ZN(new_n266));
  XNOR2_X1  g065(.A(G134gat), .B(G162gat), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G190gat), .B(G218gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT94), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n269), .B(new_n271), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n265), .A2(new_n266), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n272), .B1(new_n265), .B2(new_n266), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n229), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G230gat), .ZN(new_n278));
  INV_X1    g077(.A(G233gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT96), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n259), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n256), .A2(new_n258), .A3(KEYINPUT96), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n215), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n259), .A2(new_n282), .A3(new_n214), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT10), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n256), .A2(new_n258), .A3(KEYINPUT10), .A4(new_n214), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n281), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n285), .A2(new_n286), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n280), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G120gat), .B(G148gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(G204gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(KEYINPUT97), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n296), .B(G176gat), .Z(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT98), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n297), .B1(new_n290), .B2(new_n292), .ZN(new_n301));
  OR3_X1    g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n293), .A2(new_n300), .A3(new_n298), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n277), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT99), .ZN(new_n306));
  INV_X1    g105(.A(new_n304), .ZN(new_n307));
  NOR3_X1   g106(.A1(new_n229), .A2(new_n307), .A3(new_n276), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT99), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n239), .A2(new_n207), .ZN(new_n312));
  NAND2_X1  g111(.A1(G229gat), .A2(G233gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n207), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n238), .A2(new_n314), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n312), .A2(KEYINPUT18), .A3(new_n313), .A4(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n238), .B(new_n314), .ZN(new_n317));
  XOR2_X1   g116(.A(new_n313), .B(KEYINPUT13), .Z(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT87), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT11), .B(G169gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(G197gat), .ZN(new_n324));
  XOR2_X1   g123(.A(G113gat), .B(G141gat), .Z(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(KEYINPUT12), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n312), .A2(new_n315), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT18), .B1(new_n329), .B2(new_n313), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n322), .B(new_n328), .C1(new_n330), .C2(new_n320), .ZN(new_n331));
  INV_X1    g130(.A(new_n330), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n332), .B(new_n321), .C1(KEYINPUT87), .C2(new_n327), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT37), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT74), .B(G204gat), .ZN(new_n337));
  INV_X1    g136(.A(G197gat), .ZN(new_n338));
  OR2_X1    g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n338), .ZN(new_n340));
  INV_X1    g139(.A(G211gat), .ZN(new_n341));
  INV_X1    g140(.A(G218gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n339), .B(new_n340), .C1(KEYINPUT22), .C2(new_n343), .ZN(new_n344));
  XOR2_X1   g143(.A(G211gat), .B(G218gat), .Z(new_n345));
  XOR2_X1   g144(.A(new_n344), .B(new_n345), .Z(new_n346));
  NAND2_X1  g145(.A1(G226gat), .A2(G233gat), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT25), .ZN(new_n349));
  NAND2_X1  g148(.A1(G183gat), .A2(G190gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT66), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT66), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n352), .A2(G183gat), .A3(G190gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT65), .ZN(new_n355));
  OAI22_X1  g154(.A1(new_n355), .A2(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n349), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT23), .ZN(new_n359));
  NAND2_X1  g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n361), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n356), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(new_n351), .A3(new_n353), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n357), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT24), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n350), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(G183gat), .A2(G190gat), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n349), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n366), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT28), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(KEYINPUT67), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G190gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT67), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n382), .B1(new_n383), .B2(KEYINPUT28), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n381), .A2(KEYINPUT68), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT68), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT27), .B(G183gat), .ZN(new_n387));
  AOI21_X1  g186(.A(G190gat), .B1(new_n376), .B2(KEYINPUT67), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n378), .B1(new_n385), .B2(new_n389), .ZN(new_n390));
  OR2_X1    g189(.A1(G169gat), .A2(G176gat), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT26), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n350), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n391), .A2(new_n392), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n393), .B1(new_n360), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT68), .B1(new_n381), .B2(new_n384), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n387), .A2(new_n386), .A3(new_n388), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n377), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n390), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n375), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT29), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n348), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT69), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n390), .A2(KEYINPUT69), .A3(new_n395), .A4(new_n398), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n375), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(KEYINPUT75), .A3(new_n348), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT75), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n374), .B1(new_n404), .B2(new_n405), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n409), .B1(new_n410), .B2(new_n347), .ZN(new_n411));
  AOI211_X1 g210(.A(new_n346), .B(new_n402), .C1(new_n408), .C2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n375), .A2(new_n348), .A3(new_n399), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n347), .A2(new_n401), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n413), .B(new_n346), .C1(new_n410), .C2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n336), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n344), .B(new_n345), .ZN(new_n418));
  INV_X1    g217(.A(new_n402), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT75), .B1(new_n407), .B2(new_n348), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n410), .A2(new_n409), .A3(new_n347), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n418), .B(new_n419), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n422), .A2(KEYINPUT76), .A3(new_n415), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n335), .B1(new_n417), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n335), .A3(new_n415), .ZN(new_n425));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(new_n208), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(new_n251), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT38), .B1(new_n424), .B2(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n346), .B(new_n419), .C1(new_n420), .C2(new_n421), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n418), .B(new_n413), .C1(new_n410), .C2(new_n414), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(KEYINPUT37), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT38), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n425), .A2(new_n433), .A3(new_n434), .A4(new_n428), .ZN(new_n435));
  NAND2_X1  g234(.A1(G225gat), .A2(G233gat), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G120gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(G113gat), .ZN(new_n439));
  INV_X1    g238(.A(G113gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(G120gat), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(G127gat), .B1(new_n442), .B2(KEYINPUT1), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT1), .B1(new_n439), .B2(new_n441), .ZN(new_n444));
  INV_X1    g243(.A(G127gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n443), .A2(G134gat), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G134gat), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n444), .A2(new_n445), .ZN(new_n449));
  AOI211_X1 g248(.A(KEYINPUT1), .B(G127gat), .C1(new_n439), .C2(new_n441), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(G148gat), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n452), .A2(G141gat), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT78), .B(G148gat), .ZN(new_n455));
  INV_X1    g254(.A(G141gat), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(G155gat), .A2(G162gat), .ZN(new_n458));
  NOR2_X1   g257(.A1(G155gat), .A2(G162gat), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n458), .B1(new_n460), .B2(KEYINPUT2), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT2), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n456), .A2(G148gat), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n462), .B1(new_n453), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n458), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n465), .A2(new_n459), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n457), .A2(new_n461), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n447), .A2(new_n451), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n467), .B1(new_n447), .B2(new_n451), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n437), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT80), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT79), .B(KEYINPUT4), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n447), .A2(new_n451), .ZN(new_n475));
  INV_X1    g274(.A(new_n467), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n467), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n465), .B1(new_n462), .B2(new_n459), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n452), .A2(KEYINPUT78), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n452), .A2(KEYINPUT78), .ZN(new_n482));
  OAI21_X1  g281(.A(G141gat), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n480), .B1(new_n483), .B2(new_n454), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n464), .A2(new_n466), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT3), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n475), .A2(new_n479), .A3(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n447), .A2(new_n451), .A3(KEYINPUT4), .A4(new_n467), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n477), .A2(new_n487), .A3(new_n436), .A4(new_n488), .ZN(new_n489));
  OAI211_X1 g288(.A(KEYINPUT80), .B(new_n437), .C1(new_n468), .C2(new_n469), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n472), .A2(KEYINPUT5), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n468), .A2(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n468), .A2(new_n473), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n437), .A2(KEYINPUT5), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n492), .A2(new_n487), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(G1gat), .B(G29gat), .Z(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G57gat), .B(G85gat), .ZN(new_n500));
  XOR2_X1   g299(.A(new_n499), .B(new_n500), .Z(new_n501));
  NAND3_X1  g300(.A1(new_n496), .A2(KEYINPUT6), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT84), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n496), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(new_n501), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n496), .A2(new_n501), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT6), .ZN(new_n508));
  INV_X1    g307(.A(new_n501), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n491), .A2(new_n509), .A3(new_n495), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n435), .A2(new_n506), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n428), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n422), .A2(new_n415), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n430), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(G228gat), .A2(G233gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(G22gat), .ZN(new_n517));
  XOR2_X1   g316(.A(G78gat), .B(G106gat), .Z(new_n518));
  XOR2_X1   g317(.A(new_n517), .B(new_n518), .Z(new_n519));
  NAND2_X1  g318(.A1(new_n479), .A2(new_n401), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n346), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT3), .B1(new_n418), .B2(new_n401), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n521), .B1(new_n522), .B2(new_n467), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n523), .A2(KEYINPUT82), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(KEYINPUT82), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n519), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n523), .A2(KEYINPUT82), .ZN(new_n527));
  INV_X1    g326(.A(new_n519), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n523), .A2(KEYINPUT82), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT83), .B(G50gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT31), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n526), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n532), .B1(new_n526), .B2(new_n530), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT30), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n514), .B(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n423), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT76), .B1(new_n422), .B2(new_n415), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n428), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT77), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n513), .B1(new_n417), .B2(new_n423), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT77), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n538), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n492), .A2(new_n487), .A3(new_n493), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n437), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n548), .A2(KEYINPUT39), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n468), .A2(new_n469), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n548), .B(KEYINPUT39), .C1(new_n437), .C2(new_n550), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n549), .A2(new_n551), .A3(new_n509), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n552), .A2(KEYINPUT40), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(KEYINPUT40), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n507), .A3(new_n554), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n515), .B(new_n536), .C1(new_n546), .C2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT36), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n475), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n560), .B1(new_n406), .B2(new_n375), .ZN(new_n561));
  AOI211_X1 g360(.A(new_n475), .B(new_n374), .C1(new_n404), .C2(new_n405), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(G227gat), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n564), .A2(new_n279), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n559), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NOR4_X1   g366(.A1(new_n561), .A2(new_n562), .A3(new_n565), .A4(new_n558), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n565), .B1(new_n561), .B2(new_n562), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT32), .ZN(new_n571));
  XOR2_X1   g370(.A(KEYINPUT70), .B(KEYINPUT33), .Z(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G15gat), .B(G43gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(G71gat), .ZN(new_n576));
  INV_X1    g375(.A(G99gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n571), .A2(new_n574), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n578), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n570), .B(KEYINPUT32), .C1(new_n573), .C2(new_n580), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n569), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n568), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n563), .A2(new_n566), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(new_n558), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n579), .A2(new_n581), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n557), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT73), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT73), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n589), .B(new_n557), .C1(new_n582), .C2(new_n586), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n579), .A2(new_n581), .ZN(new_n592));
  INV_X1    g391(.A(new_n569), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n569), .A2(new_n579), .A3(new_n581), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(KEYINPUT36), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT72), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT72), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n594), .A2(new_n598), .A3(KEYINPUT36), .A4(new_n595), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n591), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n511), .A2(new_n502), .ZN(new_n602));
  INV_X1    g401(.A(new_n538), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n543), .A2(new_n544), .ZN(new_n604));
  AOI211_X1 g403(.A(KEYINPUT77), .B(new_n513), .C1(new_n417), .C2(new_n423), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n602), .B(new_n603), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n535), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n556), .A2(new_n601), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n582), .A2(new_n586), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n536), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT35), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n535), .A2(new_n582), .A3(new_n586), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT35), .B1(new_n506), .B2(new_n511), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(new_n546), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT85), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n608), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n608), .A2(new_n615), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT85), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n311), .A2(new_n334), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n617), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n616), .B1(new_n608), .B2(new_n615), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n625), .A2(KEYINPUT100), .A3(new_n334), .A4(new_n311), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n602), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G1gat), .ZN(G1324gat));
  INV_X1    g429(.A(new_n546), .ZN(new_n631));
  NAND2_X1  g430(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n203), .A2(new_n206), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n627), .A2(new_n631), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n634), .A2(KEYINPUT42), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(KEYINPUT42), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n627), .A2(new_n631), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n637), .A2(KEYINPUT101), .A3(G8gat), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT101), .B1(new_n637), .B2(G8gat), .ZN(new_n639));
  OAI22_X1  g438(.A1(new_n635), .A2(new_n636), .B1(new_n638), .B2(new_n639), .ZN(G1325gat));
  AOI21_X1  g439(.A(G15gat), .B1(new_n627), .B2(new_n609), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n641), .A2(KEYINPUT102), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(KEYINPUT102), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n601), .B(KEYINPUT103), .Z(new_n644));
  AOI21_X1  g443(.A(new_n644), .B1(new_n622), .B2(new_n626), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n642), .A2(new_n643), .B1(new_n645), .B2(G15gat), .ZN(G1326gat));
  NAND2_X1  g445(.A1(new_n627), .A2(new_n535), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT43), .B(G22gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(G1327gat));
  NAND3_X1  g448(.A1(new_n619), .A2(new_n617), .A3(new_n276), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n229), .ZN(new_n652));
  INV_X1    g451(.A(new_n334), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n652), .A2(new_n653), .A3(new_n307), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n655), .A2(G29gat), .A3(new_n602), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n650), .A2(KEYINPUT44), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n608), .A2(KEYINPUT105), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT105), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n556), .A2(new_n601), .A3(new_n661), .A4(new_n607), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n660), .A2(new_n615), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(new_n664), .A3(new_n276), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n654), .ZN(new_n667));
  OAI21_X1  g466(.A(G29gat), .B1(new_n667), .B2(new_n602), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n658), .A2(new_n668), .ZN(G1328gat));
  NAND4_X1  g468(.A1(new_n651), .A2(new_n235), .A3(new_n631), .A4(new_n654), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n670), .B(KEYINPUT46), .Z(new_n671));
  NOR2_X1   g470(.A1(new_n667), .A2(new_n546), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n671), .B1(new_n235), .B2(new_n672), .ZN(G1329gat));
  INV_X1    g472(.A(G43gat), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n651), .A2(new_n674), .A3(new_n609), .A4(new_n654), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT106), .ZN(new_n676));
  OAI21_X1  g475(.A(G43gat), .B1(new_n667), .B2(new_n601), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(KEYINPUT47), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(G43gat), .B1(new_n667), .B2(new_n644), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n678), .B1(new_n680), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g480(.A(G50gat), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n655), .B2(new_n536), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT48), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n535), .A2(G50gat), .ZN(new_n685));
  OAI221_X1 g484(.A(new_n683), .B1(KEYINPUT107), .B2(new_n684), .C1(new_n667), .C2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(KEYINPUT107), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1331gat));
  NAND3_X1  g487(.A1(new_n277), .A2(new_n653), .A3(new_n307), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT108), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n663), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n628), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g493(.A(new_n546), .B(new_n691), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n695));
  NOR2_X1   g494(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1333gat));
  INV_X1    g496(.A(G71gat), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n692), .A2(new_n698), .A3(new_n609), .ZN(new_n699));
  OAI21_X1  g498(.A(G71gat), .B1(new_n691), .B2(new_n644), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g501(.A1(new_n691), .A2(new_n536), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT109), .B(G78gat), .Z(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1335gat));
  NOR2_X1   g504(.A1(new_n652), .A2(new_n334), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n307), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n666), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(G85gat), .B1(new_n709), .B2(new_n602), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n663), .A2(new_n276), .A3(new_n706), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT51), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n304), .A2(G85gat), .A3(new_n602), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT110), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n710), .A2(new_n716), .ZN(G1336gat));
  OAI21_X1  g516(.A(G92gat), .B1(new_n709), .B2(new_n546), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n713), .A2(new_n251), .A3(new_n631), .A4(new_n307), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(KEYINPUT111), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n721), .A3(KEYINPUT52), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT52), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n718), .B(new_n719), .C1(KEYINPUT111), .C2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(G1337gat));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n644), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n713), .A2(new_n307), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n609), .A2(new_n577), .ZN(new_n728));
  OAI22_X1  g527(.A1(new_n726), .A2(new_n577), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT112), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n731));
  OAI221_X1 g530(.A(new_n731), .B1(new_n727), .B2(new_n728), .C1(new_n726), .C2(new_n577), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(G1338gat));
  INV_X1    g532(.A(KEYINPUT114), .ZN(new_n734));
  AOI211_X1 g533(.A(new_n536), .B(new_n707), .C1(new_n659), .C2(new_n665), .ZN(new_n735));
  XOR2_X1   g534(.A(KEYINPUT113), .B(G106gat), .Z(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n734), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n666), .A2(new_n535), .A3(new_n708), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n739), .A2(KEYINPUT114), .A3(new_n736), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n536), .A2(G106gat), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n307), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT115), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n713), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n738), .A2(new_n740), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(KEYINPUT53), .ZN(new_n746));
  AND4_X1   g545(.A1(KEYINPUT116), .A2(new_n666), .A3(new_n535), .A4(new_n708), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n707), .B1(new_n659), .B2(new_n665), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT116), .B1(new_n748), .B2(new_n535), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n736), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n713), .A2(new_n307), .A3(new_n741), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n746), .A2(new_n753), .ZN(G1339gat));
  OAI211_X1 g553(.A(new_n280), .B(new_n288), .C1(new_n291), .C2(KEYINPUT10), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n755), .A2(KEYINPUT54), .A3(new_n290), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT54), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n757), .B(new_n281), .C1(new_n287), .C2(new_n289), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n758), .A2(KEYINPUT117), .A3(new_n298), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT117), .B1(new_n758), .B2(new_n298), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n756), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n299), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI211_X1 g562(.A(KEYINPUT55), .B(new_n756), .C1(new_n759), .C2(new_n760), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT118), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n758), .A2(new_n298), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n758), .A2(KEYINPUT117), .A3(new_n298), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n771), .A2(KEYINPUT118), .A3(KEYINPUT55), .A4(new_n756), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n763), .A2(new_n766), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT119), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n763), .A2(new_n766), .A3(new_n772), .A4(KEYINPUT119), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(new_n334), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n332), .A2(new_n321), .A3(new_n327), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n329), .A2(new_n313), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n317), .A2(new_n318), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n326), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n304), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n276), .B1(new_n777), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n782), .A2(new_n275), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n775), .A2(new_n776), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n229), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n305), .A2(new_n334), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n610), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n631), .A2(new_n602), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n793), .A2(new_n653), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(new_n440), .ZN(G1340gat));
  NOR2_X1   g594(.A1(new_n793), .A2(new_n304), .ZN(new_n796));
  XNOR2_X1  g595(.A(KEYINPUT120), .B(G120gat), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n796), .B(new_n797), .ZN(G1341gat));
  NOR2_X1   g597(.A1(new_n793), .A2(new_n229), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(new_n445), .ZN(G1342gat));
  NAND4_X1  g599(.A1(new_n791), .A2(new_n448), .A3(new_n276), .A4(new_n792), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT56), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n790), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n805), .A2(new_n612), .A3(new_n276), .A4(new_n792), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT121), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n806), .A2(new_n807), .A3(G134gat), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n807), .B1(new_n806), .B2(G134gat), .ZN(new_n809));
  OAI22_X1  g608(.A1(new_n803), .A2(new_n804), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT122), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI221_X1 g611(.A(KEYINPUT122), .B1(new_n808), .B2(new_n809), .C1(new_n803), .C2(new_n804), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(G1343gat));
  AOI21_X1  g613(.A(new_n536), .B1(new_n788), .B2(new_n790), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n792), .A2(new_n601), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n334), .A2(new_n763), .A3(new_n766), .A4(new_n772), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n783), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n275), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n652), .B1(new_n821), .B2(new_n786), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n535), .B1(new_n822), .B2(new_n789), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n818), .B1(new_n823), .B2(KEYINPUT57), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n817), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(G141gat), .B1(new_n825), .B2(new_n653), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n815), .A2(new_n644), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n827), .A2(new_n456), .A3(new_n334), .A4(new_n792), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT58), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT58), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n826), .A2(new_n831), .A3(new_n828), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(G1344gat));
  AND2_X1   g632(.A1(new_n827), .A2(new_n792), .ZN(new_n834));
  INV_X1    g633(.A(new_n455), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n835), .A3(new_n307), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n817), .A2(new_n307), .A3(new_n824), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT123), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n835), .A2(KEYINPUT59), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n838), .B1(new_n837), .B2(new_n839), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n815), .A2(new_n816), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n276), .B1(new_n819), .B2(new_n783), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n773), .A2(new_n275), .A3(new_n782), .ZN(new_n846));
  OR3_X1    g645(.A1(new_n845), .A2(new_n846), .A3(KEYINPUT124), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT124), .B1(new_n845), .B2(new_n846), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n847), .A2(new_n229), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n311), .A2(new_n653), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n816), .A3(new_n535), .ZN(new_n852));
  INV_X1    g651(.A(new_n818), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n844), .A2(new_n852), .A3(new_n307), .A4(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n843), .B1(new_n854), .B2(G148gat), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n836), .B1(new_n842), .B2(new_n855), .ZN(G1345gat));
  INV_X1    g655(.A(G155gat), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n825), .A2(new_n857), .A3(new_n229), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n834), .A2(new_n652), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n858), .B1(new_n859), .B2(new_n857), .ZN(G1346gat));
  INV_X1    g659(.A(G162gat), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n825), .A2(new_n861), .A3(new_n275), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n834), .A2(new_n276), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(new_n861), .ZN(G1347gat));
  NOR2_X1   g663(.A1(new_n546), .A2(new_n628), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n791), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n334), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n307), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g669(.A1(new_n866), .A2(new_n652), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(G183gat), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n872), .B1(new_n381), .B2(new_n871), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT60), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT60), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n872), .B(new_n875), .C1(new_n381), .C2(new_n871), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(G1350gat));
  NAND2_X1  g676(.A1(new_n866), .A2(new_n276), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT61), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n878), .A2(new_n879), .A3(new_n382), .ZN(new_n880));
  XOR2_X1   g679(.A(KEYINPUT61), .B(G190gat), .Z(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n878), .B2(new_n881), .ZN(G1351gat));
  AND2_X1   g681(.A1(new_n644), .A2(new_n865), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n844), .A2(new_n852), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(G197gat), .B1(new_n884), .B2(new_n653), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n827), .A2(new_n865), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT125), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n827), .A2(new_n888), .A3(new_n865), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n887), .A2(new_n338), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n885), .B1(new_n890), .B2(new_n653), .ZN(G1352gat));
  NAND3_X1  g690(.A1(new_n827), .A2(new_n307), .A3(new_n865), .ZN(new_n892));
  OR3_X1    g691(.A1(new_n892), .A2(KEYINPUT62), .A3(G204gat), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n844), .A2(new_n307), .A3(new_n852), .ZN(new_n894));
  INV_X1    g693(.A(new_n883), .ZN(new_n895));
  OAI21_X1  g694(.A(G204gat), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT62), .B1(new_n892), .B2(G204gat), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n893), .A2(new_n896), .A3(new_n897), .ZN(G1353gat));
  NAND4_X1  g697(.A1(new_n887), .A2(new_n341), .A3(new_n652), .A4(new_n889), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n844), .A2(new_n852), .A3(new_n652), .A4(new_n883), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT63), .B1(new_n900), .B2(G211gat), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(G1354gat));
  NAND3_X1  g703(.A1(new_n887), .A2(new_n276), .A3(new_n889), .ZN(new_n905));
  INV_X1    g704(.A(new_n884), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n276), .A2(G218gat), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT126), .ZN(new_n908));
  AOI22_X1  g707(.A1(new_n905), .A2(new_n342), .B1(new_n906), .B2(new_n908), .ZN(G1355gat));
endmodule


