//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n834, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G8gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(G43gat), .B(G50gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(KEYINPUT93), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n208), .B(KEYINPUT15), .ZN(new_n209));
  NOR3_X1   g008(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT94), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n212), .A2(new_n213), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n209), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G29gat), .A2(G36gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n213), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n216), .B1(new_n217), .B2(new_n210), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(KEYINPUT15), .A3(new_n207), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT17), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n206), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT95), .B1(new_n220), .B2(new_n221), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NOR3_X1   g023(.A1(new_n220), .A2(KEYINPUT95), .A3(new_n221), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n222), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G229gat), .A2(G233gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n220), .A2(new_n206), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n226), .A2(KEYINPUT18), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G113gat), .B(G141gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n230), .B(G197gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT11), .B(G169gat), .ZN(new_n232));
  XOR2_X1   g031(.A(new_n231), .B(new_n232), .Z(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT92), .B(KEYINPUT12), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n233), .B(new_n234), .Z(new_n235));
  XNOR2_X1  g034(.A(new_n220), .B(new_n206), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n227), .B(KEYINPUT13), .Z(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n229), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT97), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT96), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n240), .A2(KEYINPUT96), .A3(new_n241), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n245), .A2(new_n246), .A3(new_n238), .A4(new_n229), .ZN(new_n247));
  INV_X1    g046(.A(new_n235), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n239), .A2(new_n243), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT81), .ZN(new_n250));
  OR2_X1    g049(.A1(KEYINPUT79), .A2(G141gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(KEYINPUT79), .A2(G141gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(G148gat), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G148gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(G141gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(G155gat), .A2(G162gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(G155gat), .A2(G162gat), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT2), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n253), .A2(new_n255), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G155gat), .B(G162gat), .ZN(new_n261));
  INV_X1    g060(.A(G141gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G148gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n255), .A2(new_n263), .ZN(new_n264));
  AND2_X1   g063(.A1(KEYINPUT78), .A2(KEYINPUT2), .ZN(new_n265));
  NOR2_X1   g064(.A1(KEYINPUT78), .A2(KEYINPUT2), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n261), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n250), .B1(new_n260), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n256), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n270), .A2(new_n257), .ZN(new_n271));
  XNOR2_X1  g070(.A(G141gat), .B(G148gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT78), .B(KEYINPUT2), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n255), .ZN(new_n275));
  AND2_X1   g074(.A1(KEYINPUT79), .A2(G141gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(KEYINPUT79), .A2(G141gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n275), .B1(new_n278), .B2(G148gat), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n270), .B1(new_n258), .B2(new_n257), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n274), .B(KEYINPUT81), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n269), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT67), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G134gat), .ZN(new_n285));
  INV_X1    g084(.A(G120gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G113gat), .ZN(new_n287));
  INV_X1    g086(.A(G113gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G120gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT1), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n285), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI211_X1 g091(.A(KEYINPUT1), .B(G134gat), .C1(new_n287), .C2(new_n289), .ZN(new_n293));
  OAI21_X1  g092(.A(G127gat), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G113gat), .B(G120gat), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n284), .B(G134gat), .C1(new_n295), .C2(KEYINPUT1), .ZN(new_n296));
  INV_X1    g095(.A(G134gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n290), .A2(new_n291), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G127gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n296), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n282), .A2(new_n283), .A3(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n274), .B1(new_n279), .B2(new_n280), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n292), .A2(new_n293), .A3(G127gat), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n299), .B1(new_n296), .B2(new_n298), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT4), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT5), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT3), .B1(new_n260), .B2(new_n268), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT80), .B(KEYINPUT3), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n274), .B(new_n312), .C1(new_n279), .C2(new_n280), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n311), .A2(new_n313), .A3(new_n294), .A4(new_n300), .ZN(new_n314));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n309), .A2(new_n310), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT84), .ZN(new_n318));
  INV_X1    g117(.A(new_n315), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n294), .A2(new_n303), .A3(new_n300), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n303), .B1(new_n294), .B2(new_n300), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT83), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n294), .A2(new_n303), .A3(new_n300), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT83), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n326), .A3(new_n319), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT82), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n305), .A2(new_n306), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n269), .A2(new_n281), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n329), .B(KEYINPUT4), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n283), .B1(new_n282), .B2(new_n301), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n301), .A2(new_n283), .A3(new_n304), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT82), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n332), .B(new_n316), .C1(new_n333), .C2(new_n335), .ZN(new_n336));
  AND4_X1   g135(.A1(new_n318), .A2(new_n328), .A3(new_n336), .A4(KEYINPUT5), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n310), .B1(new_n323), .B2(new_n327), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n318), .B1(new_n338), .B2(new_n336), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n317), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G1gat), .B(G29gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(G57gat), .B(G85gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT85), .B(KEYINPUT0), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT6), .ZN(new_n346));
  OR2_X1    g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n346), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n340), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n336), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n326), .B1(new_n325), .B2(new_n319), .ZN(new_n351));
  AOI211_X1 g150(.A(KEYINPUT83), .B(new_n315), .C1(new_n307), .C2(new_n324), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT5), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT84), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n318), .A3(new_n336), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n356), .A2(new_n346), .A3(new_n317), .A4(new_n345), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n349), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G226gat), .A2(G233gat), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n359), .B(KEYINPUT74), .Z(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G183gat), .A2(G190gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(G169gat), .A2(G176gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT26), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NOR3_X1   g165(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n362), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(G183gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT27), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT27), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G183gat), .ZN(new_n372));
  INV_X1    g171(.A(G190gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT28), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT27), .B(G183gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n377), .A2(KEYINPUT28), .A3(new_n373), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n368), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n362), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT64), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n382), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT64), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT65), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n364), .B2(KEYINPUT23), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT23), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n389), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(G169gat), .ZN(new_n392));
  INV_X1    g191(.A(G176gat), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT23), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n394), .A2(new_n363), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n386), .A2(new_n391), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT25), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n384), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT66), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n363), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n397), .B1(new_n364), .B2(KEYINPUT23), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n391), .A2(new_n399), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n379), .B1(new_n398), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n361), .B1(new_n406), .B2(KEYINPUT29), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT75), .B1(new_n406), .B2(new_n359), .ZN(new_n408));
  INV_X1    g207(.A(new_n368), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n376), .A2(new_n378), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n363), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n412), .B1(new_n388), .B2(new_n390), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT25), .B1(new_n413), .B2(new_n386), .ZN(new_n414));
  INV_X1    g213(.A(new_n405), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n411), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT75), .ZN(new_n417));
  INV_X1    g216(.A(new_n359), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n407), .A2(new_n408), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n421));
  OR2_X1    g220(.A1(G197gat), .A2(G204gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(G197gat), .A2(G204gat), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n424), .A2(KEYINPUT73), .ZN(new_n425));
  XOR2_X1   g224(.A(G211gat), .B(G218gat), .Z(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n420), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n359), .B1(new_n406), .B2(KEYINPUT29), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n416), .A2(new_n360), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT76), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT76), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n430), .A2(new_n434), .A3(new_n427), .A4(new_n431), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n429), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G8gat), .B(G36gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(G64gat), .B(G92gat), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n437), .B(new_n438), .Z(new_n439));
  NAND4_X1  g238(.A1(new_n436), .A2(KEYINPUT77), .A3(KEYINPUT30), .A4(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT77), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n429), .A2(new_n433), .A3(new_n435), .A4(new_n439), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT30), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n429), .A2(new_n433), .A3(new_n435), .ZN(new_n445));
  INV_X1    g244(.A(new_n439), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n442), .A2(new_n443), .ZN(new_n448));
  AND4_X1   g247(.A1(new_n440), .A2(new_n444), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n358), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G78gat), .B(G106gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(G22gat), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n313), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n428), .B1(KEYINPUT29), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT29), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT3), .B1(new_n427), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n455), .B1(new_n457), .B2(new_n304), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n458), .A2(G228gat), .A3(G233gat), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT87), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(G228gat), .A2(G233gat), .ZN(new_n462));
  OR2_X1    g261(.A1(new_n424), .A2(new_n426), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n424), .A2(new_n426), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(new_n456), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT86), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n312), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n465), .A2(new_n466), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n331), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n428), .B(KEYINPUT87), .C1(KEYINPUT29), .C2(new_n454), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n461), .A2(new_n462), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n459), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT31), .B(G50gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n473), .A2(new_n474), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n453), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n477), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n479), .A2(new_n452), .A3(new_n475), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n450), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT36), .ZN(new_n483));
  NAND2_X1  g282(.A1(G227gat), .A2(G233gat), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n394), .A2(new_n401), .A3(KEYINPUT25), .A4(new_n402), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n486), .B1(new_n388), .B2(new_n390), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n399), .A2(new_n487), .B1(new_n396), .B2(new_n397), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT68), .B1(new_n488), .B2(new_n379), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT68), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n490), .B(new_n411), .C1(new_n414), .C2(new_n415), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n301), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n330), .B1(new_n416), .B2(KEYINPUT68), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n485), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT32), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT33), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT69), .B(G71gat), .ZN(new_n498));
  INV_X1    g297(.A(G99gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(G15gat), .B(G43gat), .Z(new_n501));
  XOR2_X1   g300(.A(new_n500), .B(new_n501), .Z(new_n502));
  NAND3_X1  g301(.A1(new_n495), .A2(new_n497), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(KEYINPUT70), .A2(KEYINPUT34), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(KEYINPUT70), .A2(KEYINPUT34), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n491), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n493), .B1(new_n508), .B2(new_n330), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n507), .B1(new_n509), .B2(new_n484), .ZN(new_n510));
  NOR4_X1   g309(.A1(new_n492), .A2(new_n493), .A3(new_n485), .A4(new_n505), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n502), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n494), .B(KEYINPUT32), .C1(new_n496), .C2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n503), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT72), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n512), .B1(new_n503), .B2(new_n514), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI211_X1 g317(.A(KEYINPUT72), .B(new_n512), .C1(new_n503), .C2(new_n514), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n483), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n514), .ZN(new_n521));
  INV_X1    g320(.A(new_n512), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT71), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n515), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n517), .A2(KEYINPUT71), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT36), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n482), .A2(new_n520), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT88), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT88), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n482), .A2(new_n520), .A3(new_n526), .A4(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT37), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n439), .B1(new_n436), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT90), .B(KEYINPUT38), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n430), .A2(new_n431), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n531), .B1(new_n534), .B2(new_n428), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n420), .A2(new_n427), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n532), .A2(new_n537), .B1(new_n436), .B2(new_n439), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n436), .A2(new_n531), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n446), .B1(new_n445), .B2(KEYINPUT37), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n533), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n538), .A2(new_n349), .A3(new_n357), .A4(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n481), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT40), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n315), .B1(new_n309), .B2(new_n314), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT39), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n345), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n307), .A2(new_n315), .A3(new_n324), .ZN(new_n548));
  INV_X1    g347(.A(new_n314), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n549), .B1(new_n302), .B2(new_n308), .ZN(new_n550));
  OAI211_X1 g349(.A(KEYINPUT39), .B(new_n548), .C1(new_n550), .C2(new_n315), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n340), .A2(new_n345), .B1(new_n544), .B2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n440), .A2(new_n444), .A3(new_n447), .A4(new_n448), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT89), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n552), .B2(new_n544), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n547), .A2(new_n551), .A3(KEYINPUT89), .A4(KEYINPUT40), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n553), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n543), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n528), .A2(new_n530), .A3(new_n560), .ZN(new_n561));
  AND3_X1   g360(.A1(new_n503), .A2(new_n514), .A3(new_n512), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n562), .B1(KEYINPUT71), .B2(new_n517), .ZN(new_n563));
  INV_X1    g362(.A(new_n525), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n543), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT35), .B1(new_n565), .B2(new_n450), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT91), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n450), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n358), .A2(new_n449), .A3(KEYINPUT91), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n516), .A2(new_n517), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n521), .A2(new_n522), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n571), .A2(KEYINPUT72), .A3(new_n515), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n481), .A2(KEYINPUT35), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n568), .A2(new_n569), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n566), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n249), .B1(new_n561), .B2(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(G134gat), .B(G162gat), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n220), .A2(new_n221), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT102), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT7), .ZN(new_n582));
  NAND2_X1  g381(.A1(G85gat), .A2(G92gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n582), .B(new_n583), .Z(new_n584));
  INV_X1    g383(.A(KEYINPUT8), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n585), .B1(new_n586), .B2(KEYINPUT103), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n587), .B1(KEYINPUT103), .B2(new_n586), .ZN(new_n588));
  XOR2_X1   g387(.A(KEYINPUT104), .B(G85gat), .Z(new_n589));
  INV_X1    g388(.A(G92gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n584), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G99gat), .B(G106gat), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n584), .A2(new_n595), .A3(new_n588), .A4(new_n591), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n580), .B(new_n597), .C1(new_n224), .C2(new_n225), .ZN(new_n598));
  INV_X1    g397(.A(new_n597), .ZN(new_n599));
  NAND2_X1  g398(.A1(G232gat), .A2(G233gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT100), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n599), .A2(new_n220), .B1(KEYINPUT41), .B2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n598), .A2(KEYINPUT105), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n605), .A2(KEYINPUT101), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n602), .A2(KEYINPUT41), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT105), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n580), .A2(new_n597), .ZN(new_n610));
  INV_X1    g409(.A(new_n225), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n610), .B1(new_n611), .B2(new_n223), .ZN(new_n612));
  INV_X1    g411(.A(new_n603), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n609), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n598), .A2(KEYINPUT105), .A3(new_n603), .ZN(new_n615));
  INV_X1    g414(.A(new_n604), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n606), .A2(new_n608), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n608), .B1(new_n606), .B2(new_n617), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n579), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n606), .A2(new_n617), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n607), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n617), .A3(new_n608), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n622), .A2(new_n578), .A3(new_n623), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g424(.A1(G71gat), .A2(G78gat), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n626), .A2(KEYINPUT9), .ZN(new_n627));
  INV_X1    g426(.A(G64gat), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n628), .A2(G57gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(G57gat), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT98), .ZN(new_n632));
  NOR2_X1   g431(.A1(G71gat), .A2(G78gat), .ZN(new_n633));
  OAI22_X1  g432(.A1(new_n627), .A2(new_n632), .B1(new_n626), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n631), .B(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n635), .A2(KEYINPUT21), .ZN(new_n636));
  NAND2_X1  g435(.A1(G231gat), .A2(G233gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(G127gat), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n206), .B1(new_n635), .B2(KEYINPUT21), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G183gat), .B(G211gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT99), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n644));
  INV_X1    g443(.A(G155gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n643), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n641), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n625), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(G120gat), .B(G148gat), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT108), .ZN(new_n651));
  XNOR2_X1  g450(.A(G176gat), .B(G204gat), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n651), .B(new_n652), .Z(new_n653));
  NAND2_X1  g452(.A1(G230gat), .A2(G233gat), .ZN(new_n654));
  INV_X1    g453(.A(new_n635), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n597), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n635), .A2(new_n594), .A3(new_n596), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n597), .A2(new_n655), .A3(KEYINPUT106), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT10), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT10), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n654), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n659), .A2(G230gat), .A3(G233gat), .A4(new_n660), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n653), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT109), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT107), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n665), .A2(new_n668), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n669), .A2(new_n664), .A3(new_n670), .A4(new_n653), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n649), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n577), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n358), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g476(.A1(new_n674), .A2(new_n554), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT16), .B(G8gat), .Z(new_n679));
  AND2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(G8gat), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(KEYINPUT42), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n683), .B1(KEYINPUT42), .B2(new_n680), .ZN(G1325gat));
  INV_X1    g483(.A(G15gat), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n674), .A2(new_n685), .A3(new_n573), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n483), .B1(new_n563), .B2(new_n564), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT36), .B1(new_n572), .B2(new_n570), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n674), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n686), .B1(new_n691), .B2(new_n685), .ZN(G1326gat));
  NAND2_X1  g491(.A1(new_n674), .A2(new_n481), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT43), .B(G22gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1327gat));
  AOI21_X1  g494(.A(new_n625), .B1(new_n561), .B2(new_n576), .ZN(new_n696));
  INV_X1    g495(.A(new_n648), .ZN(new_n697));
  INV_X1    g496(.A(new_n672), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n249), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n701), .A2(G29gat), .A3(new_n358), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT45), .Z(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n689), .A2(new_n705), .A3(new_n482), .A4(new_n560), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n560), .A2(new_n482), .A3(new_n520), .A4(new_n526), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT110), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n706), .A2(new_n708), .B1(new_n566), .B2(new_n575), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n704), .B1(new_n709), .B2(new_n625), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n561), .A2(new_n576), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n620), .A2(new_n624), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(KEYINPUT44), .A3(new_n712), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n710), .A2(new_n713), .A3(new_n700), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(G29gat), .B1(new_n715), .B2(new_n358), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n703), .A2(new_n716), .ZN(G1328gat));
  NOR3_X1   g516(.A1(new_n701), .A2(G36gat), .A3(new_n449), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT46), .ZN(new_n719));
  OAI21_X1  g518(.A(G36gat), .B1(new_n715), .B2(new_n449), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(G1329gat));
  NAND4_X1  g520(.A1(new_n710), .A2(new_n713), .A3(new_n690), .A4(new_n700), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(G43gat), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT113), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT112), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n243), .A2(new_n239), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n247), .A2(new_n248), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n573), .ZN(new_n729));
  NOR4_X1   g528(.A1(new_n699), .A2(new_n625), .A3(G43gat), .A4(new_n729), .ZN(new_n730));
  AND4_X1   g529(.A1(new_n725), .A2(new_n711), .A3(new_n728), .A4(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n725), .B1(new_n577), .B2(new_n730), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n724), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n711), .A2(new_n728), .A3(new_n730), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT112), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n577), .A2(new_n725), .A3(new_n730), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(KEYINPUT113), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n723), .A2(new_n733), .A3(new_n737), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT111), .B(KEYINPUT47), .Z(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n723), .B(KEYINPUT47), .C1(new_n732), .C2(new_n731), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT114), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT114), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n740), .A2(new_n744), .A3(new_n741), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(G1330gat));
  NAND3_X1  g545(.A1(new_n714), .A2(G50gat), .A3(new_n481), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n701), .A2(new_n543), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(G50gat), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(G1331gat));
  NOR4_X1   g550(.A1(new_n709), .A2(new_n728), .A3(new_n649), .A4(new_n698), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n675), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n554), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n756));
  XOR2_X1   g555(.A(KEYINPUT49), .B(G64gat), .Z(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n755), .B2(new_n757), .ZN(G1333gat));
  NAND2_X1  g557(.A1(new_n752), .A2(new_n690), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n729), .A2(G71gat), .ZN(new_n760));
  AOI22_X1  g559(.A1(new_n759), .A2(G71gat), .B1(new_n752), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g561(.A1(new_n752), .A2(new_n481), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g563(.A1(new_n728), .A2(new_n648), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n709), .A2(new_n625), .A3(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT51), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n768), .A2(new_n675), .A3(new_n589), .A4(new_n672), .ZN(new_n769));
  AND4_X1   g568(.A1(new_n672), .A2(new_n710), .A3(new_n713), .A4(new_n765), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(new_n675), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n589), .B2(new_n771), .ZN(G1336gat));
  NAND4_X1  g571(.A1(new_n768), .A2(new_n590), .A3(new_n554), .A4(new_n672), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n554), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G92gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT52), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n773), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1337gat));
  NAND4_X1  g579(.A1(new_n768), .A2(new_n499), .A3(new_n573), .A4(new_n672), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n770), .A2(new_n690), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G99gat), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n782), .A2(new_n783), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n781), .B1(new_n785), .B2(new_n786), .ZN(G1338gat));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n481), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT53), .B1(new_n788), .B2(G106gat), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT118), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n543), .A2(G106gat), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n672), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n768), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n790), .B1(new_n768), .B2(new_n793), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n789), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797));
  XOR2_X1   g596(.A(new_n792), .B(KEYINPUT117), .Z(new_n798));
  AOI22_X1  g597(.A1(G106gat), .A2(new_n788), .B1(new_n768), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n796), .B1(new_n797), .B2(new_n799), .ZN(G1339gat));
  AOI21_X1  g599(.A(new_n227), .B1(new_n226), .B2(new_n228), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n236), .A2(new_n237), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n233), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n726), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n672), .ZN(new_n805));
  OR3_X1    g604(.A1(new_n661), .A2(new_n654), .A3(new_n663), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n806), .A2(KEYINPUT54), .A3(new_n664), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n808), .B(new_n654), .C1(new_n661), .C2(new_n663), .ZN(new_n809));
  INV_X1    g608(.A(new_n653), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n807), .A2(new_n811), .A3(KEYINPUT55), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT119), .B1(new_n812), .B2(new_n671), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT55), .B1(new_n807), .B2(new_n811), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n812), .A2(KEYINPUT119), .A3(new_n671), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(new_n728), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n712), .B1(new_n805), .B2(new_n817), .ZN(new_n818));
  AND4_X1   g617(.A1(new_n712), .A2(new_n804), .A3(new_n815), .A4(new_n816), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n697), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n673), .A2(new_n249), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n358), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n565), .A2(new_n554), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(G113gat), .B1(new_n824), .B2(new_n728), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n481), .B1(new_n820), .B2(new_n821), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n826), .A2(new_n675), .A3(new_n449), .A4(new_n573), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT120), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n249), .A2(new_n288), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n825), .B1(new_n828), .B2(new_n829), .ZN(G1340gat));
  AOI21_X1  g629(.A(G120gat), .B1(new_n824), .B2(new_n672), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n698), .A2(new_n286), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n828), .B2(new_n832), .ZN(G1341gat));
  XNOR2_X1  g632(.A(KEYINPUT67), .B(G127gat), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n697), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n824), .A2(new_n648), .ZN(new_n836));
  AOI22_X1  g635(.A1(new_n828), .A2(new_n835), .B1(new_n836), .B2(new_n834), .ZN(G1342gat));
  AOI21_X1  g636(.A(new_n297), .B1(new_n828), .B2(new_n712), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n824), .A2(new_n297), .A3(new_n712), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT56), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n838), .A2(new_n840), .ZN(G1343gat));
  NOR3_X1   g640(.A1(new_n690), .A2(new_n358), .A3(new_n554), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n671), .B(new_n812), .C1(new_n814), .C2(new_n843), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n814), .A2(new_n843), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n249), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n672), .A2(new_n726), .A3(new_n803), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n625), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n712), .A2(new_n804), .A3(new_n816), .A4(new_n815), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n648), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n649), .A2(new_n728), .A3(new_n672), .ZN(new_n851));
  OAI211_X1 g650(.A(KEYINPUT57), .B(new_n481), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n543), .B1(new_n820), .B2(new_n821), .ZN(new_n853));
  XNOR2_X1  g652(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  OAI22_X1  g654(.A1(new_n852), .A2(KEYINPUT123), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n844), .A2(new_n845), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n728), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n712), .B1(new_n859), .B2(new_n805), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n697), .B1(new_n860), .B2(new_n819), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n543), .B1(new_n861), .B2(new_n821), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n857), .B1(new_n862), .B2(KEYINPUT57), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n728), .B(new_n842), .C1(new_n856), .C2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n278), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AND4_X1   g665(.A1(new_n449), .A2(new_n822), .A3(new_n481), .A4(new_n689), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n262), .A3(new_n728), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT58), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT58), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n866), .A2(new_n871), .A3(new_n868), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(G1344gat));
  AND2_X1   g672(.A1(new_n853), .A2(new_n855), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n862), .A2(KEYINPUT57), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n842), .A2(new_n672), .ZN(new_n877));
  OAI21_X1  g676(.A(G148gat), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT59), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n254), .A2(KEYINPUT59), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n842), .B1(new_n856), .B2(new_n863), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n881), .B2(new_n698), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n867), .A2(new_n254), .A3(new_n672), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(G1345gat));
  OAI21_X1  g684(.A(G155gat), .B1(new_n881), .B2(new_n697), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n867), .A2(new_n645), .A3(new_n648), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1346gat));
  NAND2_X1  g687(.A1(new_n712), .A2(G162gat), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n881), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(G162gat), .B1(new_n867), .B2(new_n712), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(G1347gat));
  NAND2_X1  g692(.A1(new_n820), .A2(new_n821), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n675), .A2(new_n449), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n565), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(G169gat), .B1(new_n899), .B2(new_n728), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n826), .A2(new_n573), .A3(new_n895), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n249), .A2(new_n392), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(G1348gat));
  NOR3_X1   g702(.A1(new_n898), .A2(G176gat), .A3(new_n698), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n901), .A2(new_n672), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(G176gat), .ZN(new_n906));
  XOR2_X1   g705(.A(new_n906), .B(KEYINPUT124), .Z(G1349gat));
  AOI21_X1  g706(.A(new_n369), .B1(new_n901), .B2(new_n648), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n648), .A2(new_n377), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n899), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n910), .B(new_n911), .ZN(G1350gat));
  NAND3_X1  g711(.A1(new_n899), .A2(new_n373), .A3(new_n712), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n901), .A2(new_n712), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(G190gat), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n915), .A2(KEYINPUT61), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(KEYINPUT61), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(G1351gat));
  NOR2_X1   g717(.A1(new_n690), .A2(new_n896), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n853), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(G197gat), .B1(new_n920), .B2(new_n728), .ZN(new_n921));
  INV_X1    g720(.A(new_n876), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n919), .B(KEYINPUT126), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n728), .A2(G197gat), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n921), .B1(new_n925), .B2(new_n926), .ZN(G1352gat));
  OAI21_X1  g726(.A(G204gat), .B1(new_n924), .B2(new_n698), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n929));
  AOI21_X1  g728(.A(G204gat), .B1(new_n929), .B2(KEYINPUT62), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n920), .A2(new_n672), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n929), .A2(KEYINPUT62), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n931), .B(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n928), .A2(new_n933), .ZN(G1353gat));
  INV_X1    g733(.A(G211gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n920), .A2(new_n935), .A3(new_n648), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n648), .ZN(new_n937));
  OAI21_X1  g736(.A(G211gat), .B1(new_n876), .B2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT63), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n938), .A2(new_n939), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n936), .B1(new_n940), .B2(new_n941), .ZN(G1354gat));
  OAI21_X1  g741(.A(G218gat), .B1(new_n924), .B2(new_n625), .ZN(new_n943));
  INV_X1    g742(.A(G218gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n920), .A2(new_n944), .A3(new_n712), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1355gat));
endmodule


