//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n567, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162, new_n1163;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT66), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n454), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  XOR2_X1   g044(.A(new_n469), .B(KEYINPUT67), .Z(new_n470));
  AOI21_X1  g045(.A(new_n462), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n462), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n472), .B(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n464), .A2(new_n466), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G137), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n475), .A2(KEYINPUT69), .A3(new_n478), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n471), .B1(new_n481), .B2(new_n482), .ZN(G160));
  NOR2_X1   g058(.A1(new_n476), .A2(new_n462), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n477), .A2(G136), .ZN(new_n486));
  NOR2_X1   g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(new_n462), .B2(G112), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n485), .B(new_n486), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT70), .ZN(G162));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n467), .A2(new_n462), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n477), .A2(KEYINPUT4), .A3(G138), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n467), .A2(G126), .A3(G2105), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G114), .C2(new_n462), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n496), .A2(new_n500), .ZN(G164));
  XNOR2_X1  g076(.A(KEYINPUT71), .B(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT6), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(KEYINPUT5), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n504), .A2(KEYINPUT72), .A3(G543), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n511), .A2(KEYINPUT6), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n503), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  XOR2_X1   g088(.A(KEYINPUT73), .B(G88), .Z(new_n514));
  NAND3_X1  g089(.A1(new_n503), .A2(G543), .A3(new_n512), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n518), .A2(new_n502), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n517), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  INV_X1    g097(.A(G51), .ZN(new_n523));
  INV_X1    g098(.A(G89), .ZN(new_n524));
  OAI221_X1 g099(.A(new_n522), .B1(new_n515), .B2(new_n523), .C1(new_n524), .C2(new_n513), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n504), .A2(KEYINPUT72), .A3(G543), .ZN(new_n527));
  AOI21_X1  g102(.A(KEYINPUT72), .B1(new_n504), .B2(G543), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT74), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n510), .A2(KEYINPUT74), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n533), .A2(G63), .A3(G651), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n525), .A2(new_n534), .ZN(G168));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  INV_X1    g111(.A(G52), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n513), .A2(new_n536), .B1(new_n515), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT75), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n533), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n502), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  INV_X1    g118(.A(new_n502), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n545), .B1(new_n531), .B2(new_n532), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n544), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(KEYINPUT76), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n503), .A2(new_n510), .A3(new_n512), .ZN(new_n551));
  AND3_X1   g126(.A1(new_n503), .A2(G543), .A3(new_n512), .ZN(new_n552));
  AOI22_X1  g127(.A1(G81), .A2(new_n551), .B1(new_n552), .B2(G43), .ZN(new_n553));
  AOI211_X1 g128(.A(new_n530), .B(new_n505), .C1(new_n508), .C2(new_n509), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n508), .A2(new_n509), .ZN(new_n555));
  AOI21_X1  g130(.A(KEYINPUT74), .B1(new_n555), .B2(new_n526), .ZN(new_n556));
  OAI21_X1  g131(.A(G56), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(new_n547), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT76), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n558), .A2(new_n559), .A3(new_n544), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n550), .A2(new_n553), .A3(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n550), .A2(KEYINPUT77), .A3(new_n560), .A4(new_n553), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  AND3_X1   g141(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G36), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(G188));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n529), .B2(new_n573), .ZN(new_n574));
  XOR2_X1   g149(.A(new_n574), .B(KEYINPUT79), .Z(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G651), .ZN(new_n576));
  NAND2_X1  g151(.A1(KEYINPUT78), .A2(KEYINPUT9), .ZN(new_n577));
  NOR2_X1   g152(.A1(KEYINPUT78), .A2(KEYINPUT9), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n552), .A2(G53), .A3(new_n577), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n552), .A2(G53), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(new_n578), .B1(G91), .B2(new_n551), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n576), .A2(new_n580), .A3(new_n582), .ZN(G299));
  INV_X1    g158(.A(G168), .ZN(G286));
  INV_X1    g159(.A(G166), .ZN(G303));
  AOI22_X1  g160(.A1(G87), .A2(new_n551), .B1(new_n552), .B2(G49), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n533), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(new_n510), .A2(G61), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n502), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n591), .A2(KEYINPUT80), .ZN(new_n592));
  AOI22_X1  g167(.A1(G86), .A2(new_n551), .B1(new_n552), .B2(G48), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(KEYINPUT80), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n533), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT81), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(new_n544), .ZN(new_n598));
  AOI22_X1  g173(.A1(G85), .A2(new_n551), .B1(new_n552), .B2(G47), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n510), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n602));
  XOR2_X1   g177(.A(new_n602), .B(KEYINPUT83), .Z(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(G54), .B2(new_n552), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT82), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n551), .A2(new_n605), .A3(G92), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT82), .B1(new_n513), .B2(new_n607), .ZN(new_n608));
  AND3_X1   g183(.A1(new_n606), .A2(KEYINPUT10), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g184(.A(KEYINPUT10), .B1(new_n606), .B2(new_n608), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AND2_X1   g186(.A1(new_n604), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n601), .B1(new_n612), .B2(G868), .ZN(G321));
  XNOR2_X1  g188(.A(G321), .B(KEYINPUT84), .ZN(G284));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n574), .B(KEYINPUT79), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n616), .A2(new_n511), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n582), .A2(new_n580), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n615), .B1(new_n619), .B2(G868), .ZN(G297));
  OAI21_X1  g195(.A(new_n615), .B1(new_n619), .B2(G868), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n612), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n604), .A2(new_n611), .ZN(new_n624));
  OAI21_X1  g199(.A(G868), .B1(new_n624), .B2(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n565), .B2(G868), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n474), .A2(new_n467), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  INV_X1    g204(.A(G2100), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT85), .B(KEYINPUT13), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n484), .A2(G123), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n477), .A2(G135), .ZN(new_n635));
  NOR2_X1   g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  OAI21_X1  g211(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n634), .B(new_n635), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2096), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n633), .A2(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2435), .ZN(new_n642));
  XOR2_X1   g217(.A(G2427), .B(G2438), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT14), .ZN(new_n645));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT86), .B(KEYINPUT16), .Z(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2443), .B(G2446), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(G14), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT87), .ZN(G401));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  XOR2_X1   g231(.A(G2067), .B(G2678), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n656), .B1(new_n660), .B2(KEYINPUT18), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2096), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(new_n630), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n658), .A2(new_n659), .ZN(new_n665));
  AOI21_X1  g240(.A(KEYINPUT18), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n670), .A2(new_n671), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n677), .A2(new_n669), .A3(new_n672), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n675), .B(new_n678), .C1(new_n669), .C2(new_n677), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT21), .B(G1986), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT22), .B(G1981), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G229));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G6), .ZN(new_n687));
  AND3_X1   g262(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(new_n686), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT32), .B(G1981), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT92), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n686), .A2(G22), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G166), .B2(new_n686), .ZN(new_n694));
  INV_X1    g269(.A(G1971), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(G16), .A2(G23), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n586), .A2(new_n587), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(G16), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT33), .B(G1976), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n692), .A2(new_n696), .A3(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT34), .Z(new_n703));
  NAND2_X1  g278(.A1(G290), .A2(G16), .ZN(new_n704));
  INV_X1    g279(.A(G24), .ZN(new_n705));
  OAI21_X1  g280(.A(KEYINPUT90), .B1(new_n705), .B2(G16), .ZN(new_n706));
  OR3_X1    g281(.A1(new_n705), .A2(KEYINPUT90), .A3(G16), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n704), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT91), .B(G1986), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n484), .A2(G119), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n477), .A2(G131), .ZN(new_n712));
  NOR2_X1   g287(.A1(G95), .A2(G2105), .ZN(new_n713));
  OAI21_X1  g288(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n711), .B(new_n712), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  AND2_X1   g290(.A1(KEYINPUT89), .A2(G29), .ZN(new_n716));
  NOR2_X1   g291(.A1(KEYINPUT89), .A2(G29), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  MUX2_X1   g293(.A(G25), .B(new_n715), .S(new_n718), .Z(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT35), .B(G1991), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n719), .B(new_n720), .Z(new_n721));
  NAND3_X1  g296(.A1(new_n703), .A2(new_n710), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT36), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n686), .A2(KEYINPUT23), .A3(G20), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT23), .ZN(new_n725));
  INV_X1    g300(.A(G20), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(G16), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n724), .B(new_n727), .C1(new_n619), .C2(new_n686), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT97), .B(G1956), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT96), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G5), .B2(G16), .ZN(new_n732));
  OR3_X1    g307(.A1(new_n731), .A2(G5), .A3(G16), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n732), .B(new_n733), .C1(G301), .C2(new_n686), .ZN(new_n734));
  INV_X1    g309(.A(G1961), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n718), .A2(G35), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G162), .B2(new_n718), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT29), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(G2090), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n718), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n742), .A2(KEYINPUT28), .A3(G26), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n477), .A2(G140), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT93), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n484), .A2(G128), .ZN(new_n746));
  NOR2_X1   g321(.A1(G104), .A2(G2105), .ZN(new_n747));
  OAI21_X1  g322(.A(G2104), .B1(new_n462), .B2(G116), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G29), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n743), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(KEYINPUT28), .B1(new_n742), .B2(G26), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G2067), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n742), .A2(G27), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G164), .B2(new_n742), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2078), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n739), .A2(G2090), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n686), .A2(G4), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n612), .B2(new_n686), .ZN(new_n763));
  INV_X1    g338(.A(G1348), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n741), .A2(new_n760), .A3(new_n761), .A4(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n565), .A2(new_n686), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n686), .B2(G19), .ZN(new_n768));
  INV_X1    g343(.A(G1341), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  NAND2_X1  g346(.A1(G160), .A2(G29), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT24), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(G34), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(G34), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n742), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(G2084), .B1(new_n772), .B2(new_n776), .ZN(new_n777));
  AND3_X1   g352(.A1(new_n772), .A2(G2084), .A3(new_n776), .ZN(new_n778));
  NOR2_X1   g353(.A1(G16), .A2(G21), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G168), .B2(G16), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n777), .B(new_n778), .C1(G1966), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n474), .A2(G105), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n477), .A2(G141), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n484), .A2(G129), .ZN(new_n784));
  NAND3_X1  g359(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT26), .Z(new_n786));
  NAND4_X1  g361(.A1(new_n782), .A2(new_n783), .A3(new_n784), .A4(new_n786), .ZN(new_n787));
  MUX2_X1   g362(.A(G32), .B(new_n787), .S(G29), .Z(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT27), .B(G1996), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n780), .A2(G1966), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n638), .A2(new_n742), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT30), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n751), .B1(new_n793), .B2(G28), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT95), .Z(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n793), .B2(G28), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n791), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT31), .B(G11), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n781), .A2(new_n790), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NOR4_X1   g374(.A1(new_n766), .A2(new_n770), .A3(new_n771), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n477), .A2(G139), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT94), .Z(new_n802));
  NAND3_X1  g377(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT25), .Z(new_n804));
  AOI22_X1  g379(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n802), .B(new_n804), .C1(new_n462), .C2(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G33), .B(new_n806), .S(G29), .Z(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(G2072), .Z(new_n808));
  NAND4_X1  g383(.A1(new_n723), .A2(new_n730), .A3(new_n800), .A4(new_n808), .ZN(G150));
  INV_X1    g384(.A(G150), .ZN(G311));
  INV_X1    g385(.A(G93), .ZN(new_n811));
  INV_X1    g386(.A(G55), .ZN(new_n812));
  OAI22_X1  g387(.A1(new_n513), .A2(new_n811), .B1(new_n515), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n533), .A2(G67), .ZN(new_n814));
  INV_X1    g389(.A(G80), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(new_n507), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n813), .B1(new_n816), .B2(new_n544), .ZN(new_n817));
  INV_X1    g392(.A(G860), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT37), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n624), .A2(new_n622), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n561), .A2(new_n817), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT98), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n561), .A2(KEYINPUT98), .A3(new_n817), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n817), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n559), .B1(new_n558), .B2(new_n544), .ZN(new_n830));
  AOI211_X1 g405(.A(KEYINPUT76), .B(new_n502), .C1(new_n557), .C2(new_n547), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(KEYINPUT77), .B1(new_n832), .B2(new_n553), .ZN(new_n833));
  INV_X1    g408(.A(new_n564), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n829), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n828), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n823), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT39), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT100), .Z(new_n840));
  OAI21_X1  g415(.A(new_n818), .B1(new_n837), .B2(new_n838), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n820), .B1(new_n840), .B2(new_n841), .ZN(G145));
  INV_X1    g417(.A(KEYINPUT101), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n497), .B2(new_n499), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n497), .A2(new_n843), .A3(new_n499), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n496), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n750), .B(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n787), .B(KEYINPUT102), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n806), .A2(KEYINPUT103), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n806), .A2(KEYINPUT103), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n851), .B2(new_n850), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n484), .A2(G130), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n477), .A2(G142), .ZN(new_n856));
  NOR2_X1   g431(.A1(G106), .A2(G2105), .ZN(new_n857));
  OAI21_X1  g432(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n855), .B(new_n856), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n629), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n715), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n854), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n854), .A2(new_n861), .ZN(new_n863));
  XNOR2_X1  g438(.A(G160), .B(new_n638), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(G162), .Z(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n862), .A2(new_n863), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G37), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n861), .A2(KEYINPUT104), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n854), .B(new_n869), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n867), .B(new_n868), .C1(new_n870), .C2(new_n866), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g447(.A1(new_n698), .A2(G303), .ZN(new_n873));
  NAND2_X1  g448(.A1(G288), .A2(G166), .ZN(new_n874));
  AOI21_X1  g449(.A(G305), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n873), .A2(new_n874), .A3(G305), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n876), .A2(new_n599), .A3(new_n598), .A4(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n877), .ZN(new_n879));
  OAI21_X1  g454(.A(G290), .B1(new_n879), .B2(new_n875), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n878), .A2(new_n880), .A3(KEYINPUT106), .A4(new_n881), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n878), .A2(new_n880), .A3(KEYINPUT105), .ZN(new_n883));
  AOI21_X1  g458(.A(KEYINPUT105), .B1(new_n878), .B2(new_n880), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n885), .B1(KEYINPUT105), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n882), .B1(new_n887), .B2(new_n881), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n624), .A2(G559), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n836), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n612), .A2(new_n619), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n624), .A2(G299), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n891), .A2(KEYINPUT41), .A3(new_n892), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT41), .B1(new_n891), .B2(new_n892), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n894), .B1(new_n890), .B2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n888), .B(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(G868), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(G868), .B2(new_n817), .ZN(G295));
  OAI21_X1  g476(.A(new_n900), .B1(G868), .B2(new_n817), .ZN(G331));
  XNOR2_X1  g477(.A(G301), .B(G168), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n561), .A2(KEYINPUT98), .A3(new_n817), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT98), .B1(new_n561), .B2(new_n817), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n817), .B1(new_n563), .B2(new_n564), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(G301), .B(G286), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n828), .A2(new_n835), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n910), .A3(KEYINPUT107), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n828), .A2(new_n835), .A3(new_n909), .A4(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n897), .A3(new_n913), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n908), .A2(new_n910), .A3(new_n892), .A4(new_n891), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n885), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT108), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n868), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n914), .A2(new_n885), .A3(new_n915), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n885), .B1(new_n914), .B2(new_n915), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT108), .B1(new_n922), .B2(G37), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n893), .B1(new_n911), .B2(new_n913), .ZN(new_n927));
  AOI211_X1 g502(.A(new_n896), .B(new_n895), .C1(new_n910), .C2(new_n908), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n917), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(new_n868), .A3(new_n921), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT109), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n929), .A2(new_n932), .A3(new_n868), .A4(new_n921), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n925), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT44), .B1(new_n926), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n924), .A2(KEYINPUT43), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n935), .A2(new_n940), .ZN(G397));
  AND3_X1   g516(.A1(new_n497), .A2(new_n843), .A3(new_n499), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n494), .B(new_n495), .C1(new_n942), .C2(new_n844), .ZN(new_n943));
  INV_X1    g518(.A(G1384), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT45), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n471), .ZN(new_n948));
  INV_X1    g523(.A(new_n482), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT69), .B1(new_n475), .B2(new_n478), .ZN(new_n950));
  OAI211_X1 g525(.A(G40), .B(new_n948), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n750), .B(G2067), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n952), .B1(new_n954), .B2(new_n787), .ZN(new_n955));
  INV_X1    g530(.A(new_n952), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n956), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT46), .ZN(new_n958));
  INV_X1    g533(.A(G1996), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n958), .B1(new_n952), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n955), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT47), .Z(new_n962));
  NAND3_X1  g537(.A1(new_n952), .A2(G1996), .A3(new_n787), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(KEYINPUT110), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n963), .A2(KEYINPUT110), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n953), .B1(G1996), .B2(new_n787), .ZN(new_n966));
  AOI211_X1 g541(.A(new_n964), .B(new_n965), .C1(new_n952), .C2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n715), .A2(new_n720), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n750), .A2(new_n755), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n956), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n715), .A2(new_n720), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n952), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n967), .A2(new_n973), .ZN(new_n974));
  NOR3_X1   g549(.A1(G290), .A2(new_n956), .A3(G1986), .ZN(new_n975));
  XOR2_X1   g550(.A(new_n975), .B(KEYINPUT48), .Z(new_n976));
  AOI211_X1 g551(.A(new_n962), .B(new_n971), .C1(new_n974), .C2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT49), .ZN(new_n978));
  NAND2_X1  g553(.A1(G305), .A2(G1981), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(G305), .A2(G1981), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n981), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n983), .A2(KEYINPUT49), .A3(new_n979), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n945), .A2(new_n951), .ZN(new_n985));
  INV_X1    g560(.A(G8), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n982), .A2(new_n984), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1976), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT52), .B1(G288), .B2(new_n989), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n987), .B(new_n990), .C1(new_n989), .C2(G288), .ZN(new_n991));
  OAI221_X1 g566(.A(G8), .B1(G288), .B2(new_n989), .C1(new_n945), .C2(new_n951), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT52), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n988), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n988), .A2(new_n991), .A3(new_n993), .A4(KEYINPUT113), .ZN(new_n997));
  INV_X1    g572(.A(G40), .ZN(new_n998));
  AOI211_X1 g573(.A(new_n998), .B(new_n471), .C1(new_n481), .C2(new_n482), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n943), .A2(new_n1000), .A3(new_n944), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n944), .B1(new_n496), .B2(new_n500), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT50), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT111), .B(G2090), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n943), .A2(KEYINPUT45), .A3(new_n944), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1002), .A2(new_n946), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n999), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n695), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n986), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(G166), .A2(new_n986), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT55), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n996), .A2(new_n997), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT120), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1013), .A2(KEYINPUT112), .A3(new_n1015), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT45), .B1(new_n943), .B2(new_n944), .ZN(new_n1024));
  OAI211_X1 g599(.A(KEYINPUT45), .B(new_n944), .C1(new_n496), .C2(new_n500), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n1024), .A2(new_n1026), .A3(new_n951), .ZN(new_n1027));
  INV_X1    g602(.A(G2084), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .A4(new_n1028), .ZN(new_n1029));
  OAI22_X1  g604(.A1(new_n1027), .A2(G1966), .B1(new_n1029), .B2(KEYINPUT118), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(KEYINPUT118), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(G8), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1033), .A2(G286), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT120), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n996), .A2(new_n1016), .A3(new_n1035), .A4(new_n997), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1018), .A2(new_n1023), .A3(new_n1034), .A4(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT63), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n994), .A2(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n988), .A2(new_n991), .A3(new_n993), .A4(KEYINPUT117), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1015), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1000), .B(new_n944), .C1(new_n496), .C2(new_n500), .ZN(new_n1045));
  NAND3_X1  g620(.A1(G160), .A2(new_n1045), .A3(G40), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1000), .B1(new_n943), .B2(new_n944), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1047), .A2(KEYINPUT115), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1051), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(new_n1052), .A3(new_n1007), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1053), .A2(KEYINPUT116), .A3(new_n1012), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G8), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT116), .B1(new_n1053), .B2(new_n1012), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1044), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1043), .A2(new_n1023), .A3(new_n1057), .A4(new_n1034), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1058), .A2(new_n1059), .A3(new_n1038), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1059), .B1(new_n1058), .B2(new_n1038), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1039), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1023), .A2(new_n1043), .A3(new_n1057), .ZN(new_n1063));
  INV_X1    g638(.A(G2078), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n999), .A2(new_n1009), .A3(new_n1010), .A4(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1065), .A2(new_n1066), .B1(new_n1004), .B2(new_n735), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1024), .A2(new_n951), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1068), .A2(KEYINPUT53), .A3(new_n1064), .A4(new_n1009), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(G301), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(G1961), .B2(new_n1005), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n1073));
  NOR4_X1   g648(.A1(new_n1024), .A2(new_n1026), .A3(new_n951), .A4(G2078), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1073), .B1(new_n1074), .B2(KEYINPUT124), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n947), .A2(new_n1064), .A3(new_n999), .A4(new_n1025), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT124), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1072), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1070), .B1(new_n1079), .B2(G301), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT126), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1068), .A2(KEYINPUT124), .A3(new_n1064), .A4(new_n1025), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1078), .A2(KEYINPUT53), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(G301), .B1(new_n1084), .B2(new_n1067), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1070), .ZN(new_n1086));
  OAI211_X1 g661(.A(KEYINPUT126), .B(new_n1081), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1082), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1956), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT56), .B(G2072), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n999), .A2(new_n1009), .A3(new_n1010), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n576), .A2(new_n1095), .A3(new_n580), .A4(new_n582), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT57), .B1(new_n617), .B2(new_n618), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1004), .A2(new_n764), .B1(new_n985), .B2(new_n755), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1091), .A2(new_n1097), .A3(new_n1096), .A4(new_n1093), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(new_n612), .A3(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n612), .B1(new_n1100), .B2(KEYINPUT60), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT121), .B1(new_n1100), .B2(KEYINPUT60), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1100), .A2(KEYINPUT121), .A3(KEYINPUT60), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1108), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1104), .B1(new_n1110), .B2(new_n1106), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT61), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1099), .A2(new_n1113), .A3(new_n1102), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1113), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT58), .B(G1341), .ZN(new_n1116));
  OAI22_X1  g691(.A1(new_n1011), .A2(G1996), .B1(new_n985), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n565), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1118), .A2(KEYINPUT59), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1118), .A2(KEYINPUT59), .ZN(new_n1120));
  OAI22_X1  g695(.A1(new_n1114), .A2(new_n1115), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1099), .B(new_n1103), .C1(new_n1112), .C2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g697(.A(G8), .B(G286), .C1(new_n1030), .C2(new_n1032), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1123), .B(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1068), .A2(new_n1025), .ZN(new_n1126));
  INV_X1    g701(.A(G1966), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1029), .A2(KEYINPUT118), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1128), .A2(new_n1129), .A3(G168), .A4(new_n1031), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(KEYINPUT51), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1130), .A2(G8), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1132), .B1(new_n1130), .B2(G8), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1131), .A2(KEYINPUT51), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1125), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1081), .B1(new_n1079), .B2(G301), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1139));
  XOR2_X1   g714(.A(new_n1139), .B(KEYINPUT127), .Z(new_n1140));
  OAI21_X1  g715(.A(new_n1138), .B1(new_n1140), .B2(G301), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1089), .A2(new_n1122), .A3(new_n1137), .A4(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1136), .A2(new_n1133), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1123), .B(KEYINPUT122), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT62), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1125), .A2(new_n1146), .A3(new_n1133), .A4(new_n1136), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1145), .A2(new_n1147), .A3(new_n1085), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1063), .B1(new_n1142), .B2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(G288), .A2(G1976), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT114), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1151), .B1(new_n982), .B2(new_n984), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n987), .B1(new_n1152), .B2(new_n981), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n996), .A2(new_n997), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1153), .B1(new_n1023), .B2(new_n1154), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1062), .A2(new_n1149), .A3(new_n1155), .ZN(new_n1156));
  XOR2_X1   g731(.A(G290), .B(G1986), .Z(new_n1157));
  OAI21_X1  g732(.A(new_n974), .B1(new_n956), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n977), .B1(new_n1156), .B2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g734(.A1(G229), .A2(G227), .ZN(new_n1161));
  NOR2_X1   g735(.A1(G401), .A2(new_n460), .ZN(new_n1162));
  AND2_X1   g736(.A1(new_n871), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g737(.A1(new_n938), .A2(new_n1161), .A3(new_n1163), .ZN(G225));
  INV_X1    g738(.A(G225), .ZN(G308));
endmodule


