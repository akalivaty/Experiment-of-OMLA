//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n567, new_n568, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n624, new_n625, new_n626, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1200, new_n1201, new_n1202;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g026(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  XNOR2_X1  g043(.A(new_n468), .B(KEYINPUT69), .ZN(new_n469));
  OAI21_X1  g044(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g047(.A(KEYINPUT68), .B(G125), .C1(new_n461), .C2(new_n462), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n467), .B1(new_n474), .B2(new_n465), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n464), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n487), .A2(new_n465), .A3(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n486), .B1(new_n463), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n477), .A2(G126), .A3(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR3_X1   g066(.A1(new_n491), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n477), .A2(KEYINPUT4), .A3(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n489), .A2(new_n490), .A3(new_n493), .A4(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  OR2_X1    g072(.A1(KEYINPUT71), .A2(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT71), .A2(G651), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT73), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G62), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n501), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT74), .ZN(new_n510));
  OR2_X1    g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT72), .B1(new_n512), .B2(KEYINPUT6), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(new_n515), .A3(G651), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n498), .A2(KEYINPUT6), .A3(new_n499), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n506), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n517), .A2(G543), .A3(new_n518), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G50), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n509), .A2(new_n510), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n511), .A2(new_n522), .A3(new_n525), .A4(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  XNOR2_X1  g103(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n529), .B(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(G63), .A2(G651), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n531), .B1(new_n506), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n521), .A2(G89), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n524), .A2(G51), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n517), .A2(G52), .A3(G543), .A4(new_n518), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n517), .A2(G90), .A3(new_n506), .A4(new_n518), .ZN(new_n540));
  INV_X1    g115(.A(new_n505), .ZN(new_n541));
  AOI21_X1  g116(.A(G543), .B1(KEYINPUT73), .B2(KEYINPUT5), .ZN(new_n542));
  OAI21_X1  g117(.A(G64), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n501), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n539), .B(new_n540), .C1(new_n545), .C2(KEYINPUT76), .ZN(new_n546));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n504), .B2(new_n505), .ZN(new_n548));
  INV_X1    g123(.A(new_n544), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n500), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n538), .B1(new_n546), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n539), .A2(new_n540), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n545), .A2(KEYINPUT76), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n550), .A2(new_n551), .ZN(new_n556));
  NAND4_X1  g131(.A1(new_n554), .A2(KEYINPUT77), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n553), .A2(new_n557), .ZN(G171));
  NAND2_X1  g133(.A1(new_n521), .A2(G81), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n560), .A2(new_n501), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n524), .A2(G43), .ZN(new_n562));
  AND3_X1   g137(.A1(new_n559), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT78), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  AND2_X1   g144(.A1(new_n517), .A2(new_n518), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n570), .A2(new_n571), .A3(G53), .A4(G543), .ZN(new_n572));
  INV_X1    g147(.A(G53), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT9), .B1(new_n523), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G65), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n520), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n521), .A2(G91), .B1(new_n578), .B2(G651), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n575), .A2(new_n579), .ZN(G299));
  NAND3_X1  g155(.A1(new_n553), .A2(new_n557), .A3(KEYINPUT79), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(KEYINPUT79), .B1(new_n553), .B2(new_n557), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(G301));
  NAND3_X1  g159(.A1(new_n570), .A2(G87), .A3(new_n506), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AND2_X1   g162(.A1(G49), .A2(G543), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n517), .A2(new_n518), .A3(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT80), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n517), .A2(KEYINPUT80), .A3(new_n518), .A4(new_n588), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n587), .A2(new_n593), .ZN(G288));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT81), .ZN(new_n596));
  INV_X1    g171(.A(G61), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(new_n504), .B2(new_n505), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n500), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n517), .A2(G86), .A3(new_n506), .A4(new_n518), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n517), .A2(G48), .A3(G543), .A4(new_n518), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(G305));
  AOI22_X1  g177(.A1(G85), .A2(new_n521), .B1(new_n524), .B2(G47), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n501), .B2(new_n604), .ZN(G290));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n570), .A2(new_n506), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n521), .A2(KEYINPUT10), .A3(G92), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n520), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n524), .A2(G54), .B1(new_n614), .B2(G651), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n618));
  NAND2_X1  g193(.A1(G171), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n581), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n617), .B1(new_n620), .B2(G868), .ZN(G284));
  AOI21_X1  g196(.A(new_n617), .B1(new_n620), .B2(G868), .ZN(G321));
  INV_X1    g197(.A(G868), .ZN(new_n623));
  NOR2_X1   g198(.A1(G286), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g199(.A1(new_n575), .A2(new_n579), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT82), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n624), .B1(new_n626), .B2(new_n623), .ZN(G297));
  AOI21_X1  g202(.A(new_n624), .B1(new_n626), .B2(new_n623), .ZN(G280));
  INV_X1    g203(.A(new_n616), .ZN(new_n629));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G860), .ZN(G148));
  OAI21_X1  g206(.A(KEYINPUT83), .B1(new_n616), .B2(G559), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT83), .ZN(new_n634));
  NAND4_X1  g209(.A1(new_n611), .A2(new_n634), .A3(new_n630), .A4(new_n615), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  NOR3_X1   g211(.A1(new_n633), .A2(new_n623), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n623), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n477), .A2(new_n466), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT84), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(G2100), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT85), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n479), .A2(G123), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n464), .A2(G135), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n465), .A2(G111), .ZN(new_n648));
  OAI21_X1  g223(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n646), .B(new_n647), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(G2096), .Z(new_n651));
  OAI211_X1 g226(.A(new_n645), .B(new_n651), .C1(G2100), .C2(new_n643), .ZN(G156));
  INV_X1    g227(.A(KEYINPUT14), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n655), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n658), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(G14), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(G401));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT86), .Z(new_n671));
  NOR2_X1   g246(.A1(G2072), .A2(G2078), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n442), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n669), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(KEYINPUT17), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n674), .B1(new_n671), .B2(new_n675), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n669), .B(new_n670), .C1(new_n442), .C2(new_n672), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT18), .Z(new_n678));
  NAND3_X1  g253(.A1(new_n671), .A2(new_n675), .A3(new_n669), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n676), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2096), .B(G2100), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G227));
  XOR2_X1   g258(.A(G1971), .B(G1976), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n686), .A2(new_n687), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  MUX2_X1   g268(.A(new_n693), .B(new_n692), .S(new_n685), .Z(new_n694));
  NOR2_X1   g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(G229));
  NOR2_X1   g276(.A1(G29), .A2(G32), .ZN(new_n702));
  AOI22_X1  g277(.A1(new_n479), .A2(G129), .B1(new_n464), .B2(G141), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT92), .B(KEYINPUT26), .ZN(new_n704));
  AND3_X1   g279(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n706), .A2(new_n707), .B1(G105), .B2(new_n466), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT93), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n702), .B1(new_n710), .B2(G29), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT27), .B(G1996), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G26), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  INV_X1    g291(.A(G128), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n465), .ZN(new_n718));
  INV_X1    g293(.A(G140), .ZN(new_n719));
  OAI22_X1  g294(.A1(new_n717), .A2(new_n478), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(G2104), .B1(new_n465), .B2(G116), .ZN(new_n721));
  OR3_X1    g296(.A1(KEYINPUT90), .A2(G104), .A3(G2105), .ZN(new_n722));
  OAI21_X1  g297(.A(KEYINPUT90), .B1(G104), .B2(G2105), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n716), .B1(new_n725), .B2(new_n714), .ZN(new_n726));
  INV_X1    g301(.A(G2067), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT30), .B(G28), .ZN(new_n729));
  OR2_X1    g304(.A1(KEYINPUT31), .A2(G11), .ZN(new_n730));
  NAND2_X1  g305(.A1(KEYINPUT31), .A2(G11), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n729), .A2(new_n714), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G29), .A2(G35), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G162), .B2(G29), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT29), .B(G2090), .ZN(new_n735));
  OAI221_X1 g310(.A(new_n732), .B1(new_n714), .B2(new_n650), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  NOR3_X1   g311(.A1(KEYINPUT91), .A2(G29), .A3(G33), .ZN(new_n737));
  OAI21_X1  g312(.A(KEYINPUT91), .B1(G29), .B2(G33), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(new_n465), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT25), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n464), .A2(G139), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n741), .A2(new_n746), .ZN(new_n747));
  AOI211_X1 g322(.A(new_n737), .B(new_n739), .C1(new_n747), .C2(G29), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(G2072), .ZN(new_n749));
  NOR2_X1   g324(.A1(G164), .A2(new_n714), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G27), .B2(new_n714), .ZN(new_n751));
  INV_X1    g326(.A(G2078), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR3_X1   g328(.A1(new_n736), .A2(new_n749), .A3(new_n753), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n713), .A2(new_n728), .A3(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G16), .A2(G19), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n563), .B2(G16), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n757), .A2(G1341), .ZN(new_n758));
  INV_X1    g333(.A(G1966), .ZN(new_n759));
  NAND2_X1  g334(.A1(G168), .A2(G16), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G16), .B2(G21), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n758), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n748), .A2(G2072), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n734), .A2(new_n735), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n763), .B(new_n764), .C1(new_n751), .C2(new_n752), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n762), .B(new_n766), .C1(new_n759), .C2(new_n761), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n755), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G16), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G5), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G171), .B2(new_n769), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n768), .B1(G1961), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(G1961), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT94), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n769), .A2(G4), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n629), .B2(new_n769), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT89), .B(G1348), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n769), .A2(G20), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT23), .Z(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G299), .B2(G16), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT95), .B(G1956), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n714), .B1(KEYINPUT24), .B2(G34), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(KEYINPUT24), .B2(G34), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n475), .B2(G29), .ZN(new_n786));
  INV_X1    g361(.A(G2084), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G1341), .B2(new_n757), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n778), .A2(new_n783), .A3(new_n789), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n772), .A2(new_n774), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(G303), .A2(G16), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n769), .A2(G22), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n794), .A2(KEYINPUT88), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(KEYINPUT88), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(G1971), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n795), .A2(G1971), .A3(new_n796), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  MUX2_X1   g376(.A(G6), .B(G305), .S(G16), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT32), .ZN(new_n803));
  INV_X1    g378(.A(G1981), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n769), .A2(G23), .ZN(new_n806));
  INV_X1    g381(.A(G288), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(new_n769), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT33), .B(G1976), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n805), .A2(new_n810), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n801), .A2(new_n811), .A3(KEYINPUT34), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n769), .A2(G24), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G290), .B2(G16), .ZN(new_n814));
  INV_X1    g389(.A(G1986), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n479), .A2(G119), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n464), .A2(G131), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n465), .A2(G107), .ZN(new_n819));
  OAI21_X1  g394(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n817), .B(new_n818), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  MUX2_X1   g396(.A(G25), .B(new_n821), .S(G29), .Z(new_n822));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G1991), .Z(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n822), .B(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n814), .A2(new_n815), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n816), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n812), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT36), .ZN(new_n830));
  OAI21_X1  g405(.A(KEYINPUT34), .B1(new_n801), .B2(new_n811), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n830), .B1(new_n829), .B2(new_n831), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n791), .B1(new_n833), .B2(new_n834), .ZN(G150));
  INV_X1    g410(.A(G150), .ZN(G311));
  AOI22_X1  g411(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(new_n501), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT97), .B(G55), .Z(new_n839));
  INV_X1    g414(.A(G93), .ZN(new_n840));
  OAI221_X1 g415(.A(new_n838), .B1(new_n523), .B2(new_n839), .C1(new_n607), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(G860), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT37), .Z(new_n843));
  NOR2_X1   g418(.A1(new_n616), .A2(new_n630), .ZN(new_n844));
  XNOR2_X1  g419(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n841), .B1(new_n563), .B2(KEYINPUT98), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n559), .A2(new_n562), .A3(new_n561), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT98), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n841), .A2(new_n849), .A3(new_n848), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n846), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n856));
  INV_X1    g431(.A(G860), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n855), .B2(KEYINPUT39), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n843), .B1(new_n856), .B2(new_n858), .ZN(G145));
  NAND2_X1  g434(.A1(new_n479), .A2(G130), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n465), .A2(G118), .ZN(new_n861));
  OAI21_X1  g436(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(G142), .B2(new_n464), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n641), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n821), .ZN(new_n866));
  OAI21_X1  g441(.A(G164), .B1(new_n724), .B2(new_n720), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n725), .A2(new_n496), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT99), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n710), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n710), .B1(new_n871), .B2(new_n873), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n747), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n870), .A2(new_n709), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n870), .A2(new_n709), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n878), .A2(new_n879), .A3(new_n747), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n866), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n650), .B(new_n475), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n484), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n877), .A2(new_n881), .A3(new_n866), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n883), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(G37), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT100), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n887), .B1(new_n882), .B2(new_n891), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n877), .A2(KEYINPUT100), .A3(new_n881), .A4(new_n866), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n886), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT40), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(G395));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n616), .A2(G299), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n625), .A2(new_n611), .A3(new_n615), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  AND4_X1   g477(.A1(new_n632), .A2(new_n851), .A3(new_n635), .A4(new_n852), .ZN(new_n903));
  AOI22_X1  g478(.A1(new_n852), .A2(new_n851), .B1(new_n632), .B2(new_n635), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n903), .A2(new_n904), .ZN(new_n908));
  OR3_X1    g483(.A1(new_n901), .A2(KEYINPUT102), .A3(KEYINPUT41), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n616), .A2(G299), .ZN(new_n910));
  AOI22_X1  g485(.A1(new_n611), .A2(new_n615), .B1(new_n575), .B2(new_n579), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT41), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n899), .A2(new_n900), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(KEYINPUT102), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n908), .A2(new_n909), .A3(new_n915), .ZN(new_n916));
  OAI211_X1 g491(.A(KEYINPUT101), .B(new_n902), .C1(new_n903), .C2(new_n904), .ZN(new_n917));
  AND4_X1   g492(.A1(new_n898), .A2(new_n907), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  INV_X1    g494(.A(new_n907), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT103), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  XOR2_X1   g496(.A(G290), .B(G305), .Z(new_n922));
  XNOR2_X1  g497(.A(G166), .B(G288), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT42), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n924), .A2(KEYINPUT42), .A3(new_n925), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n918), .B1(new_n921), .B2(new_n931), .ZN(new_n932));
  NOR4_X1   g507(.A1(new_n930), .A2(new_n919), .A3(new_n920), .A4(KEYINPUT103), .ZN(new_n933));
  OAI21_X1  g508(.A(G868), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n841), .A2(new_n623), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(G295));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n935), .ZN(G331));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n620), .A2(G168), .ZN(new_n939));
  NOR2_X1   g514(.A1(G171), .A2(G168), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n939), .A2(new_n853), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n853), .B1(new_n939), .B2(new_n941), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n902), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(G286), .B1(new_n619), .B2(new_n581), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n852), .B(new_n851), .C1(new_n945), .C2(new_n940), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n939), .A2(new_n853), .A3(new_n941), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n909), .A2(new_n946), .A3(new_n947), .A4(new_n915), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n944), .A2(new_n948), .A3(new_n926), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n889), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n926), .B1(new_n944), .B2(new_n948), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n938), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT104), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n914), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n899), .A2(new_n900), .A3(KEYINPUT104), .A4(new_n913), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(new_n912), .A3(new_n955), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n956), .A2(new_n946), .A3(new_n947), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n901), .B1(new_n947), .B2(new_n946), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n924), .B(new_n925), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n959), .A2(KEYINPUT43), .A3(new_n889), .A4(new_n949), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n952), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT44), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT43), .B1(new_n950), .B2(new_n951), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n959), .A2(new_n938), .A3(new_n889), .A4(new_n949), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n962), .A2(new_n967), .ZN(G397));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n969));
  INV_X1    g544(.A(G8), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n467), .B(G40), .C1(new_n474), .C2(new_n465), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n496), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n972), .A2(KEYINPUT118), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT118), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT45), .B1(new_n496), .B2(new_n973), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n978), .B1(new_n971), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n973), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n977), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n974), .A2(KEYINPUT50), .ZN(new_n983));
  XNOR2_X1  g558(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n496), .A2(new_n973), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n972), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n982), .A2(new_n759), .B1(new_n987), .B2(new_n787), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n970), .B1(new_n988), .B2(G168), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n982), .A2(new_n759), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n787), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(G286), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n969), .B1(new_n989), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n990), .A2(G168), .A3(new_n991), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(G8), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(KEYINPUT51), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT62), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n988), .A2(G168), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT51), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT62), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n989), .A2(new_n969), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT108), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n971), .B1(new_n1004), .B2(new_n979), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT105), .B(G1384), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT109), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n496), .A2(new_n1009), .A3(KEYINPUT45), .A4(new_n1006), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n976), .A2(KEYINPUT108), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1005), .A2(new_n1011), .A3(new_n752), .A4(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(G2078), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n977), .A2(new_n980), .A3(new_n981), .A4(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1961), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n986), .A2(new_n1018), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n1017), .A2(new_n1019), .A3(KEYINPUT121), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT121), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1015), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1022), .A2(new_n620), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n979), .A2(new_n1004), .ZN(new_n1025));
  AOI211_X1 g600(.A(KEYINPUT108), .B(KEYINPUT45), .C1(new_n496), .C2(new_n973), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n1025), .A2(new_n1026), .A3(new_n971), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1971), .B1(new_n1027), .B2(new_n1011), .ZN(new_n1028));
  XOR2_X1   g603(.A(KEYINPUT111), .B(G2090), .Z(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n986), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1024), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT114), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G303), .A2(G8), .ZN(new_n1035));
  NAND2_X1  g610(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1036), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1034), .ZN(new_n1039));
  AOI211_X1 g614(.A(new_n1038), .B(new_n1039), .C1(G303), .C2(G8), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1005), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n798), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1031), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(new_n1044), .A3(KEYINPUT112), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1032), .A2(new_n1041), .A3(G8), .A4(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1041), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT117), .B1(new_n974), .B2(KEYINPUT50), .ZN(new_n1048));
  INV_X1    g623(.A(new_n984), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n974), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT50), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n496), .A2(new_n1051), .A3(new_n1052), .A4(new_n973), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1048), .A2(new_n972), .A3(new_n1050), .A4(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(new_n1030), .ZN(new_n1055));
  OAI21_X1  g630(.A(G8), .B1(new_n1028), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1047), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(G8), .B1(new_n971), .B2(new_n974), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  OAI211_X1 g635(.A(KEYINPUT115), .B(G8), .C1(new_n971), .C2(new_n974), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G1976), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT52), .B1(G288), .B2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n587), .A2(KEYINPUT116), .A3(G1976), .A4(new_n593), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n593), .A2(G1976), .A3(new_n586), .A4(new_n585), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1062), .A2(new_n1064), .A3(new_n1069), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1061), .ZN(new_n1072));
  NAND2_X1  g647(.A1(G305), .A2(G1981), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT49), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n599), .A2(new_n600), .A3(new_n601), .A4(new_n804), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1074), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1077));
  OAI22_X1  g652(.A1(new_n1071), .A2(new_n1072), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1070), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1080), .B1(new_n1062), .B2(new_n1069), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1046), .A2(new_n1057), .A3(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n998), .A2(new_n1003), .A3(new_n1023), .A4(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT125), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1046), .A2(new_n1057), .A3(new_n1082), .ZN(new_n1087));
  INV_X1    g662(.A(G1996), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1005), .A2(new_n1011), .A3(new_n1088), .A4(new_n1012), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT58), .B(G1341), .Z(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n971), .B2(new_n974), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n563), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1094), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1092), .A2(new_n563), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT61), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n575), .A2(new_n579), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1100), .B1(new_n575), .B2(new_n579), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT119), .B(G1956), .Z(new_n1104));
  NAND2_X1  g679(.A1(new_n1054), .A2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT56), .B(G2072), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1005), .A2(new_n1011), .A3(new_n1012), .A4(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1103), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1099), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n986), .A2(new_n777), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n972), .A2(new_n973), .A3(new_n727), .A4(new_n496), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(KEYINPUT60), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT60), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1114), .B1(new_n1115), .B2(new_n616), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1117), .A2(KEYINPUT60), .A3(new_n629), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1103), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1122), .A2(KEYINPUT61), .A3(new_n1108), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1098), .A2(new_n1111), .A3(new_n1119), .A4(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1117), .A2(new_n616), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1110), .B1(new_n1125), .B2(new_n1108), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1087), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1016), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n496), .A2(new_n1006), .ZN(new_n1130));
  OR2_X1    g705(.A1(new_n1130), .A2(KEYINPUT106), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT45), .B1(new_n1130), .B2(KEYINPUT106), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1129), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n467), .A2(G40), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n474), .A2(KEYINPUT122), .ZN(new_n1135));
  OAI21_X1  g710(.A(G2105), .B1(new_n474), .B2(KEYINPUT122), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT123), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1139), .B(new_n1134), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1133), .A2(new_n1138), .A3(new_n1011), .A4(new_n1140), .ZN(new_n1141));
  AND4_X1   g716(.A1(G301), .A2(new_n1015), .A3(new_n1019), .A4(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(KEYINPUT124), .B(new_n1128), .C1(new_n1023), .C2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1142), .B1(new_n1022), .B2(new_n620), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1144), .B1(new_n1145), .B2(KEYINPUT54), .ZN(new_n1146));
  OAI211_X1 g721(.A(G301), .B(new_n1015), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1015), .A2(new_n1141), .A3(new_n1019), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1128), .B1(new_n1148), .B2(G171), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1000), .A2(new_n1002), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1127), .A2(new_n1143), .A3(new_n1146), .A4(new_n1150), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1078), .A2(new_n1063), .A3(new_n807), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1075), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1062), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1082), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1154), .B1(new_n1155), .B2(new_n1046), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n992), .A2(G8), .A3(G168), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1157), .B1(new_n1087), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1032), .A2(G8), .A3(new_n1045), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n1047), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1158), .A2(new_n1157), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1161), .A2(new_n1162), .A3(new_n1046), .A4(new_n1082), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1156), .B1(new_n1159), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1022), .A2(new_n620), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1087), .A2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1166), .A2(KEYINPUT125), .A3(new_n998), .A4(new_n1003), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1086), .A2(new_n1151), .A3(new_n1164), .A4(new_n1167), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n972), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1170), .A2(new_n1088), .A3(new_n709), .ZN(new_n1171));
  XOR2_X1   g746(.A(new_n1171), .B(KEYINPUT107), .Z(new_n1172));
  INV_X1    g747(.A(new_n1170), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n725), .B(G2067), .ZN(new_n1174));
  INV_X1    g749(.A(new_n710), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1174), .B1(new_n1175), .B2(G1996), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1172), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n821), .A2(new_n824), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n821), .A2(new_n824), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1173), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(G290), .B(G1986), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1181), .B1(new_n1173), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1168), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1170), .B1(new_n709), .B2(new_n1174), .ZN(new_n1185));
  OR3_X1    g760(.A1(new_n1170), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1186));
  OAI21_X1  g761(.A(KEYINPUT46), .B1(new_n1170), .B2(G1996), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1185), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  XOR2_X1   g763(.A(new_n1188), .B(KEYINPUT47), .Z(new_n1189));
  NOR3_X1   g764(.A1(new_n1170), .A2(G1986), .A3(G290), .ZN(new_n1190));
  XOR2_X1   g765(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1191));
  XNOR2_X1  g766(.A(new_n1190), .B(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1189), .B1(new_n1181), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n725), .A2(new_n727), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1170), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1184), .A2(new_n1197), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g773(.A(G319), .B(new_n682), .C1(new_n666), .C2(new_n667), .ZN(new_n1200));
  NOR2_X1   g774(.A1(G229), .A2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g775(.A(new_n1201), .B1(new_n894), .B2(new_n890), .ZN(new_n1202));
  AOI21_X1  g776(.A(new_n1202), .B1(new_n963), .B2(new_n964), .ZN(G308));
  OAI211_X1 g777(.A(new_n965), .B(new_n1201), .C1(new_n894), .C2(new_n890), .ZN(G225));
endmodule


