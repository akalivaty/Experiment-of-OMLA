//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n213), .A2(KEYINPUT0), .ZN(new_n214));
  OR2_X1    g0014(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n215), .A2(G50), .A3(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n208), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n213), .A2(KEYINPUT0), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n214), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT65), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n210), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n224), .A2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT66), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  AND2_X1   g0051(.A1(new_n251), .A2(new_n219), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n252), .B(new_n253), .C1(G1), .C2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT81), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT25), .ZN(new_n258));
  INV_X1    g0058(.A(G107), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(new_n257), .B2(KEYINPUT25), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n258), .B1(new_n260), .B2(new_n253), .ZN(new_n261));
  INV_X1    g0061(.A(new_n253), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n262), .A2(new_n257), .A3(KEYINPUT25), .A4(new_n259), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n256), .A2(G107), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT24), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n208), .B(G87), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT22), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT22), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n270), .A2(new_n271), .A3(new_n208), .A4(G87), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G116), .ZN(new_n274));
  NOR3_X1   g0074(.A1(new_n254), .A2(new_n274), .A3(G20), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT23), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n276), .B1(new_n208), .B2(G107), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n259), .A2(KEYINPUT23), .A3(G20), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n265), .B1(new_n273), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n273), .A2(new_n265), .A3(new_n279), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n251), .A2(new_n219), .ZN(new_n284));
  AOI21_X1  g0084(.A(KEYINPUT80), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n282), .ZN(new_n286));
  OAI211_X1 g0086(.A(KEYINPUT80), .B(new_n284), .C1(new_n286), .C2(new_n280), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n264), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT5), .B(G41), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G1), .A3(G13), .ZN(new_n292));
  AND3_X1   g0092(.A1(new_n207), .A2(G45), .A3(G274), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G45), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(G1), .ZN(new_n297));
  AND2_X1   g0097(.A1(KEYINPUT5), .A2(G41), .ZN(new_n298));
  NOR2_X1   g0098(.A1(KEYINPUT5), .A2(G41), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n300), .A2(G264), .A3(new_n292), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT84), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT84), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n300), .A2(new_n303), .A3(G264), .A4(new_n292), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n295), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  OAI211_X1 g0105(.A(G257), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT82), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT82), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n270), .A2(new_n308), .A3(G257), .A4(G1698), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G294), .ZN(new_n310));
  INV_X1    g0110(.A(G1698), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n270), .A2(G250), .A3(new_n311), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n307), .A2(new_n309), .A3(new_n310), .A4(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n305), .B1(new_n315), .B2(KEYINPUT83), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT83), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(new_n313), .B2(new_n314), .ZN(new_n318));
  OAI21_X1  g0118(.A(G169), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n302), .A2(new_n304), .ZN(new_n320));
  AND3_X1   g0120(.A1(new_n315), .A2(KEYINPUT85), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT85), .B1(new_n315), .B2(new_n320), .ZN(new_n322));
  OAI211_X1 g0122(.A(G179), .B(new_n294), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT86), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n319), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n315), .A2(new_n320), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT85), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n315), .A2(KEYINPUT85), .A3(new_n320), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n295), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(KEYINPUT86), .B1(new_n330), .B2(G179), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n289), .B1(new_n325), .B2(new_n331), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n311), .A2(G226), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n270), .B(new_n333), .C1(G223), .C2(G1698), .ZN(new_n334));
  NAND2_X1  g0134(.A1(G33), .A2(G87), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n292), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n207), .B(G274), .C1(G41), .C2(G45), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n292), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n337), .B1(new_n339), .B2(new_n235), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G179), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(G169), .B2(new_n341), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT72), .ZN(new_n345));
  AND2_X1   g0145(.A1(KEYINPUT68), .A2(G58), .ZN(new_n346));
  NOR2_X1   g0146(.A1(KEYINPUT68), .A2(G58), .ZN(new_n347));
  OAI21_X1  g0147(.A(G68), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n208), .B1(new_n348), .B2(new_n202), .ZN(new_n349));
  NOR2_X1   g0149(.A1(G20), .A2(G33), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G159), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n345), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n353), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT68), .B(G58), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n201), .B1(new_n356), .B2(G68), .ZN(new_n357));
  OAI211_X1 g0157(.A(KEYINPUT72), .B(new_n355), .C1(new_n357), .C2(new_n208), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n266), .A2(new_n267), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT7), .B1(new_n359), .B2(new_n208), .ZN(new_n360));
  OR2_X1    g0160(.A1(KEYINPUT3), .A2(G33), .ZN(new_n361));
  NAND2_X1  g0161(.A1(KEYINPUT3), .A2(G33), .ZN(new_n362));
  AND4_X1   g0162(.A1(KEYINPUT7), .A2(new_n361), .A3(new_n208), .A4(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(G68), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n354), .A2(new_n358), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT16), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n252), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n354), .A2(new_n358), .A3(new_n364), .A4(KEYINPUT16), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(KEYINPUT8), .A2(G58), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(new_n356), .B2(KEYINPUT8), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n207), .A2(G20), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(KEYINPUT73), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n252), .A2(new_n253), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT73), .B1(new_n371), .B2(new_n372), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n376), .A2(new_n377), .B1(new_n253), .B2(new_n371), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n344), .B1(new_n369), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT18), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G200), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n341), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G190), .ZN(new_n385));
  NOR3_X1   g0185(.A1(new_n336), .A2(new_n385), .A3(new_n340), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n369), .A2(new_n379), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT17), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n378), .B1(new_n367), .B2(new_n368), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT18), .B1(new_n391), .B2(new_n344), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(KEYINPUT17), .A3(new_n387), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n382), .A2(new_n390), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n337), .ZN(new_n396));
  INV_X1    g0196(.A(new_n339), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n396), .B1(new_n397), .B2(G226), .ZN(new_n398));
  AOI21_X1  g0198(.A(G1698), .B1(new_n361), .B2(new_n362), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G222), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n400), .B(KEYINPUT67), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n359), .A2(new_n311), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n402), .A2(G223), .B1(G77), .B2(new_n359), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n398), .B1(new_n404), .B2(new_n292), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G200), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n372), .A2(G50), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G50), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n375), .A2(new_n408), .B1(new_n409), .B2(new_n262), .ZN(new_n410));
  OAI21_X1  g0210(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n411));
  INV_X1    g0211(.A(G150), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n411), .B1(new_n412), .B2(new_n351), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n208), .A2(G33), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n413), .B1(new_n415), .B2(new_n371), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n410), .B1(new_n416), .B2(new_n252), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT9), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n406), .B(new_n418), .C1(new_n405), .C2(new_n385), .ZN(new_n419));
  XNOR2_X1  g0219(.A(new_n419), .B(KEYINPUT10), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n405), .A2(G179), .ZN(new_n421));
  INV_X1    g0221(.A(G169), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n405), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(new_n417), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n235), .A2(G1698), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(G226), .B2(G1698), .ZN(new_n428));
  INV_X1    g0228(.A(G97), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n428), .A2(new_n359), .B1(new_n254), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n314), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n292), .A2(G238), .A3(new_n338), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n432), .A2(KEYINPUT70), .A3(new_n337), .ZN(new_n433));
  AOI21_X1  g0233(.A(KEYINPUT70), .B1(new_n432), .B2(new_n337), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT13), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT13), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n431), .B(new_n437), .C1(new_n433), .C2(new_n434), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G169), .ZN(new_n440));
  INV_X1    g0240(.A(new_n439), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n440), .A2(KEYINPUT14), .B1(new_n441), .B2(G179), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n422), .B1(new_n436), .B2(new_n438), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT14), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(KEYINPUT71), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT71), .B1(new_n443), .B2(new_n444), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n442), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G68), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n350), .A2(G50), .B1(G20), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G77), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(new_n414), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT11), .B1(new_n452), .B2(new_n284), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n262), .A2(new_n449), .ZN(new_n454));
  XNOR2_X1  g0254(.A(new_n454), .B(KEYINPUT12), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n452), .A2(KEYINPUT11), .A3(new_n284), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n375), .A2(G68), .A3(new_n372), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n448), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n439), .A2(G200), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n458), .A2(new_n453), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n460), .B(new_n461), .C1(new_n385), .C2(new_n439), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  XOR2_X1   g0263(.A(KEYINPUT8), .B(G58), .Z(new_n464));
  AOI22_X1  g0264(.A1(new_n464), .A2(new_n350), .B1(G20), .B2(G77), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT15), .B(G87), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n465), .B1(new_n414), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n284), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n262), .A2(new_n451), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n372), .A2(G77), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n468), .B(new_n469), .C1(new_n374), .C2(new_n470), .ZN(new_n471));
  XNOR2_X1  g0271(.A(new_n471), .B(KEYINPUT69), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n397), .A2(G244), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n402), .A2(G238), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n399), .A2(G232), .B1(new_n359), .B2(G107), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI211_X1 g0276(.A(new_n396), .B(new_n473), .C1(new_n476), .C2(new_n314), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G190), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n472), .B(new_n478), .C1(new_n383), .C2(new_n477), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n471), .B1(new_n477), .B2(G169), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n477), .A2(new_n342), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  AND4_X1   g0284(.A1(new_n395), .A2(new_n426), .A3(new_n463), .A4(new_n484), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n316), .A2(G190), .A3(new_n318), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n294), .B1(new_n321), .B2(new_n322), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n486), .B1(new_n487), .B2(new_n383), .ZN(new_n488));
  OR2_X1    g0288(.A1(new_n488), .A2(new_n289), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n262), .A2(new_n274), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(new_n255), .B2(new_n274), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G33), .A2(G283), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n492), .B(new_n208), .C1(G33), .C2(new_n429), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n493), .B(new_n284), .C1(new_n208), .C2(G116), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT20), .ZN(new_n495));
  OR2_X1    g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n495), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n491), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n314), .B1(new_n297), .B2(new_n290), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n295), .B1(G270), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n270), .A2(G257), .A3(new_n311), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n359), .A2(G303), .ZN(new_n503));
  OAI211_X1 g0303(.A(G264), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n314), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n499), .A2(G169), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT21), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n507), .A2(G200), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n511), .B(new_n498), .C1(new_n385), .C2(new_n507), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT79), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n505), .A2(new_n314), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n500), .A2(G270), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n294), .ZN(new_n516));
  OAI211_X1 g0316(.A(KEYINPUT21), .B(G169), .C1(new_n514), .C2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n501), .A2(G179), .A3(new_n506), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n513), .B1(new_n519), .B2(new_n499), .ZN(new_n520));
  AOI211_X1 g0320(.A(KEYINPUT79), .B(new_n498), .C1(new_n517), .C2(new_n518), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n510), .B(new_n512), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n402), .A2(G244), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n399), .A2(G238), .B1(G33), .B2(G116), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n292), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT77), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n207), .A2(G45), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G250), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n526), .B1(new_n314), .B2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n292), .A2(KEYINPUT77), .A3(G250), .A4(new_n527), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT76), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n293), .A2(new_n531), .A3(new_n292), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n531), .B1(new_n293), .B2(new_n292), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n529), .B(new_n530), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT78), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n207), .A2(G45), .A3(G274), .ZN(new_n536));
  OAI21_X1  g0336(.A(KEYINPUT76), .B1(new_n314), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n293), .A2(new_n292), .A3(new_n531), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT78), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n539), .A2(new_n540), .A3(new_n529), .A4(new_n530), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n525), .B1(new_n535), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G190), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n270), .A2(new_n208), .A3(G68), .ZN(new_n544));
  NAND3_X1  g0344(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n208), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n205), .B2(G87), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT19), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n414), .B2(new_n429), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n544), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(new_n284), .B1(new_n262), .B2(new_n466), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n256), .A2(G87), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n543), .B(new_n553), .C1(new_n383), .C2(new_n542), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n535), .A2(new_n541), .ZN(new_n555));
  INV_X1    g0355(.A(new_n525), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n342), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n551), .B1(new_n255), .B2(new_n466), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n557), .B(new_n558), .C1(G169), .C2(new_n542), .ZN(new_n559));
  OAI211_X1 g0359(.A(G250), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n560));
  OAI211_X1 g0360(.A(G244), .B(new_n311), .C1(new_n266), .C2(new_n267), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT4), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n492), .B(new_n560), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT4), .B1(new_n399), .B2(G244), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n314), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n300), .A2(G257), .A3(new_n292), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n294), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n568), .A3(new_n342), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n561), .A2(new_n562), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n270), .A2(KEYINPUT4), .A3(G244), .A4(new_n311), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n570), .A2(new_n571), .A3(new_n492), .A4(new_n560), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n567), .B1(new_n572), .B2(new_n314), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n569), .B1(G169), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n262), .A2(new_n429), .ZN(new_n575));
  OR2_X1    g0375(.A1(new_n575), .A2(KEYINPUT75), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(KEYINPUT75), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n576), .B(new_n577), .C1(new_n429), .C2(new_n255), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n351), .A2(new_n451), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  XNOR2_X1  g0380(.A(G97), .B(G107), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT6), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n582), .A2(new_n429), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n581), .A2(new_n582), .B1(new_n259), .B2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(KEYINPUT74), .B(new_n580), .C1(new_n584), .C2(new_n208), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT74), .ZN(new_n586));
  AND2_X1   g0386(.A1(G97), .A2(G107), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n582), .B1(new_n587), .B2(new_n204), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n259), .A2(KEYINPUT6), .A3(G97), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n208), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n586), .B1(new_n590), .B2(new_n579), .ZN(new_n591));
  OAI21_X1  g0391(.A(G107), .B1(new_n360), .B2(new_n363), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n585), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n578), .B1(new_n593), .B2(new_n284), .ZN(new_n594));
  OR2_X1    g0394(.A1(new_n574), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n565), .A2(new_n568), .A3(G190), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n594), .B(new_n596), .C1(new_n383), .C2(new_n573), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n554), .A2(new_n559), .A3(new_n595), .A4(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n522), .A2(new_n598), .ZN(new_n599));
  AND4_X1   g0399(.A1(new_n332), .A2(new_n485), .A3(new_n489), .A4(new_n599), .ZN(G372));
  NAND2_X1  g0400(.A1(new_n519), .A2(new_n499), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n510), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n330), .A2(KEYINPUT86), .A3(G179), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n323), .A2(new_n324), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n604), .A3(new_n319), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n602), .B1(new_n605), .B2(new_n289), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n553), .B1(new_n542), .B2(new_n383), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(KEYINPUT87), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT87), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n553), .B(new_n609), .C1(new_n542), .C2(new_n383), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n543), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n559), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n593), .A2(new_n284), .ZN(new_n613));
  INV_X1    g0413(.A(new_n578), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n596), .B1(new_n383), .B2(new_n573), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n574), .A2(new_n594), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n488), .B2(new_n289), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n606), .A2(new_n612), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n557), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n558), .B1(new_n542), .B2(G169), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n607), .A2(KEYINPUT87), .B1(G190), .B2(new_n542), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n624), .B1(new_n625), .B2(new_n610), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n627), .A3(new_n618), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n554), .A2(new_n559), .A3(new_n618), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n624), .B1(new_n629), .B2(KEYINPUT26), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n485), .B1(new_n621), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n424), .ZN(new_n633));
  INV_X1    g0433(.A(new_n459), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n634), .B1(new_n462), .B2(new_n482), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n390), .A2(new_n393), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n392), .B(new_n382), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n633), .B1(new_n637), .B2(new_n420), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n639), .B(KEYINPUT88), .ZN(G369));
  NAND3_X1  g0440(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(G213), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(G343), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n332), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n646), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n284), .B1(new_n286), .B2(new_n280), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT80), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n287), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n648), .B1(new_n652), .B2(new_n264), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n332), .A2(new_n489), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT90), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n605), .A2(new_n656), .A3(new_n653), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n656), .B1(new_n605), .B2(new_n653), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n655), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n510), .B1(new_n520), .B2(new_n521), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(new_n646), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n647), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n498), .A2(new_n648), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n602), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n522), .B2(new_n665), .ZN(new_n667));
  XNOR2_X1  g0467(.A(KEYINPUT89), .B(G330), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n660), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n664), .A2(new_n671), .ZN(G399));
  INV_X1    g0472(.A(new_n211), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(G41), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G1), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n217), .B2(new_n675), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT28), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT30), .ZN(new_n680));
  INV_X1    g0480(.A(new_n518), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n681), .B(new_n542), .C1(new_n321), .C2(new_n322), .ZN(new_n682));
  INV_X1    g0482(.A(new_n573), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n680), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n683), .A2(new_n507), .A3(new_n342), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT91), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n542), .A2(new_n686), .ZN(new_n687));
  AOI211_X1 g0487(.A(KEYINPUT91), .B(new_n525), .C1(new_n535), .C2(new_n541), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n487), .B(new_n685), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n328), .A2(new_n329), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n683), .A2(new_n680), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n690), .A2(new_n681), .A3(new_n542), .A4(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n684), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n693), .A2(KEYINPUT31), .A3(new_n646), .ZN(new_n694));
  AOI21_X1  g0494(.A(KEYINPUT31), .B1(new_n693), .B2(new_n646), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT92), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n693), .A2(new_n646), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT31), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT92), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n693), .A2(KEYINPUT31), .A3(new_n646), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n599), .A2(new_n332), .A3(new_n489), .A4(new_n648), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n696), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n668), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT29), .ZN(new_n706));
  OAI211_X1 g0506(.A(new_n706), .B(new_n648), .C1(new_n621), .C2(new_n631), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n620), .A2(new_n612), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n332), .A2(new_n662), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n624), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n626), .A2(KEYINPUT93), .A3(KEYINPUT26), .A4(new_n618), .ZN(new_n711));
  AND4_X1   g0511(.A1(KEYINPUT26), .A2(new_n611), .A3(new_n559), .A4(new_n618), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT93), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n713), .B1(new_n629), .B2(new_n627), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n711), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n646), .B1(new_n710), .B2(new_n715), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n705), .B(new_n707), .C1(new_n706), .C2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n679), .B1(new_n718), .B2(G1), .ZN(G364));
  AND2_X1   g0519(.A1(new_n208), .A2(G13), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n207), .B1(new_n720), .B2(G45), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n675), .A2(KEYINPUT94), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT94), .ZN(new_n723));
  INV_X1    g0523(.A(new_n721), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n674), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n211), .A2(new_n270), .ZN(new_n728));
  INV_X1    g0528(.A(G355), .ZN(new_n729));
  OAI22_X1  g0529(.A1(new_n728), .A2(new_n729), .B1(G116), .B2(new_n211), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n211), .A2(new_n359), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT95), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n296), .B2(new_n218), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n249), .A2(G45), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n730), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G13), .A2(G33), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n219), .B1(G20), .B2(new_n422), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n727), .B1(new_n735), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n208), .A2(new_n342), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(G190), .A3(G200), .ZN(new_n744));
  INV_X1    g0544(.A(new_n356), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n743), .A2(G190), .A3(new_n383), .ZN(new_n746));
  OAI221_X1 g0546(.A(new_n270), .B1(new_n744), .B2(new_n409), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n208), .A2(new_n383), .A3(G179), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n748), .A2(new_n385), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n259), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n748), .A2(G190), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI211_X1 g0553(.A(new_n747), .B(new_n751), .C1(G87), .C2(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n743), .A2(new_n385), .A3(G200), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n342), .A2(new_n383), .A3(G190), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n756), .A2(G68), .B1(G97), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(KEYINPUT97), .B(G159), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G190), .A2(G200), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n761), .A2(G20), .A3(new_n342), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g0563(.A(KEYINPUT98), .B(KEYINPUT32), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n743), .A2(new_n761), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n766), .A2(KEYINPUT96), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(KEYINPUT96), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G77), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n754), .A2(new_n759), .A3(new_n765), .A4(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(KEYINPUT33), .B(G317), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n774), .A2(KEYINPUT99), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n755), .B1(new_n774), .B2(KEYINPUT99), .ZN(new_n776));
  INV_X1    g0576(.A(new_n746), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n775), .A2(new_n776), .B1(G322), .B2(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT100), .ZN(new_n779));
  INV_X1    g0579(.A(G283), .ZN(new_n780));
  INV_X1    g0580(.A(new_n758), .ZN(new_n781));
  INV_X1    g0581(.A(G294), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n750), .A2(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G303), .ZN(new_n784));
  INV_X1    g0584(.A(G326), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n752), .A2(new_n784), .B1(new_n744), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n762), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n270), .B1(new_n788), .B2(G329), .ZN(new_n789));
  INV_X1    g0589(.A(G311), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n787), .B(new_n789), .C1(new_n790), .C2(new_n766), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n772), .B1(new_n779), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n742), .B1(new_n792), .B2(new_n739), .ZN(new_n793));
  INV_X1    g0593(.A(new_n738), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n793), .B1(new_n667), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT101), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n667), .A2(new_n668), .ZN(new_n797));
  AND3_X1   g0597(.A1(new_n797), .A2(new_n669), .A3(new_n726), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(G396));
  OAI21_X1  g0600(.A(new_n648), .B1(new_n621), .B2(new_n631), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n483), .A2(KEYINPUT103), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT103), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n482), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n471), .A2(new_n646), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n479), .A2(new_n806), .ZN(new_n807));
  AND3_X1   g0607(.A1(new_n482), .A2(KEYINPUT104), .A3(new_n646), .ZN(new_n808));
  AOI21_X1  g0608(.A(KEYINPUT104), .B1(new_n482), .B2(new_n646), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n805), .A2(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n801), .B(new_n810), .Z(new_n811));
  AOI21_X1  g0611(.A(new_n727), .B1(new_n811), .B2(new_n705), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n705), .B2(new_n811), .ZN(new_n813));
  INV_X1    g0613(.A(new_n739), .ZN(new_n814));
  INV_X1    g0614(.A(G137), .ZN(new_n815));
  XNOR2_X1  g0615(.A(KEYINPUT102), .B(G143), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n815), .A2(new_n744), .B1(new_n746), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n769), .A2(new_n760), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n817), .B(new_n818), .C1(G150), .C2(new_n756), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n819), .A2(KEYINPUT34), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(KEYINPUT34), .ZN(new_n821));
  INV_X1    g0621(.A(G132), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n270), .B1(new_n822), .B2(new_n762), .C1(new_n781), .C2(new_n745), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n750), .A2(new_n449), .B1(new_n409), .B2(new_n752), .ZN(new_n824));
  OR4_X1    g0624(.A1(new_n820), .A2(new_n821), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n770), .A2(G116), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n749), .A2(G87), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G97), .B2(new_n758), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n752), .A2(new_n259), .B1(new_n755), .B2(new_n780), .ZN(new_n829));
  INV_X1    g0629(.A(new_n744), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n829), .B1(G303), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n359), .B1(new_n762), .B2(new_n790), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(G294), .B2(new_n777), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n826), .A2(new_n828), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n814), .B1(new_n825), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n739), .A2(new_n736), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n726), .B(new_n835), .C1(new_n451), .C2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n810), .B2(new_n737), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n813), .A2(new_n838), .ZN(G384));
  INV_X1    g0639(.A(new_n584), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n840), .A2(KEYINPUT35), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(KEYINPUT35), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n841), .A2(new_n842), .A3(G116), .A4(new_n220), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT36), .Z(new_n844));
  NAND3_X1  g0644(.A1(new_n218), .A2(G77), .A3(new_n348), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n409), .A2(G68), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n207), .B(G13), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT37), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n369), .A2(new_n379), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT106), .ZN(new_n851));
  INV_X1    g0651(.A(new_n644), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT106), .B1(new_n391), .B2(new_n644), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n369), .A2(new_n379), .A3(new_n387), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n856), .A2(new_n380), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n849), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n380), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n850), .A2(new_n852), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n859), .A2(new_n860), .A3(new_n849), .A4(new_n388), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(KEYINPUT107), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT107), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n388), .B1(new_n391), .B2(new_n344), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n854), .B2(new_n853), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n864), .B(new_n861), .C1(new_n866), .C2(new_n849), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n394), .A2(new_n854), .A3(new_n853), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n863), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n863), .A2(new_n867), .A3(KEYINPUT38), .A4(new_n868), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n871), .A2(KEYINPUT39), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n459), .A2(new_n646), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n863), .A2(new_n867), .A3(new_n868), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT108), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n391), .A2(new_n644), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT37), .B1(new_n865), .B2(new_n877), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n861), .A2(new_n878), .B1(new_n394), .B2(new_n877), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n876), .B1(new_n879), .B2(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(new_n861), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n394), .A2(new_n877), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(KEYINPUT108), .A3(new_n870), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n875), .A2(KEYINPUT38), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n873), .B(new_n874), .C1(new_n885), .C2(KEYINPUT39), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n852), .B1(new_n382), .B2(new_n392), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n871), .A2(new_n872), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT105), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n461), .A2(new_n648), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n459), .A2(new_n889), .A3(new_n462), .A4(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n442), .B(new_n462), .C1(new_n446), .C2(new_n447), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n889), .B1(new_n893), .B2(new_n890), .ZN(new_n894));
  OAI22_X1  g0694(.A1(new_n443), .A2(new_n444), .B1(new_n439), .B2(new_n342), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n443), .A2(new_n444), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT71), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n895), .B1(new_n898), .B2(new_n445), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n462), .B(new_n891), .C1(new_n899), .C2(new_n461), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n894), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n892), .A2(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n648), .B(new_n810), .C1(new_n621), .C2(new_n631), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n646), .B1(new_n802), .B2(new_n804), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n902), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n887), .B1(new_n888), .B2(new_n906), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n886), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n707), .B1(new_n716), .B2(new_n706), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n485), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n638), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n908), .B(new_n911), .Z(new_n912));
  NAND3_X1  g0712(.A1(new_n703), .A2(new_n699), .A3(new_n701), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n810), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n914), .A2(new_n902), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT40), .B1(new_n888), .B2(new_n915), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n892), .A2(new_n901), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n917), .A2(KEYINPUT40), .A3(new_n810), .A4(new_n913), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n885), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n485), .A2(new_n913), .ZN(new_n920));
  OR3_X1    g0720(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n920), .B1(new_n916), .B2(new_n919), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(new_n668), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n912), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n207), .B2(new_n720), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n912), .A2(new_n923), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n848), .B1(new_n925), .B2(new_n926), .ZN(G367));
  OAI21_X1  g0727(.A(new_n619), .B1(new_n594), .B2(new_n648), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n618), .A2(new_n646), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n671), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n553), .A2(new_n648), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n624), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n612), .B2(new_n933), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT43), .Z(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT110), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT42), .ZN(new_n939));
  INV_X1    g0739(.A(new_n663), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n653), .B1(new_n325), .B2(new_n331), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT90), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n657), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n940), .B1(new_n943), .B2(new_n655), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n939), .B1(new_n944), .B2(new_n930), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n332), .A2(new_n928), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n646), .B1(new_n946), .B2(new_n595), .ZN(new_n947));
  OAI21_X1  g0747(.A(KEYINPUT109), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n660), .A2(new_n663), .A3(new_n930), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(KEYINPUT42), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT109), .ZN(new_n951));
  INV_X1    g0751(.A(new_n947), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n948), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n949), .A2(KEYINPUT42), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n938), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  AOI211_X1 g0757(.A(KEYINPUT110), .B(new_n955), .C1(new_n948), .C2(new_n953), .ZN(new_n958));
  OAI211_X1 g0758(.A(KEYINPUT111), .B(new_n937), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n951), .B1(new_n950), .B2(new_n952), .ZN(new_n960));
  AOI211_X1 g0760(.A(KEYINPUT109), .B(new_n947), .C1(new_n949), .C2(KEYINPUT42), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT110), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n954), .A2(new_n938), .A3(new_n956), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n963), .A2(KEYINPUT43), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n959), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n963), .A2(new_n964), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n937), .B1(new_n967), .B2(KEYINPUT111), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n932), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n671), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT44), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n664), .B2(new_n930), .ZN(new_n972));
  OAI211_X1 g0772(.A(KEYINPUT44), .B(new_n931), .C1(new_n944), .C2(new_n647), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n664), .A2(new_n930), .ZN(new_n976));
  XOR2_X1   g0776(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n664), .A2(new_n930), .A3(new_n977), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n970), .B1(new_n975), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n943), .A2(new_n655), .A3(new_n940), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n669), .B1(new_n984), .B2(new_n944), .ZN(new_n985));
  INV_X1    g0785(.A(new_n944), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n986), .A2(new_n670), .A3(new_n983), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n717), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n974), .A2(new_n671), .A3(new_n980), .A4(new_n979), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n982), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n718), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n674), .B(KEYINPUT41), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n721), .ZN(new_n995));
  OAI21_X1  g0795(.A(KEYINPUT111), .B1(new_n957), .B2(new_n958), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n936), .ZN(new_n997));
  INV_X1    g0797(.A(new_n932), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n997), .A2(new_n998), .A3(new_n965), .A4(new_n959), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n969), .A2(new_n995), .A3(new_n999), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n732), .A2(new_n241), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n466), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n741), .B1(new_n673), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n726), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n270), .B1(new_n746), .B2(new_n412), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n750), .A2(new_n451), .B1(new_n755), .B2(new_n760), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(G137), .C2(new_n788), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n752), .A2(new_n745), .B1(new_n744), .B2(new_n816), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(G68), .B2(new_n758), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1007), .B(new_n1009), .C1(new_n409), .C2(new_n769), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n753), .A2(G116), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT46), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n750), .A2(new_n429), .B1(new_n755), .B2(new_n782), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n781), .A2(new_n259), .B1(new_n744), .B2(new_n790), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n770), .A2(G283), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n359), .B1(new_n746), .B2(new_n784), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(G317), .B2(new_n788), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1012), .A2(new_n1015), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1010), .A2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT47), .Z(new_n1021));
  OAI221_X1 g0821(.A(new_n1004), .B1(new_n935), .B2(new_n794), .C1(new_n1021), .C2(new_n814), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1000), .A2(new_n1022), .ZN(G387));
  NOR2_X1   g0823(.A1(new_n989), .A2(new_n675), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n988), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1024), .B1(new_n718), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n943), .A2(new_n655), .A3(new_n738), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n728), .A2(new_n676), .B1(G107), .B2(new_n211), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n238), .A2(new_n296), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n464), .A2(new_n409), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT50), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n676), .B(new_n296), .C1(new_n449), .C2(new_n451), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1033), .A2(new_n732), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1028), .B1(new_n1029), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n727), .B1(new_n1035), .B2(new_n741), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n766), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n371), .A2(new_n756), .B1(new_n1037), .B2(G68), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT113), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n270), .B1(new_n762), .B2(new_n412), .C1(new_n746), .C2(new_n409), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n750), .A2(new_n429), .B1(new_n451), .B2(new_n752), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n781), .A2(new_n466), .B1(new_n744), .B2(new_n352), .ZN(new_n1042));
  OR4_X1    g0842(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n270), .B1(new_n788), .B2(G326), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n781), .A2(new_n780), .B1(new_n752), .B2(new_n782), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G311), .A2(new_n756), .B1(new_n777), .B2(G317), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(KEYINPUT114), .B(G322), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1046), .B1(new_n744), .B2(new_n1047), .C1(new_n769), .C2(new_n784), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT48), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1045), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n1049), .B2(new_n1048), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT49), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1044), .B1(new_n274), .B2(new_n750), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1043), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1036), .B1(new_n1055), .B2(new_n739), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1025), .A2(new_n724), .B1(new_n1027), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1026), .A2(new_n1057), .ZN(G393));
  NAND2_X1  g0858(.A1(new_n982), .A2(new_n990), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(KEYINPUT115), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT115), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n990), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1060), .A2(new_n724), .A3(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n777), .A2(G311), .B1(new_n830), .B2(G317), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT52), .Z(new_n1065));
  OAI221_X1 g0865(.A(new_n359), .B1(new_n1047), .B2(new_n762), .C1(new_n782), .C2(new_n766), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1066), .B(new_n751), .C1(G283), .C2(new_n753), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n756), .A2(G303), .B1(G116), .B2(new_n758), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(KEYINPUT117), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1068), .A2(KEYINPUT117), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1065), .A2(new_n1067), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n752), .A2(new_n449), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n781), .A2(new_n451), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(G50), .C2(new_n756), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n412), .A2(new_n744), .B1(new_n746), .B2(new_n352), .ZN(new_n1075));
  XOR2_X1   g0875(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n1076));
  XNOR2_X1  g0876(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n770), .A2(new_n464), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n270), .B1(new_n816), .B2(new_n762), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n827), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1074), .A2(new_n1077), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n814), .B1(new_n1071), .B2(new_n1081), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n246), .A2(new_n732), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n741), .B1(G97), .B2(new_n673), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n726), .B(new_n1082), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n930), .B2(new_n794), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n989), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n991), .A2(new_n674), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1063), .B(new_n1086), .C1(new_n1087), .C2(new_n1088), .ZN(G390));
  AND3_X1   g0889(.A1(new_n871), .A2(KEYINPUT39), .A3(new_n872), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n880), .A2(new_n884), .ZN(new_n1091));
  AOI21_X1  g0891(.A(KEYINPUT39), .B1(new_n1091), .B2(new_n872), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n1090), .A2(new_n1092), .B1(new_n874), .B2(new_n906), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n704), .A2(new_n668), .A3(new_n810), .A4(new_n917), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n874), .ZN(new_n1095));
  AOI21_X1  g0895(.A(KEYINPUT108), .B1(new_n883), .B2(new_n870), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n876), .B(KEYINPUT38), .C1(new_n881), .C2(new_n882), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n872), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n904), .B1(new_n716), .B2(new_n810), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1095), .B(new_n1098), .C1(new_n1099), .C2(new_n902), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n1093), .A2(new_n1094), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n913), .A2(G330), .A3(new_n810), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1102), .A2(new_n902), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n1093), .B2(new_n1100), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1102), .A2(new_n902), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1094), .A2(new_n1099), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(KEYINPUT118), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT118), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1094), .A2(new_n1099), .A3(new_n1106), .A4(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n704), .A2(new_n668), .A3(new_n810), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n902), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n1104), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n903), .A2(new_n905), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1108), .A2(new_n1110), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n485), .A2(G330), .A3(new_n913), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1116), .A2(new_n910), .A3(new_n638), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n1101), .A2(new_n1105), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1093), .A2(new_n1094), .A3(new_n1100), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT39), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1098), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1114), .A2(new_n917), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1124), .A2(new_n873), .B1(new_n1125), .B2(new_n1095), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n716), .A2(new_n810), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n902), .B1(new_n1127), .B2(new_n905), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1098), .A2(new_n1095), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1103), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1117), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1121), .A2(new_n1122), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1118), .A2(new_n1133), .A3(new_n674), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n836), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n727), .B1(new_n371), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n737), .B1(new_n1124), .B2(new_n873), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n744), .A2(new_n780), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1138), .B(new_n1073), .C1(G107), .C2(new_n756), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n770), .A2(G97), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n359), .B1(new_n746), .B2(new_n274), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G294), .B2(new_n788), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n753), .A2(G87), .B1(new_n749), .B2(G68), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1139), .A2(new_n1140), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(G128), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n781), .A2(new_n352), .B1(new_n744), .B2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT54), .B(G143), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n769), .A2(new_n1147), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n750), .A2(new_n409), .B1(new_n755), .B2(new_n815), .ZN(new_n1149));
  INV_X1    g0949(.A(G125), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n270), .B1(new_n762), .B2(new_n1150), .C1(new_n746), .C2(new_n822), .ZN(new_n1151));
  OR4_X1    g0951(.A1(new_n1146), .A2(new_n1148), .A3(new_n1149), .A4(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n753), .A2(G150), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT53), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1144), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1136), .B(new_n1137), .C1(new_n739), .C2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1156), .B1(new_n1157), .B2(new_n724), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1134), .A2(new_n1158), .ZN(G378));
  AOI21_X1  g0959(.A(new_n726), .B1(new_n409), .B2(new_n836), .ZN(new_n1160));
  OR2_X1    g0960(.A1(new_n270), .A2(G41), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1161), .B(new_n409), .C1(G33), .C2(G41), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n781), .A2(new_n449), .B1(new_n744), .B2(new_n274), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT119), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n746), .A2(new_n259), .B1(new_n780), .B2(new_n762), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n766), .A2(new_n466), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1165), .A2(new_n1166), .A3(new_n1161), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n749), .A2(new_n356), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n753), .A2(G77), .B1(new_n756), .B2(G97), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1164), .A2(new_n1167), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT120), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1162), .B1(new_n1171), .B2(KEYINPUT58), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT121), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1171), .A2(KEYINPUT58), .ZN(new_n1174));
  AOI211_X1 g0974(.A(G33), .B(G41), .C1(new_n788), .C2(G124), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n750), .B2(new_n760), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n1150), .A2(new_n744), .B1(new_n755), .B2(new_n822), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n777), .A2(G128), .B1(new_n1037), .B2(G137), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n752), .B2(new_n1147), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1177), .B(new_n1179), .C1(G150), .C2(new_n758), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1176), .B1(new_n1181), .B2(KEYINPUT59), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(KEYINPUT59), .B2(new_n1181), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1173), .A2(new_n1174), .A3(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n425), .A2(new_n417), .A3(new_n852), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n417), .A2(new_n852), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n420), .A2(new_n424), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1185), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1160), .B1(new_n814), .B2(new_n1184), .C1(new_n1193), .C2(new_n737), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT122), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n888), .A2(new_n915), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT40), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(G330), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n918), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n1200), .B2(new_n1098), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1198), .A2(new_n1201), .A3(new_n1193), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1193), .ZN(new_n1203));
  OAI21_X1  g1003(.A(G330), .B1(new_n885), .B2(new_n918), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1203), .B1(new_n1204), .B2(new_n916), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n908), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n908), .A2(new_n1202), .A3(new_n1205), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1195), .B1(new_n1210), .B2(new_n724), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1117), .B1(new_n1157), .B2(new_n1121), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n908), .A2(new_n1202), .A3(new_n1205), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1202), .A2(new_n1205), .B1(new_n886), .B2(new_n907), .ZN(new_n1214));
  OAI21_X1  g1014(.A(KEYINPUT57), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n674), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1131), .A2(new_n1122), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1132), .B1(new_n1217), .B2(new_n1115), .ZN(new_n1218));
  AOI21_X1  g1018(.A(KEYINPUT57), .B1(new_n1218), .B2(new_n1210), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1211), .B1(new_n1216), .B2(new_n1219), .ZN(G375));
  NOR2_X1   g1020(.A1(new_n917), .A2(new_n737), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n770), .A2(G107), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n359), .B1(new_n762), .B2(new_n784), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G283), .B2(new_n777), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n752), .A2(new_n429), .B1(new_n744), .B2(new_n782), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G116), .B2(new_n756), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n749), .A2(G77), .B1(new_n758), .B2(new_n1002), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1222), .A2(new_n1224), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n270), .B1(new_n762), .B2(new_n1145), .C1(new_n766), .C2(new_n412), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1168), .B1(new_n352), .B2(new_n752), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(G50), .C2(new_n758), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT123), .Z(new_n1232));
  NAND2_X1  g1032(.A1(new_n830), .A2(G132), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n815), .B2(new_n746), .C1(new_n755), .C2(new_n1147), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1228), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n739), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1236), .B(new_n727), .C1(G68), .C2(new_n1135), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n1115), .A2(new_n721), .B1(new_n1221), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1121), .A2(new_n1132), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n993), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1121), .A2(new_n1132), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1239), .B1(new_n1241), .B2(new_n1242), .ZN(G381));
  NAND3_X1  g1043(.A1(new_n1026), .A2(new_n799), .A3(new_n1057), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(G384), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NOR4_X1   g1047(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(G375), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT124), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(G378), .A2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1134), .A2(KEYINPUT124), .A3(new_n1158), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1248), .A2(new_n1249), .A3(new_n1253), .ZN(G407));
  NAND3_X1  g1054(.A1(new_n1249), .A2(new_n1253), .A3(new_n645), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(G407), .A2(G213), .A3(new_n1255), .ZN(G409));
  NAND3_X1  g1056(.A1(new_n1218), .A2(new_n1210), .A3(new_n993), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1211), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1251), .A2(new_n1252), .A3(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(G378), .B(new_n1211), .C1(new_n1216), .C2(new_n1219), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT125), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1115), .A2(KEYINPUT60), .A3(new_n1117), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n674), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1240), .A2(KEYINPUT60), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1242), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1265), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1246), .B1(new_n1268), .B2(new_n1238), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1242), .B1(KEYINPUT60), .B2(new_n1240), .ZN(new_n1270));
  OAI211_X1 g1070(.A(G384), .B(new_n1239), .C1(new_n1270), .C2(new_n1265), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1259), .A2(new_n1260), .A3(KEYINPUT125), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n645), .A2(G213), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1263), .A2(new_n1273), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT63), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT126), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1000), .A2(new_n1022), .A3(G390), .ZN(new_n1281));
  AOI21_X1  g1081(.A(G390), .B1(new_n1000), .B2(new_n1022), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT127), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n799), .B1(new_n1026), .B2(new_n1057), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1283), .B1(new_n1285), .B2(new_n1244), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1245), .A2(new_n1284), .A3(KEYINPUT127), .ZN(new_n1287));
  OAI22_X1  g1087(.A1(new_n1281), .A2(new_n1282), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(G390), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G387), .A2(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1000), .A2(new_n1022), .A3(G390), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1290), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1288), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1261), .A2(new_n1273), .A3(KEYINPUT63), .A4(new_n1275), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1294), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1275), .ZN(new_n1298));
  AND2_X1   g1098(.A1(new_n1298), .A2(G2897), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1269), .A2(new_n1271), .A3(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1299), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1298), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1302), .B1(new_n1303), .B2(new_n1274), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1297), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1276), .A2(KEYINPUT126), .A3(new_n1277), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1280), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1294), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1298), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1273), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(KEYINPUT62), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1311), .B(new_n1295), .C1(new_n1309), .C2(new_n1302), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1276), .A2(KEYINPUT62), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1308), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1307), .A2(new_n1314), .ZN(G405));
  NAND2_X1  g1115(.A1(new_n1253), .A2(G375), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1260), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1317), .B(new_n1272), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(new_n1318), .B(new_n1294), .ZN(G402));
endmodule


