//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n984, new_n985, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1058, new_n1059;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(KEYINPUT1), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G120gat), .ZN(new_n206));
  AND2_X1   g005(.A1(new_n206), .A2(G113gat), .ZN(new_n207));
  XOR2_X1   g006(.A(KEYINPUT68), .B(G113gat), .Z(new_n208));
  AOI21_X1  g007(.A(new_n207), .B1(new_n208), .B2(G120gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n202), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n205), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G169gat), .ZN(new_n214));
  INV_X1    g013(.A(G176gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT23), .ZN(new_n220));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT24), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n225), .B(new_n226), .C1(G183gat), .C2(G190gat), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT25), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n226), .B(new_n230), .ZN(new_n231));
  OR2_X1    g030(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n232));
  INV_X1    g031(.A(G183gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(new_n225), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n237));
  AND4_X1   g036(.A1(KEYINPUT25), .A2(new_n218), .A3(new_n220), .A4(new_n221), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n237), .B1(new_n236), .B2(new_n238), .ZN(new_n240));
  OAI211_X1 g039(.A(KEYINPUT67), .B(new_n229), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(KEYINPUT65), .B(G190gat), .Z(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT27), .B(G183gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT28), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT26), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n219), .B1(new_n247), .B2(new_n221), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n216), .A2(KEYINPUT26), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n250), .B1(G183gat), .B2(G190gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n241), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT66), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n236), .A2(new_n238), .A3(new_n237), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT67), .B1(new_n257), .B2(new_n229), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n213), .B1(new_n253), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G227gat), .ZN(new_n260));
  INV_X1    g059(.A(G233gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n229), .B1(new_n239), .B2(new_n240), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n265), .A2(new_n212), .A3(new_n241), .A4(new_n252), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n259), .A2(new_n262), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT33), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n267), .A2(KEYINPUT69), .A3(new_n268), .ZN(new_n272));
  XNOR2_X1  g071(.A(G15gat), .B(G43gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(G71gat), .B(G99gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n275), .B1(new_n267), .B2(KEYINPUT32), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n271), .A2(new_n272), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n262), .B1(new_n259), .B2(new_n266), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT34), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI211_X1 g079(.A(KEYINPUT34), .B(new_n262), .C1(new_n259), .C2(new_n266), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n267), .B(KEYINPUT32), .C1(new_n268), .C2(new_n275), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n277), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n282), .B1(new_n277), .B2(new_n283), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT36), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n277), .A2(new_n283), .ZN(new_n287));
  INV_X1    g086(.A(new_n282), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT36), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n277), .A2(new_n282), .A3(new_n283), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G78gat), .B(G106gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G155gat), .B(G162gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G155gat), .ZN(new_n298));
  INV_X1    g097(.A(G162gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(KEYINPUT73), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(KEYINPUT2), .ZN(new_n303));
  XOR2_X1   g102(.A(G141gat), .B(G148gat), .Z(new_n304));
  NAND4_X1  g103(.A1(new_n297), .A2(new_n302), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT3), .ZN(new_n306));
  XNOR2_X1  g105(.A(G141gat), .B(G148gat), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n301), .B(new_n300), .C1(new_n307), .C2(KEYINPUT2), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT71), .B(KEYINPUT29), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT80), .ZN(new_n313));
  XNOR2_X1  g112(.A(G197gat), .B(G204gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT22), .ZN(new_n315));
  XNOR2_X1  g114(.A(G211gat), .B(G218gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(KEYINPUT70), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G211gat), .ZN(new_n319));
  INV_X1    g118(.A(G218gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n316), .B(new_n314), .C1(KEYINPUT22), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT70), .B1(new_n315), .B2(new_n317), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n312), .A2(new_n313), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n305), .A2(new_n308), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n315), .A2(new_n317), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n310), .B1(new_n328), .B2(new_n322), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n327), .B1(new_n329), .B2(KEYINPUT3), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n313), .B1(new_n312), .B2(new_n325), .ZN(new_n332));
  INV_X1    g131(.A(G228gat), .ZN(new_n333));
  OAI22_X1  g132(.A1(new_n331), .A2(new_n332), .B1(new_n333), .B2(new_n261), .ZN(new_n334));
  INV_X1    g133(.A(G22gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n333), .A2(new_n261), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n312), .A2(new_n325), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n323), .A2(new_n324), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT29), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT3), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n327), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n305), .A2(KEYINPUT74), .A3(new_n308), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n336), .B(new_n337), .C1(new_n340), .C2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n334), .A2(new_n335), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n335), .B1(new_n334), .B2(new_n345), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n294), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n345), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G22gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(new_n346), .A3(new_n293), .ZN(new_n352));
  XOR2_X1   g151(.A(KEYINPUT31), .B(G50gat), .Z(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n349), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n354), .B1(new_n349), .B2(new_n352), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT81), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n349), .A2(new_n352), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n353), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT81), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n349), .A2(new_n352), .A3(new_n354), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G1gat), .B(G29gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(KEYINPUT0), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(KEYINPUT78), .ZN(new_n366));
  XNOR2_X1  g165(.A(G57gat), .B(G85gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT68), .B(G113gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n370), .A2(new_n206), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n210), .B(new_n202), .C1(new_n371), .C2(new_n207), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n372), .A2(new_n305), .A3(new_n308), .A4(new_n205), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(new_n344), .B2(new_n213), .ZN(new_n374));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT5), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n212), .A2(new_n327), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n373), .A2(KEYINPUT76), .A3(KEYINPUT4), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT76), .B1(new_n373), .B2(KEYINPUT4), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n375), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n342), .A2(KEYINPUT3), .A3(new_n343), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT75), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n342), .A2(KEYINPUT75), .A3(KEYINPUT3), .A4(new_n343), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n309), .A2(new_n212), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT77), .B1(new_n385), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT4), .B1(new_n212), .B2(new_n327), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT76), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n373), .A2(KEYINPUT76), .A3(KEYINPUT4), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n376), .B1(new_n398), .B2(new_n381), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT77), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n390), .B1(new_n386), .B2(new_n387), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n389), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n378), .B1(new_n393), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n379), .A2(KEYINPUT79), .A3(new_n380), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT79), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n406), .B1(new_n373), .B2(KEYINPUT4), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n394), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n402), .A2(new_n409), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n410), .A2(KEYINPUT5), .A3(new_n376), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n369), .B1(new_n404), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n378), .ZN(new_n413));
  AND4_X1   g212(.A1(new_n400), .A2(new_n402), .A3(new_n375), .A4(new_n384), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n400), .B1(new_n399), .B2(new_n402), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n411), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(new_n368), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT6), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n412), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(KEYINPUT6), .B(new_n369), .C1(new_n404), .C2(new_n411), .ZN(new_n421));
  XNOR2_X1  g220(.A(G8gat), .B(G36gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(G64gat), .B(G92gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n263), .A2(new_n252), .ZN(new_n425));
  NAND2_X1  g224(.A1(G226gat), .A2(G233gat), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT72), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n425), .A2(KEYINPUT72), .A3(new_n427), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n311), .B1(new_n253), .B2(new_n258), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n426), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n338), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n265), .A2(new_n427), .A3(new_n241), .A4(new_n252), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n425), .A2(new_n339), .A3(new_n426), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n325), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n424), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n438), .ZN(new_n440));
  INV_X1    g239(.A(new_n424), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n430), .A2(new_n431), .B1(new_n433), .B2(new_n426), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n440), .B(new_n441), .C1(new_n442), .C2(new_n338), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n439), .A2(KEYINPUT30), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n432), .A2(new_n434), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n438), .B1(new_n445), .B2(new_n325), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT30), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(new_n447), .A3(new_n441), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n420), .A2(new_n421), .B1(new_n444), .B2(new_n448), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n286), .B(new_n292), .C1(new_n363), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n420), .A2(new_n421), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n440), .B1(new_n442), .B2(new_n338), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n441), .B1(new_n453), .B2(KEYINPUT37), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT37), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT84), .B1(new_n446), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT84), .ZN(new_n457));
  NOR4_X1   g256(.A1(new_n435), .A2(new_n457), .A3(KEYINPUT37), .A4(new_n438), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n454), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT38), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n436), .A2(new_n437), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n455), .B1(new_n461), .B2(new_n325), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n462), .B1(new_n325), .B2(new_n442), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n441), .A2(KEYINPUT38), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n463), .B(new_n464), .C1(new_n456), .C2(new_n458), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n452), .A2(new_n460), .A3(new_n443), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n359), .A2(new_n361), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT40), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n375), .B(new_n373), .C1(new_n344), .C2(new_n213), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT39), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT83), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n389), .A2(new_n401), .B1(new_n408), .B2(new_n394), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT82), .B1(new_n474), .B2(new_n375), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT82), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n410), .A2(new_n476), .A3(new_n376), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n368), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT39), .B1(new_n475), .B2(new_n477), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n469), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n475), .A2(new_n477), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT39), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n484), .A2(KEYINPUT40), .A3(new_n368), .A4(new_n478), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n481), .A2(new_n412), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n444), .A2(new_n448), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n468), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n450), .B1(new_n466), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT85), .B1(new_n284), .B2(new_n285), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT85), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n289), .A2(new_n492), .A3(new_n291), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NOR3_X1   g293(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT35), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(new_n451), .A3(new_n487), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n284), .A2(new_n285), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n498), .A2(new_n449), .A3(new_n468), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n494), .A2(new_n497), .B1(new_n499), .B2(KEYINPUT35), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n490), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G190gat), .B(G218gat), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G99gat), .B(G106gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507));
  INV_X1    g306(.A(G85gat), .ZN(new_n508));
  INV_X1    g307(.A(G92gat), .ZN(new_n509));
  AOI22_X1  g308(.A1(KEYINPUT8), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT93), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT7), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n512), .B1(new_n513), .B2(KEYINPUT92), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT94), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT92), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT7), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT94), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(new_n512), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g319(.A(G85gat), .B(G92gat), .C1(new_n512), .C2(new_n513), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n511), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G85gat), .A2(G92gat), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n523), .B1(KEYINPUT93), .B2(KEYINPUT7), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n515), .A2(new_n519), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n506), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n518), .B1(new_n517), .B2(new_n512), .ZN(new_n527));
  AOI211_X1 g326(.A(KEYINPUT93), .B(KEYINPUT94), .C1(new_n516), .C2(KEYINPUT7), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n521), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AND4_X1   g328(.A1(new_n506), .A2(new_n529), .A3(new_n525), .A4(new_n510), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G29gat), .A2(G36gat), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NOR3_X1   g333(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT15), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G43gat), .B(G50gat), .ZN(new_n539));
  INV_X1    g338(.A(new_n532), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT14), .ZN(new_n541));
  INV_X1    g340(.A(G29gat), .ZN(new_n542));
  INV_X1    g341(.A(G36gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n540), .B1(new_n544), .B2(new_n533), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT15), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n538), .A2(new_n539), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n539), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n545), .A2(new_n548), .A3(KEYINPUT15), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n505), .B1(new_n531), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n529), .A2(new_n525), .A3(new_n510), .ZN(new_n552));
  INV_X1    g351(.A(new_n506), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n529), .A2(new_n506), .A3(new_n525), .A4(new_n510), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT17), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n547), .A2(new_n557), .A3(new_n549), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n547), .B2(new_n549), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n556), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n503), .B1(new_n551), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT95), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n539), .B1(new_n545), .B2(KEYINPUT15), .ZN(new_n564));
  AOI211_X1 g363(.A(new_n537), .B(new_n540), .C1(new_n544), .C2(new_n533), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n549), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT17), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n547), .A2(new_n557), .A3(new_n549), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n568), .A2(new_n569), .B1(new_n555), .B2(new_n554), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n550), .A2(new_n554), .A3(new_n555), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n504), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n563), .B1(new_n573), .B2(new_n503), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n551), .A2(new_n563), .A3(new_n560), .A4(new_n503), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n562), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n560), .A2(new_n504), .A3(new_n571), .A4(new_n503), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT95), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n575), .ZN(new_n582));
  INV_X1    g381(.A(new_n578), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n582), .A2(new_n583), .A3(new_n562), .ZN(new_n584));
  XOR2_X1   g383(.A(G134gat), .B(G162gat), .Z(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n579), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n583), .B1(new_n582), .B2(new_n562), .ZN(new_n588));
  AOI211_X1 g387(.A(new_n578), .B(new_n561), .C1(new_n581), .C2(new_n575), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n585), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT87), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n335), .A2(G15gat), .ZN(new_n594));
  INV_X1    g393(.A(G15gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(G22gat), .ZN(new_n596));
  INV_X1    g395(.A(G1gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT16), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n594), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT86), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(G1gat), .B1(new_n594), .B2(new_n596), .ZN(new_n602));
  OAI21_X1  g401(.A(G8gat), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G15gat), .B(G22gat), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT86), .B1(new_n604), .B2(new_n598), .ZN(new_n605));
  INV_X1    g404(.A(new_n602), .ZN(new_n606));
  INV_X1    g405(.A(G8gat), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n550), .A2(new_n593), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n593), .B1(new_n550), .B2(new_n609), .ZN(new_n611));
  OAI22_X1  g410(.A1(new_n610), .A2(new_n611), .B1(new_n609), .B2(new_n550), .ZN(new_n612));
  NAND2_X1  g411(.A1(G229gat), .A2(G233gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(KEYINPUT13), .Z(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n609), .B1(new_n566), .B2(new_n567), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT87), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n550), .A2(new_n593), .A3(new_n609), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n609), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n620), .B1(new_n558), .B2(new_n559), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n619), .A2(KEYINPUT18), .A3(new_n613), .A4(new_n621), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n619), .A2(new_n613), .A3(new_n621), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT18), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G113gat), .B(G141gat), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT11), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n214), .ZN(new_n630));
  INV_X1    g429(.A(G197gat), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n629), .B(G169gat), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n633), .A2(G197gat), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT12), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(G197gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n630), .A2(new_n631), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT12), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n623), .B(new_n626), .C1(KEYINPUT88), .C2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n615), .A2(new_n622), .A3(KEYINPUT88), .ZN(new_n642));
  INV_X1    g441(.A(new_n640), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n615), .A2(new_n622), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n568), .A2(new_n569), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n617), .A2(new_n618), .B1(new_n645), .B2(new_n620), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT18), .B1(new_n646), .B2(new_n613), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n642), .B(new_n643), .C1(new_n644), .C2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n641), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(G230gat), .A2(G233gat), .ZN(new_n651));
  NAND2_X1  g450(.A1(G71gat), .A2(G78gat), .ZN(new_n652));
  OR2_X1    g451(.A1(G71gat), .A2(G78gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(G57gat), .B(G64gat), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT9), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n652), .B(new_n653), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(KEYINPUT89), .A2(G57gat), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT90), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT90), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n659), .A2(KEYINPUT89), .A3(G57gat), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n658), .A2(new_n660), .A3(G64gat), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n652), .B1(new_n653), .B2(new_n655), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(G64gat), .B1(new_n658), .B2(new_n660), .ZN(new_n664));
  OAI211_X1 g463(.A(KEYINPUT96), .B(new_n656), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n656), .B1(new_n663), .B2(new_n664), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT96), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n665), .B(new_n668), .C1(new_n526), .C2(new_n530), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n554), .A2(new_n667), .A3(new_n666), .A4(new_n555), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT10), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT10), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n556), .A2(new_n672), .A3(new_n666), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n651), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n651), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n669), .A2(new_n670), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(G120gat), .B(G148gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(G176gat), .B(G204gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n674), .A2(new_n676), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n680), .B1(new_n674), .B2(new_n676), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n650), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g485(.A(G183gat), .B(G211gat), .Z(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT21), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n666), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(G231gat), .A2(G233gat), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n690), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(G127gat), .B(G155gat), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n693), .A2(new_n695), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n699));
  NOR3_X1   g498(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n699), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n693), .A2(new_n695), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(new_n696), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n688), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n620), .B1(new_n689), .B2(new_n666), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT91), .Z(new_n706));
  OAI21_X1  g505(.A(new_n699), .B1(new_n697), .B2(new_n698), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n696), .A2(new_n702), .A3(new_n701), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(new_n708), .A3(new_n687), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n704), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n706), .B1(new_n704), .B2(new_n709), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n592), .A2(new_n686), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n501), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n452), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(G1gat), .ZN(G1324gat));
  INV_X1    g515(.A(new_n487), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT16), .B(G8gat), .Z(new_n718));
  NAND3_X1  g517(.A1(new_n714), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(KEYINPUT42), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT42), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n714), .A2(new_n717), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n721), .B1(new_n722), .B2(G8gat), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n720), .B1(new_n719), .B2(new_n723), .ZN(G1325gat));
  NAND3_X1  g523(.A1(new_n714), .A2(new_n595), .A3(new_n494), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n286), .A2(new_n292), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n501), .A2(new_n727), .A3(new_n713), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n725), .B1(new_n728), .B2(new_n595), .ZN(G1326gat));
  INV_X1    g528(.A(new_n363), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(KEYINPUT43), .B(G22gat), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1327gat));
  NAND2_X1  g532(.A1(new_n489), .A2(new_n466), .ZN(new_n734));
  INV_X1    g533(.A(new_n450), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n737));
  INV_X1    g536(.A(new_n494), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n738), .B2(new_n496), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n592), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n712), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n686), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n744), .A2(G29gat), .A3(new_n451), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT97), .B(KEYINPUT45), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(new_n747));
  OAI211_X1 g546(.A(KEYINPUT98), .B(new_n591), .C1(new_n490), .C2(new_n500), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n463), .A2(new_n464), .ZN(new_n751));
  INV_X1    g550(.A(new_n458), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n457), .B1(new_n453), .B2(KEYINPUT37), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n443), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n754), .A2(new_n451), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n488), .B1(new_n756), .B2(new_n460), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n496), .B1(new_n491), .B2(new_n493), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT35), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n467), .A2(new_n284), .A3(new_n285), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n759), .B1(new_n760), .B2(new_n449), .ZN(new_n761));
  OAI22_X1  g560(.A1(new_n757), .A2(new_n450), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n762), .A2(KEYINPUT98), .A3(KEYINPUT44), .A4(new_n591), .ZN(new_n763));
  AND4_X1   g562(.A1(new_n452), .A2(new_n750), .A3(new_n763), .A4(new_n743), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n747), .B1(new_n542), .B2(new_n764), .ZN(G1328gat));
  NOR3_X1   g564(.A1(new_n744), .A2(G36gat), .A3(new_n487), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT46), .ZN(new_n767));
  AND4_X1   g566(.A1(new_n717), .A2(new_n750), .A3(new_n763), .A4(new_n743), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n543), .B2(new_n768), .ZN(G1329gat));
  NAND4_X1  g568(.A1(new_n750), .A2(new_n726), .A3(new_n763), .A4(new_n743), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G43gat), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n738), .A2(G43gat), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n762), .A2(new_n772), .A3(new_n591), .A4(new_n743), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT99), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(KEYINPUT47), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n771), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT100), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(KEYINPUT99), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT100), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n771), .A2(new_n781), .A3(new_n776), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n778), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n780), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n781), .B1(new_n771), .B2(new_n776), .ZN(new_n785));
  AOI211_X1 g584(.A(KEYINPUT100), .B(new_n775), .C1(new_n770), .C2(G43gat), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n783), .A2(new_n787), .ZN(G1330gat));
  NAND3_X1  g587(.A1(new_n750), .A2(new_n763), .A3(new_n743), .ZN(new_n789));
  OAI21_X1  g588(.A(G50gat), .B1(new_n789), .B2(new_n468), .ZN(new_n790));
  INV_X1    g589(.A(G50gat), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n740), .A2(new_n791), .A3(new_n730), .A4(new_n743), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(KEYINPUT48), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(G50gat), .B1(new_n789), .B2(new_n363), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n794), .A2(new_n792), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n795), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g595(.A1(new_n592), .A2(new_n712), .A3(new_n650), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n501), .A2(new_n684), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT101), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n451), .B(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g601(.A(KEYINPUT102), .B(G57gat), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n802), .B(new_n803), .ZN(G1332gat));
  INV_X1    g603(.A(KEYINPUT49), .ZN(new_n805));
  INV_X1    g604(.A(G64gat), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n717), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n798), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT103), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n798), .A2(KEYINPUT103), .A3(new_n808), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT104), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT104), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n811), .A2(new_n815), .A3(new_n812), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n814), .A2(new_n805), .A3(new_n806), .A4(new_n816), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n811), .A2(new_n815), .A3(new_n812), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n815), .B1(new_n811), .B2(new_n812), .ZN(new_n819));
  OAI22_X1  g618(.A1(new_n818), .A2(new_n819), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n817), .A2(new_n820), .ZN(G1333gat));
  NAND2_X1  g620(.A1(new_n798), .A2(new_n726), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n738), .A2(G71gat), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n822), .A2(G71gat), .B1(new_n798), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g624(.A1(new_n798), .A2(new_n730), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g626(.A1(new_n712), .A2(new_n649), .A3(new_n684), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n750), .A2(new_n763), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(G85gat), .B1(new_n829), .B2(new_n451), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n712), .A2(new_n649), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n762), .A2(new_n591), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n834), .A2(KEYINPUT105), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n740), .A2(KEYINPUT51), .A3(new_n831), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n836), .B1(new_n834), .B2(KEYINPUT105), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n452), .A2(new_n508), .A3(new_n685), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n830), .B1(new_n838), .B2(new_n839), .ZN(G1336gat));
  INV_X1    g639(.A(KEYINPUT52), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n750), .A2(new_n717), .A3(new_n763), .A4(new_n828), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(G92gat), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n717), .A2(new_n509), .A3(new_n685), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n841), .B(new_n843), .C1(new_n838), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n834), .A2(new_n836), .ZN(new_n846));
  INV_X1    g645(.A(new_n844), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT106), .B1(new_n849), .B2(KEYINPUT52), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT106), .ZN(new_n851));
  AOI211_X1 g650(.A(new_n851), .B(new_n841), .C1(new_n843), .C2(new_n848), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n845), .B1(new_n850), .B2(new_n852), .ZN(G1337gat));
  OR2_X1    g652(.A1(new_n829), .A2(new_n727), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT107), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(G99gat), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n854), .A2(KEYINPUT107), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n684), .A2(G99gat), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n494), .A2(new_n858), .ZN(new_n859));
  OAI22_X1  g658(.A1(new_n856), .A2(new_n857), .B1(new_n838), .B2(new_n859), .ZN(G1338gat));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n861));
  OAI21_X1  g660(.A(G106gat), .B1(new_n829), .B2(new_n468), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n468), .A2(G106gat), .A3(new_n684), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n861), .B(new_n862), .C1(new_n838), .C2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT109), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n750), .A2(new_n730), .A3(new_n763), .A4(new_n828), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n867), .A2(G106gat), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n863), .B(KEYINPUT108), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n846), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n866), .B(KEYINPUT53), .C1(new_n868), .C2(new_n870), .ZN(new_n871));
  AOI22_X1  g670(.A1(G106gat), .A2(new_n867), .B1(new_n846), .B2(new_n869), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT109), .B1(new_n872), .B2(new_n861), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n865), .A2(new_n871), .A3(new_n873), .ZN(G1339gat));
  NOR2_X1   g673(.A1(new_n797), .A2(new_n685), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n668), .A2(new_n665), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n670), .B1(new_n531), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n672), .ZN(new_n878));
  INV_X1    g677(.A(new_n673), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n879), .A3(new_n675), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n674), .A3(KEYINPUT54), .ZN(new_n881));
  XOR2_X1   g680(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n882));
  OAI211_X1 g681(.A(new_n651), .B(new_n882), .C1(new_n671), .C2(new_n673), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n881), .A2(KEYINPUT55), .A3(new_n679), .A4(new_n883), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n884), .A2(new_n681), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n626), .A2(new_n615), .A3(new_n622), .A4(new_n640), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n636), .A2(new_n637), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n646), .A2(new_n613), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n612), .A2(new_n614), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT55), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n881), .A2(new_n679), .A3(new_n883), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n588), .A2(new_n589), .A3(new_n585), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n586), .B1(new_n579), .B2(new_n584), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n885), .B(new_n894), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT111), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n880), .A2(KEYINPUT54), .A3(new_n674), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n679), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n892), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n649), .A2(new_n681), .A3(new_n901), .A4(new_n884), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n684), .A2(new_n891), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n592), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT111), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n591), .A2(new_n907), .A3(new_n885), .A4(new_n894), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n898), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n875), .B1(new_n909), .B2(new_n741), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n730), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n717), .A2(new_n451), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n494), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(G113gat), .B1(new_n913), .B2(new_n650), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n909), .A2(new_n741), .ZN(new_n915));
  INV_X1    g714(.A(new_n875), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(new_n487), .A3(new_n801), .ZN(new_n918));
  INV_X1    g717(.A(new_n760), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT112), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n649), .A2(new_n208), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n914), .B1(new_n921), .B2(new_n922), .ZN(G1340gat));
  OAI21_X1  g722(.A(G120gat), .B1(new_n913), .B2(new_n684), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n684), .A2(G120gat), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT113), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n924), .B1(new_n921), .B2(new_n926), .ZN(G1341gat));
  INV_X1    g726(.A(G127gat), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n913), .A2(new_n928), .A3(new_n741), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n920), .A2(new_n712), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n930), .A2(KEYINPUT114), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n931), .A2(G127gat), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(KEYINPUT114), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(G1342gat));
  NOR4_X1   g733(.A1(new_n918), .A2(G134gat), .A3(new_n919), .A4(new_n592), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT56), .ZN(new_n936));
  OAI21_X1  g735(.A(G134gat), .B1(new_n913), .B2(new_n592), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1343gat));
  INV_X1    g737(.A(G141gat), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n727), .A2(new_n912), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n917), .A2(KEYINPUT57), .A3(new_n730), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT57), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n942), .B1(new_n910), .B2(new_n468), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n940), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n939), .B1(new_n944), .B2(new_n649), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n727), .A2(new_n467), .ZN(new_n946));
  NOR4_X1   g745(.A1(new_n918), .A2(G141gat), .A3(new_n650), .A4(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(KEYINPUT58), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  OR2_X1    g747(.A1(new_n948), .A2(KEYINPUT115), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(KEYINPUT115), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n947), .A2(KEYINPUT116), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n947), .A2(KEYINPUT116), .ZN(new_n952));
  OR3_X1    g751(.A1(new_n951), .A2(new_n952), .A3(KEYINPUT58), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT117), .ZN(new_n954));
  INV_X1    g753(.A(new_n944), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(new_n650), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n944), .A2(KEYINPUT117), .A3(new_n649), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n939), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI211_X1 g757(.A(new_n949), .B(new_n950), .C1(new_n953), .C2(new_n958), .ZN(G1344gat));
  NOR2_X1   g758(.A1(new_n918), .A2(new_n946), .ZN(new_n960));
  INV_X1    g759(.A(G148gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n960), .A2(new_n961), .A3(new_n685), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n962), .A2(KEYINPUT118), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(KEYINPUT118), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT59), .ZN(new_n965));
  AOI22_X1  g764(.A1(new_n641), .A2(new_n648), .B1(new_n893), .B2(new_n892), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n903), .B1(new_n966), .B2(new_n885), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n897), .B1(new_n967), .B2(new_n591), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n712), .B1(new_n968), .B2(KEYINPUT119), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT119), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n897), .B(new_n970), .C1(new_n967), .C2(new_n591), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n875), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n942), .B1(new_n972), .B2(new_n363), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n917), .A2(KEYINPUT57), .A3(new_n467), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n975), .A2(new_n727), .A3(new_n685), .A4(new_n912), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n965), .B1(new_n976), .B2(G148gat), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n965), .A2(G148gat), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n978), .B1(new_n944), .B2(new_n685), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n963), .B(new_n964), .C1(new_n977), .C2(new_n979), .ZN(G1345gat));
  OAI21_X1  g779(.A(G155gat), .B1(new_n955), .B2(new_n741), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n960), .A2(new_n298), .A3(new_n712), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1346gat));
  OAI21_X1  g782(.A(G162gat), .B1(new_n955), .B2(new_n592), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n960), .A2(new_n299), .A3(new_n591), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(G1347gat));
  NAND4_X1  g785(.A1(new_n911), .A2(new_n717), .A3(new_n494), .A4(new_n800), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n987), .A2(new_n214), .A3(new_n650), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n917), .A2(KEYINPUT120), .A3(new_n451), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT120), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n990), .B1(new_n910), .B2(new_n452), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n487), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n992), .A2(new_n760), .A3(new_n649), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n988), .B1(new_n993), .B2(new_n214), .ZN(G1348gat));
  NAND3_X1  g793(.A1(new_n992), .A2(new_n760), .A3(new_n685), .ZN(new_n995));
  AND3_X1   g794(.A1(new_n995), .A2(KEYINPUT121), .A3(new_n215), .ZN(new_n996));
  AOI21_X1  g795(.A(KEYINPUT121), .B1(new_n995), .B2(new_n215), .ZN(new_n997));
  NOR3_X1   g796(.A1(new_n987), .A2(new_n215), .A3(new_n684), .ZN(new_n998));
  NOR3_X1   g797(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(G1349gat));
  NAND4_X1  g798(.A1(new_n992), .A2(new_n243), .A3(new_n760), .A4(new_n712), .ZN(new_n1000));
  OAI21_X1  g799(.A(G183gat), .B1(new_n987), .B2(new_n741), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g801(.A(KEYINPUT122), .B(KEYINPUT60), .Z(new_n1003));
  OR3_X1    g802(.A1(new_n1002), .A2(KEYINPUT123), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g803(.A(KEYINPUT123), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1002), .A2(KEYINPUT60), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(G1350gat));
  OAI21_X1  g806(.A(G190gat), .B1(new_n987), .B2(new_n592), .ZN(new_n1008));
  XNOR2_X1  g807(.A(new_n1008), .B(KEYINPUT61), .ZN(new_n1009));
  NAND4_X1  g808(.A1(new_n992), .A2(new_n242), .A3(new_n760), .A4(new_n591), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1009), .A2(new_n1010), .ZN(G1351gat));
  NAND3_X1  g810(.A1(new_n727), .A2(new_n800), .A3(new_n717), .ZN(new_n1012));
  AOI21_X1  g811(.A(new_n1012), .B1(new_n973), .B2(new_n974), .ZN(new_n1013));
  INV_X1    g812(.A(new_n1013), .ZN(new_n1014));
  OAI21_X1  g813(.A(G197gat), .B1(new_n1014), .B2(new_n650), .ZN(new_n1015));
  AOI211_X1 g814(.A(new_n487), .B(new_n946), .C1(new_n989), .C2(new_n991), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n1016), .A2(new_n631), .A3(new_n649), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1015), .A2(new_n1017), .ZN(G1352gat));
  NOR2_X1   g817(.A1(new_n684), .A2(G204gat), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g819(.A(new_n1012), .ZN(new_n1021));
  NAND3_X1  g820(.A1(new_n975), .A2(new_n685), .A3(new_n1021), .ZN(new_n1022));
  AOI22_X1  g821(.A1(new_n1020), .A2(KEYINPUT62), .B1(G204gat), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g822(.A(KEYINPUT62), .ZN(new_n1024));
  INV_X1    g823(.A(new_n946), .ZN(new_n1025));
  NAND4_X1  g824(.A1(new_n992), .A2(new_n1024), .A3(new_n1025), .A4(new_n1019), .ZN(new_n1026));
  INV_X1    g825(.A(KEYINPUT124), .ZN(new_n1027));
  NAND2_X1  g826(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g827(.A1(new_n1016), .A2(KEYINPUT124), .A3(new_n1024), .A4(new_n1019), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g829(.A1(new_n1023), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g830(.A(KEYINPUT125), .ZN(new_n1032));
  NAND2_X1  g831(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g832(.A1(new_n1023), .A2(new_n1030), .A3(KEYINPUT125), .ZN(new_n1034));
  NAND2_X1  g833(.A1(new_n1033), .A2(new_n1034), .ZN(G1353gat));
  INV_X1    g834(.A(KEYINPUT63), .ZN(new_n1036));
  AOI21_X1  g835(.A(new_n591), .B1(new_n904), .B2(new_n902), .ZN(new_n1037));
  AND2_X1   g836(.A1(new_n886), .A2(new_n890), .ZN(new_n1038));
  NAND4_X1  g837(.A1(new_n901), .A2(new_n1038), .A3(new_n681), .A4(new_n884), .ZN(new_n1039));
  AOI21_X1  g838(.A(new_n1039), .B1(new_n587), .B2(new_n590), .ZN(new_n1040));
  OAI21_X1  g839(.A(KEYINPUT119), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g840(.A1(new_n1041), .A2(new_n741), .A3(new_n971), .ZN(new_n1042));
  NAND2_X1  g841(.A1(new_n1042), .A2(new_n916), .ZN(new_n1043));
  AOI21_X1  g842(.A(KEYINPUT57), .B1(new_n1043), .B2(new_n730), .ZN(new_n1044));
  NOR3_X1   g843(.A1(new_n910), .A2(new_n942), .A3(new_n468), .ZN(new_n1045));
  OAI211_X1 g844(.A(new_n712), .B(new_n1021), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g845(.A(KEYINPUT126), .ZN(new_n1047));
  OAI21_X1  g846(.A(G211gat), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g847(.A(KEYINPUT126), .B1(new_n1013), .B2(new_n712), .ZN(new_n1049));
  OAI21_X1  g848(.A(new_n1036), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g849(.A1(new_n1050), .A2(KEYINPUT127), .ZN(new_n1051));
  INV_X1    g850(.A(KEYINPUT127), .ZN(new_n1052));
  OAI211_X1 g851(.A(new_n1052), .B(new_n1036), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1053));
  OR3_X1    g852(.A1(new_n1048), .A2(new_n1049), .A3(new_n1036), .ZN(new_n1054));
  NAND3_X1  g853(.A1(new_n1051), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g854(.A1(new_n1016), .A2(new_n319), .A3(new_n712), .ZN(new_n1056));
  NAND2_X1  g855(.A1(new_n1055), .A2(new_n1056), .ZN(G1354gat));
  OAI21_X1  g856(.A(G218gat), .B1(new_n1014), .B2(new_n592), .ZN(new_n1058));
  NAND3_X1  g857(.A1(new_n1016), .A2(new_n320), .A3(new_n591), .ZN(new_n1059));
  NAND2_X1  g858(.A1(new_n1058), .A2(new_n1059), .ZN(G1355gat));
endmodule


