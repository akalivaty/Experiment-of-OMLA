//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 0 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n609, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  OR2_X1    g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(new_n461), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n467), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT64), .B1(new_n471), .B2(new_n461), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AND2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT64), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n478), .A2(new_n479), .A3(G2105), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n470), .B1(new_n472), .B2(new_n480), .ZN(G160));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n468), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT65), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G112), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n476), .A2(new_n461), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G124), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n484), .A2(new_n495), .A3(G138), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n461), .C1(new_n474), .C2(new_n475), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n500), .B1(new_n461), .B2(G114), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(KEYINPUT66), .A3(G2105), .ZN(new_n503));
  OR2_X1    g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n501), .A2(new_n503), .A3(new_n504), .A4(G2104), .ZN(new_n505));
  OAI211_X1 g080(.A(G126), .B(G2105), .C1(new_n474), .C2(new_n475), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n499), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  XOR2_X1   g085(.A(KEYINPUT5), .B(G543), .Z(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G651), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n517), .B(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(G543), .A3(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G50), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n519), .A2(new_n520), .A3(new_n512), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G88), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n515), .A2(new_n523), .A3(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND3_X1  g103(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n524), .B2(new_n533), .ZN(new_n534));
  OAI221_X1 g109(.A(new_n529), .B1(new_n530), .B2(new_n521), .C1(new_n534), .C2(KEYINPUT68), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(KEYINPUT68), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n537), .ZN(G168));
  AOI22_X1  g113(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n514), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n525), .A2(G90), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n522), .A2(G52), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  AOI22_X1  g119(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n514), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n525), .A2(G81), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n522), .A2(G43), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND4_X1  g130(.A1(new_n519), .A2(G53), .A3(G543), .A4(new_n520), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  XNOR2_X1  g133(.A(KEYINPUT69), .B(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n511), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n525), .A2(G91), .B1(G651), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(G299));
  INV_X1    g137(.A(KEYINPUT70), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n563), .B1(new_n535), .B2(new_n537), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n534), .A2(KEYINPUT68), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n529), .B1(new_n521), .B2(new_n530), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n567), .A2(KEYINPUT70), .A3(new_n536), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G286));
  NAND4_X1  g145(.A1(new_n519), .A2(G49), .A3(G543), .A4(new_n520), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n519), .A2(new_n512), .A3(G87), .A4(new_n520), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  NAND4_X1  g149(.A1(new_n519), .A2(G48), .A3(G543), .A4(new_n520), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n519), .A2(new_n512), .A3(G86), .A4(new_n520), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n575), .B(new_n576), .C1(new_n577), .C2(new_n514), .ZN(G305));
  AOI22_X1  g153(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n514), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT71), .ZN(new_n581));
  XOR2_X1   g156(.A(KEYINPUT72), .B(G47), .Z(new_n582));
  AOI22_X1  g157(.A1(G85), .A2(new_n525), .B1(new_n522), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(G290));
  INV_X1    g159(.A(G868), .ZN(new_n585));
  NOR2_X1   g160(.A1(G301), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n525), .A2(KEYINPUT10), .A3(G92), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n588));
  INV_X1    g163(.A(G92), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n524), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g166(.A(KEYINPUT74), .B(G66), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n512), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT73), .Z(new_n595));
  AOI21_X1  g170(.A(new_n514), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(new_n522), .B2(G54), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT75), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n591), .A2(KEYINPUT75), .A3(new_n597), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n586), .B1(new_n603), .B2(new_n585), .ZN(G284));
  XNOR2_X1  g179(.A(G284), .B(KEYINPUT76), .ZN(G321));
  NOR2_X1   g180(.A1(G299), .A2(G868), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(new_n569), .B2(G868), .ZN(G297));
  AOI21_X1  g182(.A(new_n606), .B1(new_n569), .B2(G868), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n603), .B1(new_n609), .B2(G860), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT77), .ZN(G148));
  NAND3_X1  g186(.A1(new_n600), .A2(new_n609), .A3(new_n601), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n467), .A2(new_n463), .ZN(new_n616));
  XOR2_X1   g191(.A(KEYINPUT78), .B(KEYINPUT12), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n491), .A2(G123), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n461), .A2(G111), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n483), .A2(new_n485), .ZN(new_n624));
  INV_X1    g199(.A(G135), .ZN(new_n625));
  OAI221_X1 g200(.A(new_n621), .B1(new_n622), .B2(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n620), .A2(G2100), .B1(G2096), .B2(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(G2096), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n627), .B(new_n628), .C1(G2100), .C2(new_n620), .ZN(G156));
  XOR2_X1   g204(.A(KEYINPUT15), .B(G2435), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2427), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT80), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT79), .B(KEYINPUT14), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n631), .A2(new_n633), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT81), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n638), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2443), .B(G2446), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT82), .Z(new_n646));
  INV_X1    g221(.A(G14), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n647), .B1(new_n643), .B2(new_n644), .ZN(new_n648));
  AND2_X1   g223(.A1(new_n646), .A2(new_n648), .ZN(G401));
  XOR2_X1   g224(.A(KEYINPUT83), .B(KEYINPUT18), .Z(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT17), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  INV_X1    g232(.A(new_n650), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n657), .B1(new_n653), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2096), .B(G2100), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(G1971), .B(G1976), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1956), .B(G2474), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1961), .B(G1966), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  NOR3_X1   g243(.A1(new_n664), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n664), .A2(new_n667), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT20), .Z(new_n671));
  AOI211_X1 g246(.A(new_n669), .B(new_n671), .C1(new_n664), .C2(new_n668), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G1981), .ZN(new_n673));
  XOR2_X1   g248(.A(G1991), .B(G1996), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT86), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n673), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n673), .A2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT87), .B(G1986), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  OR3_X1    g258(.A1(new_n680), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n680), .B2(new_n681), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(G229));
  NAND2_X1  g261(.A1(new_n486), .A2(G139), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT94), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT25), .ZN(new_n690));
  NAND2_X1  g265(.A1(G115), .A2(G2104), .ZN(new_n691));
  INV_X1    g266(.A(G127), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n476), .B2(new_n692), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n693), .A2(KEYINPUT95), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n461), .B1(new_n693), .B2(KEYINPUT95), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n690), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n688), .A2(new_n696), .ZN(new_n697));
  MUX2_X1   g272(.A(G33), .B(new_n697), .S(G29), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT96), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G2072), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G4), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(new_n603), .B2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(G1348), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G26), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n491), .A2(G128), .ZN(new_n710));
  NOR2_X1   g285(.A1(G104), .A2(G2105), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT92), .Z(new_n712));
  OAI21_X1  g287(.A(G2104), .B1(new_n461), .B2(G116), .ZN(new_n713));
  INV_X1    g288(.A(G140), .ZN(new_n714));
  OAI221_X1 g289(.A(new_n710), .B1(new_n712), .B2(new_n713), .C1(new_n624), .C2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT93), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n709), .B1(new_n717), .B2(new_n707), .ZN(new_n718));
  INV_X1    g293(.A(G2067), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT98), .B(KEYINPUT23), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n701), .A2(G20), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G299), .B2(G16), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1956), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n701), .A2(G21), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G168), .B2(new_n701), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G1966), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(G1966), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n720), .A2(new_n725), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n550), .A2(G16), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G16), .B2(G19), .ZN(new_n732));
  INV_X1    g307(.A(G1341), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n701), .A2(G5), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G171), .B2(new_n701), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1961), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT24), .ZN(new_n738));
  INV_X1    g313(.A(G34), .ZN(new_n739));
  AOI21_X1  g314(.A(G29), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n738), .B2(new_n739), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G160), .B2(new_n707), .ZN(new_n742));
  AOI211_X1 g317(.A(new_n734), .B(new_n737), .C1(G2084), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(G162), .A2(G29), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G29), .B2(G35), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT29), .B(G2090), .Z(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n707), .A2(G27), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G164), .B2(new_n707), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(G2078), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT31), .B(G11), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n752), .A2(G28), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n707), .B1(new_n752), .B2(G28), .ZN(new_n754));
  OAI221_X1 g329(.A(new_n751), .B1(new_n753), .B2(new_n754), .C1(new_n626), .C2(new_n707), .ZN(new_n755));
  AOI211_X1 g330(.A(new_n750), .B(new_n755), .C1(new_n732), .C2(new_n733), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n749), .A2(G2078), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n745), .A2(new_n746), .ZN(new_n758));
  AND4_X1   g333(.A1(new_n747), .A2(new_n756), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n742), .A2(G2084), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT97), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n486), .A2(G141), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT26), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n463), .A2(G105), .ZN(new_n765));
  AOI211_X1 g340(.A(new_n764), .B(new_n765), .C1(G129), .C2(new_n491), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  MUX2_X1   g342(.A(G32), .B(new_n767), .S(G29), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT27), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1996), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n743), .A2(new_n759), .A3(new_n761), .A4(new_n770), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n706), .A2(new_n730), .A3(new_n771), .ZN(new_n772));
  MUX2_X1   g347(.A(G6), .B(G305), .S(G16), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT89), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT32), .B(G1981), .Z(new_n775));
  OR2_X1    g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G16), .A2(G23), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT90), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G288), .B2(new_n701), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT33), .ZN(new_n780));
  INV_X1    g355(.A(G1976), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n701), .A2(G22), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G166), .B2(new_n701), .ZN(new_n784));
  INV_X1    g359(.A(G1971), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n774), .A2(new_n775), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n776), .A2(new_n782), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(KEYINPUT34), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(KEYINPUT34), .ZN(new_n790));
  MUX2_X1   g365(.A(G24), .B(G290), .S(G16), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1986), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n707), .A2(G25), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT88), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n486), .A2(G131), .ZN(new_n795));
  OAI21_X1  g370(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n796));
  INV_X1    g371(.A(G107), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(G2105), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n491), .B2(G119), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n794), .B1(new_n800), .B2(G29), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT35), .B(G1991), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n792), .A2(KEYINPUT91), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n789), .A2(new_n790), .A3(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT36), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n805), .A2(new_n806), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n772), .A2(new_n808), .A3(new_n809), .ZN(G150));
  INV_X1    g385(.A(G150), .ZN(G311));
  NAND2_X1  g386(.A1(new_n603), .A2(G559), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT38), .ZN(new_n813));
  NAND2_X1  g388(.A1(G80), .A2(G543), .ZN(new_n814));
  INV_X1    g389(.A(G67), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n511), .B2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT99), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n818), .A2(new_n819), .A3(new_n514), .ZN(new_n820));
  INV_X1    g395(.A(G55), .ZN(new_n821));
  INV_X1    g396(.A(G93), .ZN(new_n822));
  OAI22_X1  g397(.A1(new_n821), .A2(new_n521), .B1(new_n524), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n550), .B(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n813), .B(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT39), .ZN(new_n827));
  AOI21_X1  g402(.A(G860), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n827), .B2(new_n826), .ZN(new_n829));
  OAI21_X1  g404(.A(G860), .B1(new_n820), .B2(new_n823), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT37), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(G145));
  XNOR2_X1  g407(.A(new_n493), .B(new_n626), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT100), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(G160), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n800), .B(new_n618), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n697), .A2(KEYINPUT102), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n507), .A2(KEYINPUT101), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT101), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n505), .A2(new_n839), .A3(new_n506), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(new_n499), .A3(new_n840), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n837), .A2(new_n841), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n836), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n837), .A2(new_n841), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n837), .A2(new_n841), .ZN(new_n846));
  INV_X1    g421(.A(new_n836), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n716), .B(new_n767), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n491), .A2(G130), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n461), .A2(G118), .ZN(new_n852));
  OAI21_X1  g427(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n853));
  INV_X1    g428(.A(G142), .ZN(new_n854));
  OAI221_X1 g429(.A(new_n851), .B1(new_n852), .B2(new_n853), .C1(new_n624), .C2(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n850), .B(new_n855), .Z(new_n856));
  NAND2_X1  g431(.A1(new_n849), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n850), .B(new_n855), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n858), .A2(new_n848), .A3(new_n844), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n835), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(G37), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n857), .A2(new_n835), .A3(new_n859), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n862), .A2(new_n863), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g442(.A(G290), .B(G305), .ZN(new_n868));
  INV_X1    g443(.A(G288), .ZN(new_n869));
  XNOR2_X1  g444(.A(G303), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n868), .B(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT42), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n603), .A2(new_n825), .A3(new_n609), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n824), .B(new_n549), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n612), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n598), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(G299), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n598), .A2(new_n557), .A3(new_n561), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT104), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(new_n878), .B2(G299), .ZN(new_n883));
  XNOR2_X1  g458(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n884));
  NOR3_X1   g459(.A1(new_n881), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n879), .A2(new_n880), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n877), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n881), .A2(new_n883), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n890), .B(KEYINPUT105), .C1(new_n877), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n886), .A2(new_n882), .ZN(new_n893));
  INV_X1    g468(.A(new_n883), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n895), .A2(new_n896), .A3(new_n874), .A4(new_n876), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n873), .B1(new_n892), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n884), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n893), .A2(new_n894), .A3(new_n899), .ZN(new_n900));
  AOI22_X1  g475(.A1(new_n900), .A2(new_n888), .B1(new_n874), .B2(new_n876), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT105), .B1(new_n877), .B2(new_n891), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n897), .B(new_n873), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n872), .B1(new_n898), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n897), .B1(new_n901), .B2(new_n902), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT42), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(new_n871), .A3(new_n903), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n585), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n824), .A2(G868), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT107), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n907), .A2(new_n871), .A3(new_n903), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n871), .B1(new_n907), .B2(new_n903), .ZN(new_n913));
  OAI21_X1  g488(.A(G868), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n915));
  INV_X1    g490(.A(new_n910), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n911), .A2(new_n917), .ZN(G295));
  NAND2_X1  g493(.A1(new_n914), .A2(new_n916), .ZN(G331));
  AOI21_X1  g494(.A(G301), .B1(new_n564), .B2(new_n568), .ZN(new_n920));
  NOR2_X1   g495(.A1(G168), .A2(G171), .ZN(new_n921));
  OR3_X1    g496(.A1(new_n920), .A2(new_n825), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n825), .B1(new_n920), .B2(new_n921), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n895), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n925), .B(new_n884), .C1(new_n881), .C2(new_n883), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(new_n887), .B2(new_n886), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n925), .B1(new_n895), .B2(new_n884), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n923), .A2(KEYINPUT108), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n931), .B(new_n825), .C1(new_n920), .C2(new_n921), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n930), .A2(new_n922), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n924), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n871), .ZN(new_n935));
  INV_X1    g510(.A(new_n923), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n920), .A2(new_n825), .A3(new_n921), .ZN(new_n937));
  OAI22_X1  g512(.A1(new_n936), .A2(new_n937), .B1(new_n885), .B2(new_n889), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n930), .A2(new_n922), .A3(new_n895), .A4(new_n932), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n938), .A2(new_n939), .A3(new_n872), .A4(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n938), .A2(new_n939), .A3(new_n872), .ZN(new_n942));
  AOI21_X1  g517(.A(G37), .B1(new_n942), .B2(KEYINPUT109), .ZN(new_n943));
  AND4_X1   g518(.A1(KEYINPUT43), .A2(new_n935), .A3(new_n941), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(KEYINPUT109), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n939), .A2(new_n938), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n871), .ZN(new_n947));
  INV_X1    g522(.A(G37), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n945), .A2(new_n947), .A3(new_n948), .A4(new_n941), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT44), .B1(new_n944), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n935), .A2(new_n950), .A3(new_n941), .A4(new_n943), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n952), .A2(new_n957), .ZN(G397));
  INV_X1    g533(.A(G1384), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n495), .B1(new_n484), .B2(G138), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n840), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n839), .B1(new_n505), .B2(new_n506), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(G160), .A2(G40), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n716), .B(new_n719), .ZN(new_n969));
  INV_X1    g544(.A(G1996), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n767), .B(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n800), .B(new_n802), .Z(new_n974));
  OAI21_X1  g549(.A(new_n968), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(G290), .A2(G1986), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT111), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(G1986), .B2(G290), .ZN(new_n979));
  INV_X1    g554(.A(new_n968), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n975), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT112), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n509), .A2(new_n959), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n965), .ZN(new_n984));
  INV_X1    g559(.A(G40), .ZN(new_n985));
  AOI211_X1 g560(.A(new_n985), .B(new_n470), .C1(new_n472), .C2(new_n480), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n841), .A2(KEYINPUT45), .A3(new_n959), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n984), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(KEYINPUT56), .B(G2072), .Z(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT119), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT57), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n557), .A2(new_n992), .A3(new_n561), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n992), .B1(new_n557), .B2(new_n561), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n986), .B1(KEYINPUT50), .B2(new_n983), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n964), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n841), .A2(KEYINPUT113), .A3(new_n959), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n996), .B1(new_n1000), .B2(KEYINPUT50), .ZN(new_n1001));
  XNOR2_X1  g576(.A(KEYINPUT118), .B(G1956), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n991), .B(new_n995), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n1003), .A2(new_n878), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n998), .A2(new_n1005), .A3(new_n999), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1005), .B1(new_n509), .B2(new_n959), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n967), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT120), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1006), .A2(KEYINPUT120), .A3(new_n1008), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(new_n704), .A3(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n998), .A2(new_n999), .A3(new_n986), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1014), .A2(G2067), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n995), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n991), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n1004), .A2(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT58), .B(G1341), .Z(new_n1020));
  NAND2_X1  g595(.A1(new_n1014), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n984), .A2(new_n986), .A3(new_n987), .A4(new_n970), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n1021), .A2(KEYINPUT121), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT121), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n550), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT59), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT59), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1027), .B(new_n550), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n996), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n841), .A2(KEYINPUT113), .A3(new_n959), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT113), .B1(new_n841), .B2(new_n959), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT50), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1002), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n988), .A2(new_n990), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1017), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT123), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1036), .A2(new_n1003), .A3(new_n1037), .A4(KEYINPUT61), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1036), .A2(new_n1003), .A3(KEYINPUT122), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT61), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT122), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1018), .A2(new_n1041), .A3(new_n1017), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1036), .A2(new_n1003), .A3(KEYINPUT61), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT123), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1029), .A2(new_n1038), .A3(new_n1043), .A4(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT60), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n878), .B1(new_n1016), .B2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1013), .A2(KEYINPUT60), .A3(new_n598), .A4(new_n1015), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n1048), .A2(new_n1049), .B1(new_n1047), .B2(new_n1016), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1019), .B1(new_n1046), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1006), .A2(KEYINPUT120), .A3(new_n1008), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT120), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n1053), .A2(new_n1054), .A3(G1961), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n965), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1056));
  INV_X1    g631(.A(new_n983), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n967), .B1(KEYINPUT45), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1059), .A2(new_n1060), .A3(G2078), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT125), .B1(new_n1055), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G1961), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1011), .A2(new_n1063), .A3(new_n1012), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT125), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n986), .B1(new_n965), .B2(new_n983), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n1000), .B2(new_n965), .ZN(new_n1067));
  INV_X1    g642(.A(G2078), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(KEYINPUT53), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1064), .A2(new_n1065), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1062), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1060), .B1(new_n988), .B2(G2078), .ZN(new_n1072));
  AOI21_X1  g647(.A(G301), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n478), .A2(G2105), .ZN(new_n1074));
  NOR4_X1   g649(.A1(new_n470), .A2(new_n1060), .A3(new_n985), .A4(G2078), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n966), .A2(new_n1074), .A3(new_n987), .A4(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1064), .A2(new_n1072), .A3(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(G171), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1052), .B1(new_n1073), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT124), .ZN(new_n1080));
  INV_X1    g655(.A(G1966), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT45), .B1(new_n998), .B2(new_n999), .ZN(new_n1082));
  OAI211_X1 g657(.A(KEYINPUT117), .B(new_n1081), .C1(new_n1082), .C2(new_n1066), .ZN(new_n1083));
  INV_X1    g658(.A(G2084), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1006), .A2(new_n1084), .A3(new_n1008), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT117), .B1(new_n1059), .B2(new_n1081), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1080), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n1067), .B2(G1966), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1090), .A2(KEYINPUT124), .A3(new_n1085), .A4(new_n1083), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(new_n1091), .A3(G168), .ZN(new_n1092));
  AND2_X1   g667(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1090), .A2(new_n1085), .A3(new_n1083), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(G8), .ZN(new_n1096));
  INV_X1    g671(.A(G8), .ZN(new_n1097));
  NOR2_X1   g672(.A1(G168), .A2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1098), .A2(KEYINPUT51), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1094), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n1098), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n988), .A2(new_n785), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1009), .B2(G2090), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(G8), .ZN(new_n1107));
  NAND2_X1  g682(.A1(G303), .A2(G8), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(KEYINPUT55), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1014), .B(G8), .C1(new_n781), .C2(G288), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT52), .ZN(new_n1112));
  AND2_X1   g687(.A1(G305), .A2(G1981), .ZN(new_n1113));
  NOR2_X1   g688(.A1(G305), .A2(G1981), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT49), .ZN(new_n1115));
  OR3_X1    g690(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1115), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1116), .A2(new_n1117), .A3(G8), .A4(new_n1014), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT52), .B1(G288), .B2(new_n781), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1119), .B(KEYINPUT114), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1112), .B(new_n1118), .C1(new_n1111), .C2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1110), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1109), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1105), .B1(new_n1124), .B2(G2090), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1123), .B1(new_n1125), .B2(G8), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1071), .A2(G301), .A3(new_n1072), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1052), .B1(new_n1077), .B2(G171), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1051), .A2(new_n1079), .A3(new_n1104), .A4(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1101), .A2(new_n1133), .A3(new_n1103), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1092), .A2(new_n1093), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1102), .A2(new_n1098), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT62), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1126), .A2(new_n1110), .A3(new_n1121), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1138), .A2(new_n1139), .A3(G171), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1134), .A2(new_n1137), .A3(new_n1140), .A4(KEYINPUT126), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1096), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n569), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1142), .B1(new_n1128), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1142), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1122), .A2(new_n1143), .A3(new_n569), .A4(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1123), .A2(G8), .A3(new_n1106), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n1114), .B(KEYINPUT115), .Z(new_n1149));
  NOR2_X1   g724(.A1(G288), .A2(G1976), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n1118), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1014), .A2(G8), .ZN(new_n1152));
  OAI22_X1  g727(.A1(new_n1121), .A2(new_n1148), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT116), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1153), .A2(KEYINPUT116), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1145), .A2(new_n1147), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1132), .A2(new_n1141), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1073), .A2(new_n1139), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1158), .B1(new_n1104), .B2(KEYINPUT62), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT126), .B1(new_n1159), .B2(new_n1134), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n982), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n795), .A2(new_n802), .A3(new_n799), .ZN(new_n1162));
  OAI22_X1  g737(.A1(new_n973), .A2(new_n1162), .B1(G2067), .B2(new_n716), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1163), .A2(new_n968), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n767), .B1(KEYINPUT46), .B2(new_n970), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n969), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT46), .B1(new_n968), .B2(new_n970), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1167), .A2(KEYINPUT127), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1167), .A2(KEYINPUT127), .ZN(new_n1169));
  OAI22_X1  g744(.A1(new_n1166), .A2(new_n980), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n1170), .B(KEYINPUT47), .Z(new_n1171));
  NAND2_X1  g746(.A1(new_n978), .A2(new_n968), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT48), .ZN(new_n1173));
  AOI211_X1 g748(.A(new_n1164), .B(new_n1171), .C1(new_n975), .C2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1161), .A2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g750(.A1(G227), .A2(new_n459), .ZN(new_n1177));
  NAND3_X1  g751(.A1(new_n684), .A2(new_n685), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g752(.A(new_n1178), .B1(new_n646), .B2(new_n648), .ZN(new_n1179));
  NAND3_X1  g753(.A1(new_n1179), .A2(new_n955), .A3(new_n866), .ZN(G225));
  INV_X1    g754(.A(G225), .ZN(G308));
endmodule


