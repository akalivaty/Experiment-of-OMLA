

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775;

  AND2_X1 U372 ( .A1(n560), .A2(n571), .ZN(n569) );
  INV_X1 U373 ( .A(n548), .ZN(n710) );
  NOR2_X1 U374 ( .A1(n712), .A2(n711), .ZN(n706) );
  XNOR2_X1 U375 ( .A(n470), .B(n401), .ZN(n391) );
  NAND2_X1 U376 ( .A1(n689), .A2(n726), .ZN(n602) );
  INV_X1 U377 ( .A(G469), .ZN(n351) );
  XNOR2_X1 U378 ( .A(n481), .B(n480), .ZN(n390) );
  XNOR2_X1 U379 ( .A(n608), .B(KEYINPUT19), .ZN(n369) );
  INV_X1 U380 ( .A(G953), .ZN(n483) );
  NOR2_X2 U381 ( .A1(n646), .A2(n702), .ZN(n650) );
  XNOR2_X2 U382 ( .A(n393), .B(n424), .ZN(n761) );
  XNOR2_X2 U383 ( .A(n474), .B(G472), .ZN(n589) );
  BUF_X1 U384 ( .A(n560), .Z(n576) );
  AND2_X1 U385 ( .A1(n559), .A2(n681), .ZN(n571) );
  XNOR2_X1 U386 ( .A(n386), .B(n542), .ZN(n568) );
  OR2_X1 U387 ( .A1(n562), .A2(n550), .ZN(n552) );
  AND2_X1 U388 ( .A1(n623), .A2(n369), .ZN(n689) );
  OR2_X1 U389 ( .A1(n617), .A2(n721), .ZN(n619) );
  NOR2_X1 U390 ( .A1(n721), .A2(n720), .ZN(n621) );
  XNOR2_X1 U391 ( .A(n590), .B(KEYINPUT1), .ZN(n543) );
  OR2_X1 U392 ( .A1(n418), .A2(KEYINPUT93), .ZN(n356) );
  XNOR2_X1 U393 ( .A(n422), .B(n421), .ZN(n445) );
  XNOR2_X1 U394 ( .A(n425), .B(n423), .ZN(n422) );
  XOR2_X1 U395 ( .A(KEYINPUT59), .B(n670), .Z(n671) );
  XOR2_X1 U396 ( .A(KEYINPUT68), .B(n648), .Z(n649) );
  XNOR2_X1 U397 ( .A(KEYINPUT16), .B(G122), .ZN(n480) );
  INV_X1 U398 ( .A(KEYINPUT123), .ZN(n354) );
  XNOR2_X1 U399 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n485) );
  NOR2_X1 U400 ( .A1(G902), .A2(G237), .ZN(n475) );
  XNOR2_X1 U401 ( .A(G902), .B(KEYINPUT15), .ZN(n490) );
  INV_X1 U402 ( .A(KEYINPUT63), .ZN(n355) );
  BUF_X1 U403 ( .A(n676), .Z(n348) );
  XOR2_X1 U404 ( .A(n352), .B(n351), .Z(n349) );
  NOR2_X2 U405 ( .A1(n374), .A2(G902), .ZN(n352) );
  NAND2_X1 U406 ( .A1(n388), .A2(n387), .ZN(n386) );
  BUF_X1 U407 ( .A(n761), .Z(n350) );
  XNOR2_X2 U408 ( .A(n552), .B(n551), .ZN(n684) );
  XNOR2_X2 U409 ( .A(n352), .B(n351), .ZN(n590) );
  NAND2_X1 U410 ( .A1(n353), .A2(n570), .ZN(n578) );
  AND2_X1 U411 ( .A1(n577), .A2(n576), .ZN(n353) );
  NOR2_X2 U412 ( .A1(n658), .A2(n749), .ZN(n659) );
  BUF_X1 U413 ( .A(n651), .Z(n750) );
  NOR2_X2 U414 ( .A1(n664), .A2(n749), .ZN(n665) );
  XNOR2_X1 U415 ( .A(n659), .B(n354), .ZN(G63) );
  XNOR2_X1 U416 ( .A(n665), .B(n355), .ZN(G57) );
  AND2_X2 U417 ( .A1(n543), .A2(n706), .ZN(n561) );
  AND2_X1 U418 ( .A1(n590), .A2(n706), .ZN(n549) );
  AND2_X2 U419 ( .A1(n660), .A2(n568), .ZN(n577) );
  XNOR2_X2 U420 ( .A(n384), .B(n567), .ZN(n660) );
  NOR2_X1 U421 ( .A1(n720), .A2(n412), .ZN(n411) );
  OR2_X1 U422 ( .A1(n604), .A2(n383), .ZN(n381) );
  INV_X1 U423 ( .A(n699), .ZN(n382) );
  AND2_X1 U424 ( .A1(n367), .A2(KEYINPUT93), .ZN(n357) );
  NAND2_X1 U425 ( .A1(n411), .A2(n414), .ZN(n367) );
  NOR2_X1 U426 ( .A1(n406), .A2(n405), .ZN(n404) );
  INV_X1 U427 ( .A(G140), .ZN(n439) );
  INV_X1 U428 ( .A(KEYINPUT2), .ZN(n398) );
  XNOR2_X1 U429 ( .A(n370), .B(n629), .ZN(n399) );
  INV_X1 U430 ( .A(KEYINPUT28), .ZN(n427) );
  XNOR2_X1 U431 ( .A(n710), .B(n540), .ZN(n607) );
  NOR2_X1 U432 ( .A1(G953), .A2(G237), .ZN(n496) );
  XOR2_X1 U433 ( .A(KEYINPUT5), .B(G137), .Z(n472) );
  XNOR2_X1 U434 ( .A(G116), .B(G113), .ZN(n402) );
  XNOR2_X1 U435 ( .A(KEYINPUT79), .B(KEYINPUT98), .ZN(n441) );
  XNOR2_X1 U436 ( .A(G128), .B(KEYINPUT74), .ZN(n442) );
  XNOR2_X1 U437 ( .A(n436), .B(n435), .ZN(n519) );
  XNOR2_X1 U438 ( .A(n434), .B(n433), .ZN(n436) );
  XNOR2_X1 U439 ( .A(n486), .B(KEYINPUT10), .ZN(n760) );
  XNOR2_X1 U440 ( .A(n510), .B(n509), .ZN(n555) );
  XNOR2_X1 U441 ( .A(n508), .B(G475), .ZN(n509) );
  NAND2_X1 U442 ( .A1(n416), .A2(n415), .ZN(n414) );
  INV_X1 U443 ( .A(n647), .ZN(n415) );
  INV_X1 U444 ( .A(n411), .ZN(n406) );
  NOR2_X1 U445 ( .A1(n493), .A2(n408), .ZN(n405) );
  INV_X1 U446 ( .A(n490), .ZN(n647) );
  INV_X1 U447 ( .A(KEYINPUT72), .ZN(n371) );
  NAND2_X1 U448 ( .A1(n493), .A2(n647), .ZN(n417) );
  XNOR2_X1 U449 ( .A(G116), .B(G107), .ZN(n511) );
  NAND2_X1 U450 ( .A1(G237), .A2(G234), .ZN(n462) );
  AND2_X1 U451 ( .A1(n469), .A2(n468), .ZN(n395) );
  NAND2_X1 U452 ( .A1(n368), .A2(n357), .ZN(n409) );
  INV_X1 U453 ( .A(G902), .ZN(n444) );
  NAND2_X1 U454 ( .A1(n399), .A2(n419), .ZN(n702) );
  XNOR2_X1 U455 ( .A(G143), .B(G122), .ZN(n503) );
  XOR2_X1 U456 ( .A(G140), .B(G104), .Z(n504) );
  XNOR2_X1 U457 ( .A(n481), .B(n460), .ZN(n461) );
  XOR2_X1 U458 ( .A(G101), .B(G146), .Z(n459) );
  NOR2_X1 U459 ( .A1(n645), .A2(n398), .ZN(n397) );
  AND2_X1 U460 ( .A1(n429), .A2(n426), .ZN(n623) );
  XNOR2_X1 U461 ( .A(n428), .B(n427), .ZN(n426) );
  XNOR2_X1 U462 ( .A(n549), .B(KEYINPUT112), .ZN(n469) );
  XNOR2_X1 U463 ( .A(n431), .B(n482), .ZN(n430) );
  XNOR2_X1 U464 ( .A(n473), .B(n471), .ZN(n431) );
  BUF_X1 U465 ( .A(n483), .Z(n767) );
  XNOR2_X1 U466 ( .A(n702), .B(n375), .ZN(n768) );
  INV_X1 U467 ( .A(n766), .ZN(n375) );
  XNOR2_X1 U468 ( .A(n760), .B(n443), .ZN(n421) );
  XNOR2_X1 U469 ( .A(n636), .B(n635), .ZN(n638) );
  XNOR2_X1 U470 ( .A(n634), .B(n633), .ZN(n635) );
  AND2_X1 U471 ( .A1(n541), .A2(n557), .ZN(n387) );
  XNOR2_X1 U472 ( .A(n348), .B(n675), .ZN(n677) );
  INV_X1 U473 ( .A(n645), .ZN(n419) );
  NAND2_X1 U474 ( .A1(n644), .A2(n771), .ZN(n645) );
  NOR2_X1 U475 ( .A1(n707), .A2(n710), .ZN(n358) );
  AND2_X1 U476 ( .A1(n558), .A2(n557), .ZN(n359) );
  AND2_X1 U477 ( .A1(n413), .A2(n417), .ZN(n360) );
  AND2_X1 U478 ( .A1(n381), .A2(n382), .ZN(n361) );
  NAND2_X1 U479 ( .A1(n604), .A2(n383), .ZN(n362) );
  XOR2_X1 U480 ( .A(n534), .B(KEYINPUT67), .Z(n363) );
  XOR2_X1 U481 ( .A(n580), .B(KEYINPUT45), .Z(n364) );
  INV_X1 U482 ( .A(KEYINPUT76), .ZN(n383) );
  XNOR2_X2 U483 ( .A(n547), .B(n546), .ZN(n696) );
  BUF_X1 U484 ( .A(n561), .Z(n365) );
  BUF_X1 U485 ( .A(n374), .Z(n366) );
  XNOR2_X1 U486 ( .A(n761), .B(n461), .ZN(n374) );
  BUF_X1 U487 ( .A(n666), .Z(n743) );
  OR2_X1 U488 ( .A1(n676), .A2(n414), .ZN(n413) );
  NAND2_X1 U489 ( .A1(n676), .A2(n411), .ZN(n368) );
  XNOR2_X2 U490 ( .A(n389), .B(n755), .ZN(n676) );
  NAND2_X1 U491 ( .A1(n388), .A2(n358), .ZN(n537) );
  NAND2_X1 U492 ( .A1(n388), .A2(n359), .ZN(n681) );
  XNOR2_X2 U493 ( .A(n535), .B(n363), .ZN(n388) );
  NAND2_X1 U494 ( .A1(n369), .A2(n529), .ZN(n530) );
  XNOR2_X1 U495 ( .A(n372), .B(n371), .ZN(n420) );
  NAND2_X1 U496 ( .A1(n628), .A2(n420), .ZN(n370) );
  NAND2_X1 U497 ( .A1(n376), .A2(n361), .ZN(n372) );
  NAND2_X2 U498 ( .A1(n373), .A2(n356), .ZN(n608) );
  NAND2_X1 U499 ( .A1(n410), .A2(n409), .ZN(n373) );
  XNOR2_X1 U500 ( .A(n366), .B(KEYINPUT122), .ZN(n744) );
  NAND2_X1 U501 ( .A1(n378), .A2(n377), .ZN(n376) );
  NAND2_X1 U502 ( .A1(n380), .A2(n362), .ZN(n377) );
  NAND2_X1 U503 ( .A1(n379), .A2(n383), .ZN(n378) );
  INV_X1 U504 ( .A(n380), .ZN(n379) );
  XNOR2_X2 U505 ( .A(n600), .B(n599), .ZN(n380) );
  NAND2_X1 U506 ( .A1(n385), .A2(n566), .ZN(n384) );
  XNOR2_X1 U507 ( .A(n565), .B(n564), .ZN(n385) );
  XNOR2_X1 U508 ( .A(n489), .B(n488), .ZN(n389) );
  XNOR2_X2 U509 ( .A(n517), .B(n455), .ZN(n489) );
  XNOR2_X2 U510 ( .A(n454), .B(G143), .ZN(n517) );
  XNOR2_X2 U511 ( .A(n482), .B(n390), .ZN(n755) );
  XNOR2_X2 U512 ( .A(n400), .B(G110), .ZN(n481) );
  XNOR2_X2 U513 ( .A(n391), .B(n402), .ZN(n482) );
  XNOR2_X2 U514 ( .A(n392), .B(KEYINPUT33), .ZN(n563) );
  NAND2_X1 U515 ( .A1(n561), .A2(n607), .ZN(n392) );
  XNOR2_X1 U516 ( .A(n393), .B(n430), .ZN(n661) );
  XNOR2_X2 U517 ( .A(n489), .B(n456), .ZN(n393) );
  NAND2_X1 U518 ( .A1(n394), .A2(n469), .ZN(n495) );
  AND2_X1 U519 ( .A1(n494), .A2(n468), .ZN(n394) );
  NAND2_X1 U520 ( .A1(n395), .A2(n614), .ZN(n617) );
  NAND2_X1 U521 ( .A1(n399), .A2(n397), .ZN(n396) );
  XNOR2_X1 U522 ( .A(n396), .B(KEYINPUT86), .ZN(n652) );
  XNOR2_X2 U523 ( .A(G107), .B(G104), .ZN(n400) );
  XNOR2_X2 U524 ( .A(G101), .B(KEYINPUT94), .ZN(n401) );
  NAND2_X1 U525 ( .A1(n676), .A2(n493), .ZN(n418) );
  NAND2_X1 U526 ( .A1(n403), .A2(n413), .ZN(n410) );
  AND2_X2 U527 ( .A1(n407), .A2(n404), .ZN(n403) );
  OR2_X2 U528 ( .A1(n676), .A2(n408), .ZN(n407) );
  INV_X1 U529 ( .A(KEYINPUT93), .ZN(n408) );
  NAND2_X1 U530 ( .A1(n360), .A2(n418), .ZN(n616) );
  INV_X1 U531 ( .A(n417), .ZN(n412) );
  INV_X1 U532 ( .A(n493), .ZN(n416) );
  XNOR2_X2 U533 ( .A(n451), .B(n450), .ZN(n712) );
  INV_X1 U534 ( .A(n445), .ZN(n667) );
  XNOR2_X1 U535 ( .A(n440), .B(n424), .ZN(n423) );
  INV_X1 U536 ( .A(n457), .ZN(n424) );
  NAND2_X1 U537 ( .A1(n519), .A2(G221), .ZN(n425) );
  NAND2_X1 U538 ( .A1(n588), .A2(n589), .ZN(n428) );
  INV_X1 U539 ( .A(n349), .ZN(n429) );
  AND2_X1 U540 ( .A1(n724), .A2(n532), .ZN(n432) );
  INV_X1 U541 ( .A(KEYINPUT11), .ZN(n499) );
  XNOR2_X1 U542 ( .A(n472), .B(G146), .ZN(n473) );
  XNOR2_X1 U543 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U544 ( .A(n502), .B(n501), .ZN(n507) );
  INV_X1 U545 ( .A(KEYINPUT110), .ZN(n633) );
  AND2_X1 U546 ( .A1(n614), .A2(n637), .ZN(n494) );
  INV_X1 U547 ( .A(KEYINPUT34), .ZN(n564) );
  NAND2_X1 U548 ( .A1(n483), .A2(G234), .ZN(n434) );
  INV_X1 U549 ( .A(KEYINPUT71), .ZN(n433) );
  XOR2_X1 U550 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n435) );
  XNOR2_X1 U551 ( .A(G119), .B(G110), .ZN(n438) );
  XNOR2_X1 U552 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n437) );
  XNOR2_X1 U553 ( .A(n438), .B(n437), .ZN(n440) );
  XNOR2_X1 U554 ( .A(n439), .B(G137), .ZN(n457) );
  XNOR2_X1 U555 ( .A(G146), .B(G125), .ZN(n486) );
  XNOR2_X1 U556 ( .A(n442), .B(n441), .ZN(n443) );
  NAND2_X1 U557 ( .A1(n445), .A2(n444), .ZN(n451) );
  XOR2_X1 U558 ( .A(KEYINPUT100), .B(KEYINPUT20), .Z(n447) );
  NAND2_X1 U559 ( .A1(G234), .A2(n490), .ZN(n446) );
  XNOR2_X1 U560 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U561 ( .A(n448), .B(KEYINPUT99), .ZN(n452) );
  NAND2_X1 U562 ( .A1(n452), .A2(G217), .ZN(n449) );
  XNOR2_X1 U563 ( .A(n449), .B(KEYINPUT25), .ZN(n450) );
  NAND2_X1 U564 ( .A1(n452), .A2(G221), .ZN(n453) );
  XNOR2_X1 U565 ( .A(n453), .B(KEYINPUT21), .ZN(n711) );
  XNOR2_X2 U566 ( .A(G128), .B(KEYINPUT65), .ZN(n454) );
  INV_X1 U567 ( .A(KEYINPUT4), .ZN(n455) );
  XNOR2_X1 U568 ( .A(G134), .B(G131), .ZN(n456) );
  NAND2_X1 U569 ( .A1(G227), .A2(n767), .ZN(n458) );
  XNOR2_X1 U570 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U571 ( .A(n462), .B(KEYINPUT14), .ZN(n463) );
  NAND2_X1 U572 ( .A1(G952), .A2(n463), .ZN(n734) );
  NOR2_X1 U573 ( .A1(G953), .A2(n734), .ZN(n527) );
  AND2_X1 U574 ( .A1(G902), .A2(n463), .ZN(n524) );
  NAND2_X1 U575 ( .A1(G953), .A2(n524), .ZN(n464) );
  NOR2_X1 U576 ( .A1(G900), .A2(n464), .ZN(n465) );
  NOR2_X1 U577 ( .A1(n527), .A2(n465), .ZN(n467) );
  INV_X1 U578 ( .A(KEYINPUT81), .ZN(n466) );
  XNOR2_X1 U579 ( .A(n467), .B(n466), .ZN(n585) );
  INV_X1 U580 ( .A(n585), .ZN(n468) );
  XNOR2_X2 U581 ( .A(KEYINPUT3), .B(G119), .ZN(n470) );
  NAND2_X1 U582 ( .A1(n496), .A2(G210), .ZN(n471) );
  NAND2_X1 U583 ( .A1(n661), .A2(n444), .ZN(n474) );
  XNOR2_X1 U584 ( .A(n475), .B(KEYINPUT78), .ZN(n492) );
  INV_X1 U585 ( .A(G214), .ZN(n476) );
  OR2_X1 U586 ( .A1(n492), .A2(n476), .ZN(n477) );
  XNOR2_X1 U587 ( .A(n477), .B(KEYINPUT95), .ZN(n720) );
  INV_X1 U588 ( .A(n720), .ZN(n478) );
  AND2_X1 U589 ( .A1(n589), .A2(n478), .ZN(n479) );
  XNOR2_X1 U590 ( .A(n479), .B(KEYINPUT30), .ZN(n614) );
  NAND2_X1 U591 ( .A1(n483), .A2(G224), .ZN(n484) );
  XNOR2_X1 U592 ( .A(n485), .B(n484), .ZN(n487) );
  XNOR2_X1 U593 ( .A(n487), .B(n486), .ZN(n488) );
  INV_X1 U594 ( .A(G210), .ZN(n491) );
  OR2_X1 U595 ( .A1(n492), .A2(n491), .ZN(n493) );
  INV_X1 U596 ( .A(n616), .ZN(n637) );
  XNOR2_X1 U597 ( .A(n495), .B(KEYINPUT113), .ZN(n523) );
  XOR2_X1 U598 ( .A(KEYINPUT12), .B(KEYINPUT102), .Z(n498) );
  NAND2_X1 U599 ( .A1(G214), .A2(n496), .ZN(n497) );
  XNOR2_X1 U600 ( .A(n498), .B(n497), .ZN(n502) );
  XNOR2_X1 U601 ( .A(G113), .B(G131), .ZN(n500) );
  XNOR2_X1 U602 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U603 ( .A(n760), .B(n505), .ZN(n506) );
  XNOR2_X1 U604 ( .A(n507), .B(n506), .ZN(n670) );
  NOR2_X1 U605 ( .A1(G902), .A2(n670), .ZN(n510) );
  XNOR2_X1 U606 ( .A(KEYINPUT103), .B(KEYINPUT13), .ZN(n508) );
  XOR2_X1 U607 ( .A(G134), .B(G122), .Z(n512) );
  XNOR2_X1 U608 ( .A(n512), .B(n511), .ZN(n516) );
  XOR2_X1 U609 ( .A(KEYINPUT9), .B(KEYINPUT105), .Z(n514) );
  XNOR2_X1 U610 ( .A(KEYINPUT7), .B(KEYINPUT104), .ZN(n513) );
  XNOR2_X1 U611 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U612 ( .A(n516), .B(n515), .Z(n518) );
  XNOR2_X1 U613 ( .A(n517), .B(n518), .ZN(n521) );
  NAND2_X1 U614 ( .A1(n519), .A2(G217), .ZN(n520) );
  XNOR2_X1 U615 ( .A(n521), .B(n520), .ZN(n654) );
  NAND2_X1 U616 ( .A1(n654), .A2(n444), .ZN(n522) );
  XNOR2_X1 U617 ( .A(n522), .B(G478), .ZN(n554) );
  INV_X1 U618 ( .A(n554), .ZN(n531) );
  NOR2_X1 U619 ( .A1(n555), .A2(n531), .ZN(n566) );
  NAND2_X1 U620 ( .A1(n523), .A2(n566), .ZN(n584) );
  XNOR2_X1 U621 ( .A(n584), .B(G143), .ZN(G45) );
  NOR2_X1 U622 ( .A1(G898), .A2(n767), .ZN(n756) );
  NAND2_X1 U623 ( .A1(n524), .A2(n756), .ZN(n525) );
  XOR2_X1 U624 ( .A(KEYINPUT96), .B(n525), .Z(n526) );
  NOR2_X1 U625 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U626 ( .A(n528), .B(KEYINPUT97), .ZN(n529) );
  XNOR2_X2 U627 ( .A(n530), .B(KEYINPUT0), .ZN(n562) );
  INV_X1 U628 ( .A(n562), .ZN(n533) );
  AND2_X1 U629 ( .A1(n555), .A2(n531), .ZN(n724) );
  INV_X1 U630 ( .A(n711), .ZN(n532) );
  NAND2_X1 U631 ( .A1(n533), .A2(n432), .ZN(n535) );
  XNOR2_X1 U632 ( .A(KEYINPUT75), .B(KEYINPUT22), .ZN(n534) );
  BUF_X1 U633 ( .A(n543), .Z(n707) );
  INV_X1 U634 ( .A(n589), .ZN(n548) );
  INV_X1 U635 ( .A(KEYINPUT66), .ZN(n536) );
  XNOR2_X1 U636 ( .A(n537), .B(n536), .ZN(n538) );
  NAND2_X1 U637 ( .A1(n538), .A2(n712), .ZN(n560) );
  XNOR2_X1 U638 ( .A(n576), .B(G110), .ZN(G12) );
  NAND2_X1 U639 ( .A1(n707), .A2(n712), .ZN(n539) );
  XNOR2_X1 U640 ( .A(n539), .B(KEYINPUT107), .ZN(n541) );
  INV_X1 U641 ( .A(KEYINPUT6), .ZN(n540) );
  INV_X1 U642 ( .A(n607), .ZN(n557) );
  XNOR2_X1 U643 ( .A(KEYINPUT80), .B(KEYINPUT32), .ZN(n542) );
  XNOR2_X1 U644 ( .A(n568), .B(G119), .ZN(G21) );
  NAND2_X1 U645 ( .A1(n365), .A2(n710), .ZN(n717) );
  INV_X1 U646 ( .A(n717), .ZN(n545) );
  INV_X1 U647 ( .A(n562), .ZN(n544) );
  NAND2_X1 U648 ( .A1(n545), .A2(n544), .ZN(n547) );
  INV_X1 U649 ( .A(KEYINPUT31), .ZN(n546) );
  NAND2_X1 U650 ( .A1(n549), .A2(n548), .ZN(n550) );
  INV_X1 U651 ( .A(KEYINPUT101), .ZN(n551) );
  NAND2_X1 U652 ( .A1(n696), .A2(n684), .ZN(n556) );
  NAND2_X1 U653 ( .A1(n555), .A2(n554), .ZN(n553) );
  XNOR2_X1 U654 ( .A(n553), .B(KEYINPUT106), .ZN(n640) );
  OR2_X1 U655 ( .A1(n555), .A2(n554), .ZN(n694) );
  NAND2_X1 U656 ( .A1(n640), .A2(n694), .ZN(n726) );
  NAND2_X1 U657 ( .A1(n556), .A2(n726), .ZN(n559) );
  NOR2_X1 U658 ( .A1(n707), .A2(n712), .ZN(n558) );
  NAND2_X1 U659 ( .A1(n563), .A2(n544), .ZN(n565) );
  XNOR2_X1 U660 ( .A(KEYINPUT87), .B(KEYINPUT35), .ZN(n567) );
  NAND2_X1 U661 ( .A1(n577), .A2(n569), .ZN(n573) );
  INV_X1 U662 ( .A(KEYINPUT44), .ZN(n570) );
  NAND2_X1 U663 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U664 ( .A1(n573), .A2(n572), .ZN(n575) );
  INV_X1 U665 ( .A(KEYINPUT91), .ZN(n574) );
  XNOR2_X1 U666 ( .A(n575), .B(n574), .ZN(n579) );
  NAND2_X1 U667 ( .A1(n579), .A2(n578), .ZN(n581) );
  INV_X1 U668 ( .A(KEYINPUT64), .ZN(n580) );
  XNOR2_X2 U669 ( .A(n581), .B(n364), .ZN(n651) );
  NAND2_X1 U670 ( .A1(n651), .A2(n647), .ZN(n583) );
  INV_X1 U671 ( .A(KEYINPUT85), .ZN(n582) );
  XNOR2_X1 U672 ( .A(n583), .B(n582), .ZN(n646) );
  XNOR2_X1 U673 ( .A(n584), .B(KEYINPUT84), .ZN(n598) );
  OR2_X1 U674 ( .A1(n585), .A2(n711), .ZN(n586) );
  XNOR2_X1 U675 ( .A(n586), .B(KEYINPUT73), .ZN(n587) );
  NAND2_X1 U676 ( .A1(n587), .A2(n712), .ZN(n605) );
  INV_X1 U677 ( .A(n605), .ZN(n588) );
  NAND2_X1 U678 ( .A1(n602), .A2(KEYINPUT47), .ZN(n592) );
  INV_X1 U679 ( .A(KEYINPUT83), .ZN(n591) );
  NAND2_X1 U680 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U681 ( .A1(KEYINPUT83), .A2(KEYINPUT47), .ZN(n593) );
  NOR2_X1 U682 ( .A1(n726), .A2(n593), .ZN(n594) );
  NAND2_X1 U683 ( .A1(n689), .A2(n594), .ZN(n595) );
  NAND2_X1 U684 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U685 ( .A1(n598), .A2(n597), .ZN(n600) );
  INV_X1 U686 ( .A(KEYINPUT82), .ZN(n599) );
  XOR2_X1 U687 ( .A(KEYINPUT47), .B(KEYINPUT69), .Z(n601) );
  NOR2_X1 U688 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U689 ( .A(n603), .B(KEYINPUT77), .ZN(n604) );
  NOR2_X1 U690 ( .A1(n694), .A2(n605), .ZN(n606) );
  NAND2_X1 U691 ( .A1(n607), .A2(n606), .ZN(n630) );
  BUF_X1 U692 ( .A(n608), .Z(n609) );
  NOR2_X1 U693 ( .A1(n630), .A2(n609), .ZN(n611) );
  XOR2_X1 U694 ( .A(KEYINPUT92), .B(KEYINPUT36), .Z(n610) );
  XNOR2_X1 U695 ( .A(n611), .B(n610), .ZN(n613) );
  INV_X1 U696 ( .A(n707), .ZN(n612) );
  NOR2_X1 U697 ( .A1(n613), .A2(n612), .ZN(n699) );
  INV_X1 U698 ( .A(KEYINPUT38), .ZN(n615) );
  XNOR2_X1 U699 ( .A(n616), .B(n615), .ZN(n721) );
  XOR2_X1 U700 ( .A(KEYINPUT90), .B(KEYINPUT39), .Z(n618) );
  XNOR2_X1 U701 ( .A(n619), .B(n618), .ZN(n641) );
  NOR2_X1 U702 ( .A1(n694), .A2(n641), .ZN(n620) );
  XNOR2_X1 U703 ( .A(n620), .B(KEYINPUT40), .ZN(n774) );
  XOR2_X1 U704 ( .A(KEYINPUT114), .B(KEYINPUT42), .Z(n625) );
  NAND2_X1 U705 ( .A1(n621), .A2(n724), .ZN(n622) );
  XNOR2_X1 U706 ( .A(n622), .B(KEYINPUT41), .ZN(n737) );
  NAND2_X1 U707 ( .A1(n623), .A2(n737), .ZN(n624) );
  XNOR2_X1 U708 ( .A(n625), .B(n624), .ZN(n773) );
  NOR2_X1 U709 ( .A1(n774), .A2(n773), .ZN(n627) );
  XOR2_X1 U710 ( .A(KEYINPUT89), .B(KEYINPUT46), .Z(n626) );
  XNOR2_X1 U711 ( .A(n627), .B(n626), .ZN(n628) );
  XOR2_X1 U712 ( .A(KEYINPUT88), .B(KEYINPUT48), .Z(n629) );
  NOR2_X1 U713 ( .A1(n720), .A2(n630), .ZN(n631) );
  XOR2_X1 U714 ( .A(KEYINPUT108), .B(n631), .Z(n632) );
  NOR2_X1 U715 ( .A1(n707), .A2(n632), .ZN(n636) );
  XNOR2_X1 U716 ( .A(KEYINPUT43), .B(KEYINPUT109), .ZN(n634) );
  NOR2_X1 U717 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U718 ( .A(KEYINPUT111), .B(n639), .Z(n772) );
  INV_X1 U719 ( .A(n772), .ZN(n644) );
  OR2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n643) );
  INV_X1 U721 ( .A(KEYINPUT115), .ZN(n642) );
  XNOR2_X1 U722 ( .A(n643), .B(n642), .ZN(n771) );
  NAND2_X1 U723 ( .A1(n647), .A2(KEYINPUT2), .ZN(n648) );
  NOR2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n653) );
  INV_X1 U725 ( .A(n750), .ZN(n701) );
  NOR2_X1 U726 ( .A1(n652), .A2(n701), .ZN(n705) );
  NOR2_X2 U727 ( .A1(n653), .A2(n705), .ZN(n666) );
  NAND2_X1 U728 ( .A1(n666), .A2(G478), .ZN(n656) );
  INV_X1 U729 ( .A(n654), .ZN(n655) );
  XNOR2_X1 U730 ( .A(n656), .B(n655), .ZN(n658) );
  INV_X1 U731 ( .A(G952), .ZN(n657) );
  AND2_X1 U732 ( .A1(n657), .A2(G953), .ZN(n749) );
  XNOR2_X1 U733 ( .A(n660), .B(G122), .ZN(G24) );
  NAND2_X1 U734 ( .A1(n666), .A2(G472), .ZN(n663) );
  XOR2_X1 U735 ( .A(KEYINPUT62), .B(n661), .Z(n662) );
  XNOR2_X1 U736 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U737 ( .A1(n743), .A2(G217), .ZN(n668) );
  XNOR2_X1 U738 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X1 U739 ( .A1(n669), .A2(n749), .ZN(G66) );
  NAND2_X1 U740 ( .A1(n666), .A2(G475), .ZN(n672) );
  XNOR2_X1 U741 ( .A(n672), .B(n671), .ZN(n673) );
  NOR2_X2 U742 ( .A1(n673), .A2(n749), .ZN(n674) );
  XNOR2_X1 U743 ( .A(n674), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U744 ( .A1(n666), .A2(G210), .ZN(n678) );
  XOR2_X1 U745 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n675) );
  XNOR2_X1 U746 ( .A(n678), .B(n677), .ZN(n679) );
  NOR2_X2 U747 ( .A1(n679), .A2(n749), .ZN(n680) );
  XNOR2_X1 U748 ( .A(n680), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U749 ( .A(n681), .B(G101), .ZN(n682) );
  XNOR2_X1 U750 ( .A(KEYINPUT116), .B(n682), .ZN(G3) );
  NOR2_X1 U751 ( .A1(n694), .A2(n684), .ZN(n683) );
  XOR2_X1 U752 ( .A(G104), .B(n683), .Z(G6) );
  NOR2_X1 U753 ( .A1(n684), .A2(n640), .ZN(n688) );
  XOR2_X1 U754 ( .A(KEYINPUT27), .B(KEYINPUT117), .Z(n686) );
  XNOR2_X1 U755 ( .A(G107), .B(KEYINPUT26), .ZN(n685) );
  XNOR2_X1 U756 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U757 ( .A(n688), .B(n687), .ZN(G9) );
  INV_X1 U758 ( .A(n689), .ZN(n692) );
  NOR2_X1 U759 ( .A1(n692), .A2(n640), .ZN(n691) );
  XNOR2_X1 U760 ( .A(G128), .B(KEYINPUT29), .ZN(n690) );
  XNOR2_X1 U761 ( .A(n691), .B(n690), .ZN(G30) );
  NOR2_X1 U762 ( .A1(n692), .A2(n694), .ZN(n693) );
  XOR2_X1 U763 ( .A(G146), .B(n693), .Z(G48) );
  NOR2_X1 U764 ( .A1(n694), .A2(n696), .ZN(n695) );
  XOR2_X1 U765 ( .A(G113), .B(n695), .Z(G15) );
  NOR2_X1 U766 ( .A1(n640), .A2(n696), .ZN(n697) );
  XOR2_X1 U767 ( .A(KEYINPUT118), .B(n697), .Z(n698) );
  XNOR2_X1 U768 ( .A(G116), .B(n698), .ZN(G18) );
  XNOR2_X1 U769 ( .A(G125), .B(n699), .ZN(n700) );
  XNOR2_X1 U770 ( .A(n700), .B(KEYINPUT37), .ZN(G27) );
  NOR2_X1 U771 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U772 ( .A1(n703), .A2(KEYINPUT2), .ZN(n704) );
  NOR2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n736) );
  NOR2_X1 U774 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U775 ( .A(n708), .B(KEYINPUT50), .ZN(n709) );
  NOR2_X1 U776 ( .A1(n710), .A2(n709), .ZN(n715) );
  NAND2_X1 U777 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U778 ( .A(KEYINPUT49), .B(n713), .Z(n714) );
  NAND2_X1 U779 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U780 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U781 ( .A(KEYINPUT51), .B(n718), .Z(n719) );
  NAND2_X1 U782 ( .A1(n737), .A2(n719), .ZN(n731) );
  NAND2_X1 U783 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U784 ( .A(KEYINPUT119), .B(n722), .Z(n723) );
  NAND2_X1 U785 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U786 ( .A(n725), .B(KEYINPUT120), .ZN(n728) );
  NAND2_X1 U787 ( .A1(n621), .A2(n726), .ZN(n727) );
  NAND2_X1 U788 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U789 ( .A1(n563), .A2(n729), .ZN(n730) );
  NAND2_X1 U790 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U791 ( .A(KEYINPUT52), .B(n732), .Z(n733) );
  NOR2_X1 U792 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U793 ( .A1(n736), .A2(n735), .ZN(n740) );
  AND2_X1 U794 ( .A1(n563), .A2(n737), .ZN(n738) );
  XNOR2_X1 U795 ( .A(n738), .B(KEYINPUT121), .ZN(n739) );
  NAND2_X1 U796 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U797 ( .A1(n741), .A2(G953), .ZN(n742) );
  XNOR2_X1 U798 ( .A(n742), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U799 ( .A1(n743), .A2(G469), .ZN(n747) );
  XOR2_X1 U800 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n745) );
  XNOR2_X1 U801 ( .A(n745), .B(n744), .ZN(n746) );
  XNOR2_X1 U802 ( .A(n747), .B(n746), .ZN(n748) );
  NOR2_X1 U803 ( .A1(n749), .A2(n748), .ZN(G54) );
  NAND2_X1 U804 ( .A1(n750), .A2(n767), .ZN(n754) );
  NAND2_X1 U805 ( .A1(G953), .A2(G224), .ZN(n751) );
  XNOR2_X1 U806 ( .A(KEYINPUT61), .B(n751), .ZN(n752) );
  NAND2_X1 U807 ( .A1(n752), .A2(G898), .ZN(n753) );
  NAND2_X1 U808 ( .A1(n754), .A2(n753), .ZN(n759) );
  XNOR2_X1 U809 ( .A(n755), .B(KEYINPUT124), .ZN(n757) );
  NOR2_X1 U810 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U811 ( .A(n759), .B(n758), .ZN(G69) );
  XNOR2_X1 U812 ( .A(n350), .B(n760), .ZN(n766) );
  XOR2_X1 U813 ( .A(G227), .B(n766), .Z(n762) );
  NAND2_X1 U814 ( .A1(n762), .A2(G900), .ZN(n763) );
  XOR2_X1 U815 ( .A(KEYINPUT125), .B(n763), .Z(n764) );
  NAND2_X1 U816 ( .A1(G953), .A2(n764), .ZN(n765) );
  XNOR2_X1 U817 ( .A(n765), .B(KEYINPUT126), .ZN(n770) );
  NAND2_X1 U818 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U819 ( .A1(n770), .A2(n769), .ZN(G72) );
  XNOR2_X1 U820 ( .A(G134), .B(n771), .ZN(G36) );
  XOR2_X1 U821 ( .A(n772), .B(G140), .Z(G42) );
  XOR2_X1 U822 ( .A(G137), .B(n773), .Z(G39) );
  XNOR2_X1 U823 ( .A(G131), .B(KEYINPUT127), .ZN(n775) );
  XNOR2_X1 U824 ( .A(n775), .B(n774), .ZN(G33) );
endmodule

