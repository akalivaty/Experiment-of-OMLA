

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U551 ( .A(KEYINPUT66), .B(n535), .ZN(n872) );
  NOR2_X1 U552 ( .A1(G168), .A2(n518), .ZN(n703) );
  NOR2_X2 U553 ( .A1(n785), .A2(n787), .ZN(n517) );
  XOR2_X1 U554 ( .A(KEYINPUT99), .B(n699), .Z(n518) );
  INV_X1 U555 ( .A(KEYINPUT100), .ZN(n704) );
  XNOR2_X1 U556 ( .A(n704), .B(KEYINPUT31), .ZN(n705) );
  NOR2_X1 U557 ( .A1(n703), .A2(n702), .ZN(n706) );
  XNOR2_X1 U558 ( .A(n706), .B(n705), .ZN(n749) );
  NAND2_X1 U559 ( .A1(n757), .A2(n756), .ZN(n805) );
  INV_X1 U560 ( .A(KEYINPUT64), .ZN(n689) );
  NOR2_X1 U561 ( .A1(G164), .A2(G1384), .ZN(n690) );
  XNOR2_X1 U562 ( .A(n690), .B(n689), .ZN(n785) );
  XNOR2_X1 U563 ( .A(n536), .B(KEYINPUT65), .ZN(n547) );
  BUF_X1 U564 ( .A(n547), .Z(n865) );
  NOR2_X1 U565 ( .A1(G651), .A2(n637), .ZN(n657) );
  AND2_X1 U566 ( .A1(n544), .A2(n543), .ZN(G164) );
  NOR2_X1 U567 ( .A1(G651), .A2(G543), .ZN(n651) );
  NAND2_X1 U568 ( .A1(n651), .A2(G89), .ZN(n519) );
  XNOR2_X1 U569 ( .A(n519), .B(KEYINPUT4), .ZN(n521) );
  XOR2_X1 U570 ( .A(G543), .B(KEYINPUT0), .Z(n637) );
  INV_X1 U571 ( .A(G651), .ZN(n524) );
  NOR2_X1 U572 ( .A1(n637), .A2(n524), .ZN(n652) );
  NAND2_X1 U573 ( .A1(G76), .A2(n652), .ZN(n520) );
  NAND2_X1 U574 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U575 ( .A(KEYINPUT5), .B(n522), .ZN(n532) );
  XNOR2_X1 U576 ( .A(KEYINPUT77), .B(KEYINPUT78), .ZN(n530) );
  NAND2_X1 U577 ( .A1(n657), .A2(G51), .ZN(n523) );
  XNOR2_X1 U578 ( .A(n523), .B(KEYINPUT76), .ZN(n527) );
  NOR2_X1 U579 ( .A1(G543), .A2(n524), .ZN(n525) );
  XOR2_X1 U580 ( .A(KEYINPUT1), .B(n525), .Z(n656) );
  NAND2_X1 U581 ( .A1(G63), .A2(n656), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U583 ( .A(n528), .B(KEYINPUT6), .ZN(n529) );
  XNOR2_X1 U584 ( .A(n530), .B(n529), .ZN(n531) );
  NAND2_X1 U585 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U586 ( .A(KEYINPUT7), .B(n533), .ZN(G168) );
  NOR2_X1 U587 ( .A1(G2105), .A2(G2104), .ZN(n534) );
  XOR2_X1 U588 ( .A(n534), .B(KEYINPUT17), .Z(n535) );
  NAND2_X1 U589 ( .A1(n872), .A2(G138), .ZN(n544) );
  NAND2_X1 U590 ( .A1(G2104), .A2(G2105), .ZN(n536) );
  NAND2_X1 U591 ( .A1(G114), .A2(n547), .ZN(n537) );
  XNOR2_X1 U592 ( .A(n537), .B(KEYINPUT88), .ZN(n539) );
  INV_X1 U593 ( .A(G2104), .ZN(n540) );
  AND2_X1 U594 ( .A1(n540), .A2(G2105), .ZN(n864) );
  NAND2_X1 U595 ( .A1(n864), .A2(G126), .ZN(n538) );
  AND2_X1 U596 ( .A1(n539), .A2(n538), .ZN(n542) );
  NOR2_X1 U597 ( .A1(G2105), .A2(n540), .ZN(n869) );
  NAND2_X1 U598 ( .A1(n869), .A2(G102), .ZN(n541) );
  AND2_X1 U599 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U600 ( .A1(G101), .A2(n869), .ZN(n545) );
  XOR2_X1 U601 ( .A(KEYINPUT23), .B(n545), .Z(n691) );
  NAND2_X1 U602 ( .A1(G137), .A2(n872), .ZN(n546) );
  XOR2_X1 U603 ( .A(KEYINPUT67), .B(n546), .Z(n551) );
  NAND2_X1 U604 ( .A1(G125), .A2(n864), .ZN(n549) );
  NAND2_X1 U605 ( .A1(G113), .A2(n865), .ZN(n548) );
  AND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(n550) );
  AND2_X1 U607 ( .A1(n551), .A2(n550), .ZN(n692) );
  AND2_X1 U608 ( .A1(n691), .A2(n692), .ZN(G160) );
  XOR2_X1 U609 ( .A(G2446), .B(G2430), .Z(n553) );
  XNOR2_X1 U610 ( .A(G2451), .B(G2454), .ZN(n552) );
  XNOR2_X1 U611 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U612 ( .A(n554), .B(G2427), .Z(n556) );
  XNOR2_X1 U613 ( .A(G1341), .B(G1348), .ZN(n555) );
  XNOR2_X1 U614 ( .A(n556), .B(n555), .ZN(n560) );
  XOR2_X1 U615 ( .A(G2443), .B(KEYINPUT104), .Z(n558) );
  XNOR2_X1 U616 ( .A(G2438), .B(G2435), .ZN(n557) );
  XNOR2_X1 U617 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U618 ( .A(n560), .B(n559), .Z(n561) );
  AND2_X1 U619 ( .A1(G14), .A2(n561), .ZN(G401) );
  AND2_X1 U620 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U621 ( .A1(n872), .A2(G135), .ZN(n562) );
  XNOR2_X1 U622 ( .A(n562), .B(KEYINPUT80), .ZN(n569) );
  NAND2_X1 U623 ( .A1(G99), .A2(n869), .ZN(n564) );
  NAND2_X1 U624 ( .A1(G111), .A2(n865), .ZN(n563) );
  NAND2_X1 U625 ( .A1(n564), .A2(n563), .ZN(n567) );
  NAND2_X1 U626 ( .A1(n864), .A2(G123), .ZN(n565) );
  XOR2_X1 U627 ( .A(KEYINPUT18), .B(n565), .Z(n566) );
  NOR2_X1 U628 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(n997) );
  XNOR2_X1 U630 ( .A(G2096), .B(n997), .ZN(n570) );
  OR2_X1 U631 ( .A1(G2100), .A2(n570), .ZN(G156) );
  INV_X1 U632 ( .A(G57), .ZN(G237) );
  INV_X1 U633 ( .A(G132), .ZN(G219) );
  INV_X1 U634 ( .A(G82), .ZN(G220) );
  XOR2_X1 U635 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U636 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n572) );
  NAND2_X1 U637 ( .A1(G7), .A2(G661), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G223) );
  INV_X1 U639 ( .A(G223), .ZN(n836) );
  NAND2_X1 U640 ( .A1(n836), .A2(G567), .ZN(n573) );
  XOR2_X1 U641 ( .A(KEYINPUT11), .B(n573), .Z(G234) );
  XOR2_X1 U642 ( .A(KEYINPUT12), .B(KEYINPUT72), .Z(n575) );
  NAND2_X1 U643 ( .A1(G81), .A2(n651), .ZN(n574) );
  XNOR2_X1 U644 ( .A(n575), .B(n574), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n652), .A2(G68), .ZN(n576) );
  XNOR2_X1 U646 ( .A(KEYINPUT73), .B(n576), .ZN(n577) );
  NOR2_X1 U647 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U648 ( .A(KEYINPUT74), .B(KEYINPUT13), .ZN(n579) );
  XNOR2_X1 U649 ( .A(n580), .B(n579), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n656), .A2(G56), .ZN(n581) );
  XOR2_X1 U651 ( .A(KEYINPUT14), .B(n581), .Z(n582) );
  NOR2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n657), .A2(G43), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n949) );
  INV_X1 U655 ( .A(G860), .ZN(n613) );
  OR2_X1 U656 ( .A1(n949), .A2(n613), .ZN(G153) );
  NAND2_X1 U657 ( .A1(G64), .A2(n656), .ZN(n586) );
  XNOR2_X1 U658 ( .A(n586), .B(KEYINPUT69), .ZN(n591) );
  NAND2_X1 U659 ( .A1(G90), .A2(n651), .ZN(n588) );
  NAND2_X1 U660 ( .A1(G77), .A2(n652), .ZN(n587) );
  NAND2_X1 U661 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U662 ( .A(KEYINPUT9), .B(n589), .Z(n590) );
  NOR2_X1 U663 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n657), .A2(G52), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n593), .A2(n592), .ZN(G301) );
  NAND2_X1 U666 ( .A1(G868), .A2(G301), .ZN(n603) );
  NAND2_X1 U667 ( .A1(G66), .A2(n656), .ZN(n600) );
  NAND2_X1 U668 ( .A1(G92), .A2(n651), .ZN(n595) );
  NAND2_X1 U669 ( .A1(G79), .A2(n652), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U671 ( .A1(G54), .A2(n657), .ZN(n596) );
  XNOR2_X1 U672 ( .A(KEYINPUT75), .B(n596), .ZN(n597) );
  NOR2_X1 U673 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U675 ( .A(n601), .B(KEYINPUT15), .ZN(n888) );
  INV_X1 U676 ( .A(n888), .ZN(n941) );
  INV_X1 U677 ( .A(G868), .ZN(n670) );
  NAND2_X1 U678 ( .A1(n941), .A2(n670), .ZN(n602) );
  NAND2_X1 U679 ( .A1(n603), .A2(n602), .ZN(G284) );
  NAND2_X1 U680 ( .A1(G91), .A2(n651), .ZN(n605) );
  NAND2_X1 U681 ( .A1(G78), .A2(n652), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U683 ( .A1(n657), .A2(G53), .ZN(n606) );
  XOR2_X1 U684 ( .A(KEYINPUT70), .B(n606), .Z(n607) );
  NOR2_X1 U685 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n656), .A2(G65), .ZN(n609) );
  NAND2_X1 U687 ( .A1(n610), .A2(n609), .ZN(G299) );
  NOR2_X1 U688 ( .A1(G286), .A2(n670), .ZN(n612) );
  NOR2_X1 U689 ( .A1(G868), .A2(G299), .ZN(n611) );
  NOR2_X1 U690 ( .A1(n612), .A2(n611), .ZN(G297) );
  NAND2_X1 U691 ( .A1(n613), .A2(G559), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n614), .A2(n888), .ZN(n615) );
  XNOR2_X1 U693 ( .A(n615), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U694 ( .A1(G868), .A2(n949), .ZN(n616) );
  XOR2_X1 U695 ( .A(KEYINPUT79), .B(n616), .Z(n619) );
  NAND2_X1 U696 ( .A1(G868), .A2(n888), .ZN(n617) );
  NOR2_X1 U697 ( .A1(G559), .A2(n617), .ZN(n618) );
  NOR2_X1 U698 ( .A1(n619), .A2(n618), .ZN(G282) );
  NAND2_X1 U699 ( .A1(n888), .A2(G559), .ZN(n668) );
  XNOR2_X1 U700 ( .A(n949), .B(n668), .ZN(n620) );
  NOR2_X1 U701 ( .A1(n620), .A2(G860), .ZN(n628) );
  NAND2_X1 U702 ( .A1(G67), .A2(n656), .ZN(n622) );
  NAND2_X1 U703 ( .A1(G55), .A2(n657), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n627) );
  NAND2_X1 U705 ( .A1(G93), .A2(n651), .ZN(n624) );
  NAND2_X1 U706 ( .A1(G80), .A2(n652), .ZN(n623) );
  NAND2_X1 U707 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U708 ( .A(KEYINPUT81), .B(n625), .Z(n626) );
  OR2_X1 U709 ( .A1(n627), .A2(n626), .ZN(n671) );
  XOR2_X1 U710 ( .A(n628), .B(n671), .Z(G145) );
  NAND2_X1 U711 ( .A1(G73), .A2(n652), .ZN(n629) );
  XNOR2_X1 U712 ( .A(n629), .B(KEYINPUT2), .ZN(n636) );
  NAND2_X1 U713 ( .A1(G86), .A2(n651), .ZN(n631) );
  NAND2_X1 U714 ( .A1(G61), .A2(n656), .ZN(n630) );
  NAND2_X1 U715 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U716 ( .A1(G48), .A2(n657), .ZN(n632) );
  XNOR2_X1 U717 ( .A(KEYINPUT83), .B(n632), .ZN(n633) );
  NOR2_X1 U718 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n636), .A2(n635), .ZN(G305) );
  NAND2_X1 U720 ( .A1(G74), .A2(G651), .ZN(n642) );
  NAND2_X1 U721 ( .A1(G49), .A2(n657), .ZN(n639) );
  NAND2_X1 U722 ( .A1(G87), .A2(n637), .ZN(n638) );
  NAND2_X1 U723 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U724 ( .A1(n656), .A2(n640), .ZN(n641) );
  NAND2_X1 U725 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U726 ( .A(n643), .B(KEYINPUT82), .ZN(G288) );
  NAND2_X1 U727 ( .A1(G88), .A2(n651), .ZN(n645) );
  NAND2_X1 U728 ( .A1(G75), .A2(n652), .ZN(n644) );
  NAND2_X1 U729 ( .A1(n645), .A2(n644), .ZN(n650) );
  NAND2_X1 U730 ( .A1(G50), .A2(n657), .ZN(n646) );
  XNOR2_X1 U731 ( .A(n646), .B(KEYINPUT84), .ZN(n648) );
  NAND2_X1 U732 ( .A1(n656), .A2(G62), .ZN(n647) );
  NAND2_X1 U733 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U734 ( .A1(n650), .A2(n649), .ZN(G166) );
  NAND2_X1 U735 ( .A1(G85), .A2(n651), .ZN(n654) );
  NAND2_X1 U736 ( .A1(G72), .A2(n652), .ZN(n653) );
  NAND2_X1 U737 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U738 ( .A(KEYINPUT68), .B(n655), .Z(n661) );
  NAND2_X1 U739 ( .A1(G60), .A2(n656), .ZN(n659) );
  NAND2_X1 U740 ( .A1(G47), .A2(n657), .ZN(n658) );
  AND2_X1 U741 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U742 ( .A1(n661), .A2(n660), .ZN(G290) );
  INV_X1 U743 ( .A(G299), .ZN(n944) );
  XNOR2_X1 U744 ( .A(n944), .B(G305), .ZN(n667) );
  XOR2_X1 U745 ( .A(KEYINPUT19), .B(n671), .Z(n663) );
  XNOR2_X1 U746 ( .A(n949), .B(G166), .ZN(n662) );
  XNOR2_X1 U747 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U748 ( .A(G288), .B(n664), .ZN(n665) );
  XNOR2_X1 U749 ( .A(n665), .B(G290), .ZN(n666) );
  XNOR2_X1 U750 ( .A(n667), .B(n666), .ZN(n887) );
  XNOR2_X1 U751 ( .A(n887), .B(n668), .ZN(n669) );
  NOR2_X1 U752 ( .A1(n670), .A2(n669), .ZN(n673) );
  NOR2_X1 U753 ( .A1(G868), .A2(n671), .ZN(n672) );
  NOR2_X1 U754 ( .A1(n673), .A2(n672), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2084), .A2(G2078), .ZN(n674) );
  XNOR2_X1 U756 ( .A(n674), .B(KEYINPUT85), .ZN(n675) );
  XNOR2_X1 U757 ( .A(n675), .B(KEYINPUT20), .ZN(n676) );
  NAND2_X1 U758 ( .A1(n676), .A2(G2090), .ZN(n677) );
  XNOR2_X1 U759 ( .A(n677), .B(KEYINPUT21), .ZN(n678) );
  XNOR2_X1 U760 ( .A(n678), .B(KEYINPUT86), .ZN(n679) );
  NAND2_X1 U761 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U763 ( .A1(G220), .A2(G219), .ZN(n680) );
  XOR2_X1 U764 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U765 ( .A1(G218), .A2(n681), .ZN(n682) );
  NAND2_X1 U766 ( .A1(G96), .A2(n682), .ZN(n840) );
  NAND2_X1 U767 ( .A1(n840), .A2(G2106), .ZN(n686) );
  NAND2_X1 U768 ( .A1(G69), .A2(G120), .ZN(n683) );
  NOR2_X1 U769 ( .A1(G237), .A2(n683), .ZN(n684) );
  NAND2_X1 U770 ( .A1(G108), .A2(n684), .ZN(n841) );
  NAND2_X1 U771 ( .A1(n841), .A2(G567), .ZN(n685) );
  NAND2_X1 U772 ( .A1(n686), .A2(n685), .ZN(n917) );
  NAND2_X1 U773 ( .A1(G483), .A2(G661), .ZN(n687) );
  NOR2_X1 U774 ( .A1(n917), .A2(n687), .ZN(n688) );
  XOR2_X1 U775 ( .A(KEYINPUT87), .B(n688), .Z(n839) );
  NAND2_X1 U776 ( .A1(n839), .A2(G36), .ZN(G176) );
  XNOR2_X1 U777 ( .A(KEYINPUT89), .B(G166), .ZN(G303) );
  INV_X1 U778 ( .A(G301), .ZN(G171) );
  AND2_X1 U779 ( .A1(n691), .A2(G40), .ZN(n693) );
  NAND2_X1 U780 ( .A1(n693), .A2(n692), .ZN(n787) );
  NOR2_X1 U781 ( .A1(n517), .A2(G1966), .ZN(n694) );
  NAND2_X1 U782 ( .A1(n694), .A2(G8), .ZN(n697) );
  INV_X1 U783 ( .A(n697), .ZN(n737) );
  INV_X1 U784 ( .A(G2084), .ZN(n738) );
  NAND2_X1 U785 ( .A1(n738), .A2(n517), .ZN(n695) );
  AND2_X1 U786 ( .A1(n695), .A2(G8), .ZN(n696) );
  NAND2_X1 U787 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U788 ( .A(KEYINPUT30), .B(n698), .ZN(n699) );
  INV_X1 U789 ( .A(n517), .ZN(n743) );
  XNOR2_X1 U790 ( .A(G2078), .B(KEYINPUT25), .ZN(n926) );
  NOR2_X1 U791 ( .A1(n743), .A2(n926), .ZN(n701) );
  AND2_X1 U792 ( .A1(n743), .A2(G1961), .ZN(n700) );
  NOR2_X1 U793 ( .A1(n701), .A2(n700), .ZN(n707) );
  NOR2_X1 U794 ( .A1(G171), .A2(n707), .ZN(n702) );
  NAND2_X1 U795 ( .A1(n707), .A2(G171), .ZN(n735) );
  NAND2_X1 U796 ( .A1(n517), .A2(G2072), .ZN(n708) );
  XNOR2_X1 U797 ( .A(n708), .B(KEYINPUT27), .ZN(n710) );
  AND2_X1 U798 ( .A1(G1956), .A2(n743), .ZN(n709) );
  NOR2_X1 U799 ( .A1(n710), .A2(n709), .ZN(n712) );
  NOR2_X1 U800 ( .A1(n944), .A2(n712), .ZN(n711) );
  XOR2_X1 U801 ( .A(n711), .B(KEYINPUT28), .Z(n732) );
  NAND2_X1 U802 ( .A1(n944), .A2(n712), .ZN(n730) );
  NAND2_X1 U803 ( .A1(G2067), .A2(n517), .ZN(n714) );
  NAND2_X1 U804 ( .A1(G1348), .A2(n743), .ZN(n713) );
  NAND2_X1 U805 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U806 ( .A1(n715), .A2(n941), .ZN(n728) );
  OR2_X1 U807 ( .A1(n715), .A2(n941), .ZN(n726) );
  INV_X1 U808 ( .A(G1341), .ZN(n970) );
  NOR2_X1 U809 ( .A1(n517), .A2(n970), .ZN(n719) );
  AND2_X1 U810 ( .A1(n719), .A2(KEYINPUT26), .ZN(n716) );
  NOR2_X1 U811 ( .A1(KEYINPUT98), .A2(n716), .ZN(n717) );
  NOR2_X1 U812 ( .A1(n949), .A2(n717), .ZN(n724) );
  NAND2_X1 U813 ( .A1(n517), .A2(G1996), .ZN(n718) );
  XNOR2_X1 U814 ( .A(KEYINPUT26), .B(n718), .ZN(n721) );
  INV_X1 U815 ( .A(n719), .ZN(n720) );
  NAND2_X1 U816 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U817 ( .A1(KEYINPUT98), .A2(n722), .ZN(n723) );
  NAND2_X1 U818 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U819 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U820 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U821 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U822 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U823 ( .A(KEYINPUT29), .B(n733), .Z(n734) );
  NAND2_X1 U824 ( .A1(n735), .A2(n734), .ZN(n747) );
  AND2_X1 U825 ( .A1(n749), .A2(n747), .ZN(n736) );
  NOR2_X1 U826 ( .A1(n737), .A2(n736), .ZN(n742) );
  AND2_X1 U827 ( .A1(n738), .A2(n517), .ZN(n739) );
  NAND2_X1 U828 ( .A1(G8), .A2(n739), .ZN(n740) );
  XOR2_X1 U829 ( .A(KEYINPUT97), .B(n740), .Z(n741) );
  NAND2_X1 U830 ( .A1(n742), .A2(n741), .ZN(n757) );
  NAND2_X1 U831 ( .A1(G8), .A2(n743), .ZN(n810) );
  NOR2_X1 U832 ( .A1(G1971), .A2(n810), .ZN(n745) );
  NOR2_X1 U833 ( .A1(G2090), .A2(n743), .ZN(n744) );
  NOR2_X1 U834 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n746), .A2(G303), .ZN(n750) );
  AND2_X1 U836 ( .A1(n747), .A2(n750), .ZN(n748) );
  NAND2_X1 U837 ( .A1(n749), .A2(n748), .ZN(n754) );
  INV_X1 U838 ( .A(n750), .ZN(n751) );
  OR2_X1 U839 ( .A1(n751), .A2(G286), .ZN(n752) );
  AND2_X1 U840 ( .A1(n752), .A2(G8), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U842 ( .A(n755), .B(KEYINPUT32), .ZN(n756) );
  NOR2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n938) );
  NOR2_X1 U844 ( .A1(G1971), .A2(G303), .ZN(n758) );
  NOR2_X1 U845 ( .A1(n938), .A2(n758), .ZN(n759) );
  NAND2_X1 U846 ( .A1(n805), .A2(n759), .ZN(n761) );
  NAND2_X1 U847 ( .A1(G288), .A2(G1976), .ZN(n760) );
  XOR2_X1 U848 ( .A(KEYINPUT101), .B(n760), .Z(n939) );
  NAND2_X1 U849 ( .A1(n761), .A2(n939), .ZN(n762) );
  NOR2_X1 U850 ( .A1(n762), .A2(n810), .ZN(n763) );
  NOR2_X1 U851 ( .A1(KEYINPUT33), .A2(n763), .ZN(n766) );
  NAND2_X1 U852 ( .A1(n938), .A2(KEYINPUT33), .ZN(n764) );
  NOR2_X1 U853 ( .A1(n764), .A2(n810), .ZN(n765) );
  NOR2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n802) );
  XOR2_X1 U855 ( .A(G1981), .B(G305), .Z(n958) );
  XOR2_X1 U856 ( .A(KEYINPUT92), .B(KEYINPUT38), .Z(n768) );
  NAND2_X1 U857 ( .A1(G105), .A2(n869), .ZN(n767) );
  XNOR2_X1 U858 ( .A(n768), .B(n767), .ZN(n772) );
  NAND2_X1 U859 ( .A1(G129), .A2(n864), .ZN(n770) );
  NAND2_X1 U860 ( .A1(G117), .A2(n865), .ZN(n769) );
  NAND2_X1 U861 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U862 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U863 ( .A(KEYINPUT93), .B(n773), .Z(n775) );
  NAND2_X1 U864 ( .A1(G141), .A2(n872), .ZN(n774) );
  NAND2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n850) );
  NAND2_X1 U866 ( .A1(n850), .A2(G1996), .ZN(n784) );
  NAND2_X1 U867 ( .A1(G95), .A2(n869), .ZN(n777) );
  NAND2_X1 U868 ( .A1(G119), .A2(n864), .ZN(n776) );
  NAND2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U870 ( .A1(G131), .A2(n872), .ZN(n778) );
  XNOR2_X1 U871 ( .A(KEYINPUT91), .B(n778), .ZN(n779) );
  NOR2_X1 U872 ( .A1(n780), .A2(n779), .ZN(n782) );
  NAND2_X1 U873 ( .A1(n865), .A2(G107), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n877) );
  NAND2_X1 U875 ( .A1(n877), .A2(G1991), .ZN(n783) );
  AND2_X1 U876 ( .A1(n784), .A2(n783), .ZN(n1002) );
  INV_X1 U877 ( .A(n785), .ZN(n786) );
  NOR2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n818) );
  XOR2_X1 U879 ( .A(n818), .B(KEYINPUT94), .Z(n788) );
  NOR2_X1 U880 ( .A1(n1002), .A2(n788), .ZN(n824) );
  XNOR2_X1 U881 ( .A(KEYINPUT95), .B(n824), .ZN(n800) );
  INV_X1 U882 ( .A(n818), .ZN(n831) );
  NAND2_X1 U883 ( .A1(G128), .A2(n864), .ZN(n790) );
  NAND2_X1 U884 ( .A1(G116), .A2(n865), .ZN(n789) );
  NAND2_X1 U885 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U886 ( .A(KEYINPUT35), .B(n791), .ZN(n797) );
  NAND2_X1 U887 ( .A1(n869), .A2(G104), .ZN(n792) );
  XNOR2_X1 U888 ( .A(n792), .B(KEYINPUT90), .ZN(n794) );
  NAND2_X1 U889 ( .A1(G140), .A2(n872), .ZN(n793) );
  NAND2_X1 U890 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U891 ( .A(KEYINPUT34), .B(n795), .Z(n796) );
  NAND2_X1 U892 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U893 ( .A(KEYINPUT36), .B(n798), .ZN(n883) );
  XOR2_X1 U894 ( .A(KEYINPUT37), .B(G2067), .Z(n821) );
  NAND2_X1 U895 ( .A1(n883), .A2(n821), .ZN(n1015) );
  NOR2_X1 U896 ( .A1(n831), .A2(n1015), .ZN(n828) );
  INV_X1 U897 ( .A(n828), .ZN(n799) );
  AND2_X1 U898 ( .A1(n800), .A2(n799), .ZN(n814) );
  AND2_X1 U899 ( .A1(n958), .A2(n814), .ZN(n801) );
  NAND2_X1 U900 ( .A1(n802), .A2(n801), .ZN(n816) );
  NOR2_X1 U901 ( .A1(G2090), .A2(G303), .ZN(n803) );
  NAND2_X1 U902 ( .A1(G8), .A2(n803), .ZN(n804) );
  NAND2_X1 U903 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U904 ( .A1(n806), .A2(n810), .ZN(n812) );
  NOR2_X1 U905 ( .A1(G1981), .A2(G305), .ZN(n807) );
  XOR2_X1 U906 ( .A(n807), .B(KEYINPUT96), .Z(n808) );
  XNOR2_X1 U907 ( .A(KEYINPUT24), .B(n808), .ZN(n809) );
  OR2_X1 U908 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U909 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U912 ( .A(n817), .B(KEYINPUT102), .ZN(n820) );
  XNOR2_X1 U913 ( .A(G1986), .B(G290), .ZN(n943) );
  NAND2_X1 U914 ( .A1(n943), .A2(n818), .ZN(n819) );
  NAND2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n834) );
  NOR2_X1 U916 ( .A1(n883), .A2(n821), .ZN(n1018) );
  NOR2_X1 U917 ( .A1(G1996), .A2(n850), .ZN(n1009) );
  NOR2_X1 U918 ( .A1(G1986), .A2(G290), .ZN(n822) );
  NOR2_X1 U919 ( .A1(G1991), .A2(n877), .ZN(n1000) );
  NOR2_X1 U920 ( .A1(n822), .A2(n1000), .ZN(n823) );
  NOR2_X1 U921 ( .A1(n824), .A2(n823), .ZN(n825) );
  NOR2_X1 U922 ( .A1(n1009), .A2(n825), .ZN(n826) );
  XOR2_X1 U923 ( .A(KEYINPUT39), .B(n826), .Z(n827) );
  NOR2_X1 U924 ( .A1(n828), .A2(n827), .ZN(n829) );
  NOR2_X1 U925 ( .A1(n1018), .A2(n829), .ZN(n830) );
  NOR2_X1 U926 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U927 ( .A(KEYINPUT103), .B(n832), .ZN(n833) );
  NAND2_X1 U928 ( .A1(n834), .A2(n833), .ZN(n835) );
  XNOR2_X1 U929 ( .A(n835), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n836), .ZN(G217) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U932 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U934 ( .A1(n839), .A2(n838), .ZN(G188) );
  NOR2_X1 U935 ( .A1(n841), .A2(n840), .ZN(G325) );
  XNOR2_X1 U936 ( .A(KEYINPUT105), .B(G325), .ZN(G261) );
  INV_X1 U938 ( .A(G120), .ZN(G236) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  INV_X1 U940 ( .A(G69), .ZN(G235) );
  NAND2_X1 U941 ( .A1(G124), .A2(n864), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n842), .B(KEYINPUT44), .ZN(n845) );
  NAND2_X1 U943 ( .A1(G100), .A2(n869), .ZN(n843) );
  XOR2_X1 U944 ( .A(KEYINPUT107), .B(n843), .Z(n844) );
  NAND2_X1 U945 ( .A1(n845), .A2(n844), .ZN(n849) );
  NAND2_X1 U946 ( .A1(n865), .A2(G112), .ZN(n847) );
  NAND2_X1 U947 ( .A1(G136), .A2(n872), .ZN(n846) );
  NAND2_X1 U948 ( .A1(n847), .A2(n846), .ZN(n848) );
  NOR2_X1 U949 ( .A1(n849), .A2(n848), .ZN(G162) );
  XNOR2_X1 U950 ( .A(G164), .B(n850), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n851), .B(n997), .ZN(n863) );
  NAND2_X1 U952 ( .A1(G130), .A2(n864), .ZN(n853) );
  NAND2_X1 U953 ( .A1(G118), .A2(n865), .ZN(n852) );
  NAND2_X1 U954 ( .A1(n853), .A2(n852), .ZN(n861) );
  NAND2_X1 U955 ( .A1(G142), .A2(n872), .ZN(n854) );
  XNOR2_X1 U956 ( .A(KEYINPUT109), .B(n854), .ZN(n857) );
  NAND2_X1 U957 ( .A1(n869), .A2(G106), .ZN(n855) );
  XOR2_X1 U958 ( .A(n855), .B(KEYINPUT108), .Z(n856) );
  NOR2_X1 U959 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U960 ( .A(KEYINPUT110), .B(n858), .Z(n859) );
  XOR2_X1 U961 ( .A(n859), .B(KEYINPUT45), .Z(n860) );
  NOR2_X1 U962 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U963 ( .A(n863), .B(n862), .Z(n879) );
  NAND2_X1 U964 ( .A1(G127), .A2(n864), .ZN(n867) );
  NAND2_X1 U965 ( .A1(G115), .A2(n865), .ZN(n866) );
  NAND2_X1 U966 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n868), .B(KEYINPUT47), .ZN(n871) );
  NAND2_X1 U968 ( .A1(G103), .A2(n869), .ZN(n870) );
  NAND2_X1 U969 ( .A1(n871), .A2(n870), .ZN(n875) );
  NAND2_X1 U970 ( .A1(G139), .A2(n872), .ZN(n873) );
  XNOR2_X1 U971 ( .A(KEYINPUT111), .B(n873), .ZN(n874) );
  NOR2_X1 U972 ( .A1(n875), .A2(n874), .ZN(n1004) );
  XOR2_X1 U973 ( .A(G160), .B(n1004), .Z(n876) );
  XNOR2_X1 U974 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U975 ( .A(n879), .B(n878), .Z(n885) );
  XOR2_X1 U976 ( .A(KEYINPUT48), .B(KEYINPUT112), .Z(n881) );
  XNOR2_X1 U977 ( .A(G162), .B(KEYINPUT46), .ZN(n880) );
  XNOR2_X1 U978 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U979 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U980 ( .A(n885), .B(n884), .ZN(n886) );
  NOR2_X1 U981 ( .A1(G37), .A2(n886), .ZN(G395) );
  XOR2_X1 U982 ( .A(n887), .B(G286), .Z(n890) );
  XNOR2_X1 U983 ( .A(G171), .B(n888), .ZN(n889) );
  XNOR2_X1 U984 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U985 ( .A1(G37), .A2(n891), .ZN(G397) );
  XOR2_X1 U986 ( .A(G1976), .B(G1981), .Z(n893) );
  XNOR2_X1 U987 ( .A(G1966), .B(G1971), .ZN(n892) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U989 ( .A(n894), .B(KEYINPUT41), .Z(n896) );
  XNOR2_X1 U990 ( .A(G1996), .B(G1991), .ZN(n895) );
  XNOR2_X1 U991 ( .A(n896), .B(n895), .ZN(n900) );
  XOR2_X1 U992 ( .A(G2474), .B(G1956), .Z(n898) );
  XNOR2_X1 U993 ( .A(G1986), .B(G1961), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(G229) );
  XOR2_X1 U996 ( .A(G2096), .B(KEYINPUT43), .Z(n902) );
  XNOR2_X1 U997 ( .A(G2072), .B(G2678), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U999 ( .A(n903), .B(KEYINPUT42), .Z(n905) );
  XNOR2_X1 U1000 ( .A(G2067), .B(G2090), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n909) );
  XOR2_X1 U1002 ( .A(KEYINPUT106), .B(G2100), .Z(n907) );
  XNOR2_X1 U1003 ( .A(G2084), .B(G2078), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(G227) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(KEYINPUT114), .B(n910), .ZN(n916) );
  NOR2_X1 U1008 ( .A1(n917), .A2(G401), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n911), .B(KEYINPUT113), .ZN(n914) );
  NOR2_X1 U1010 ( .A1(G229), .A2(G227), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n912), .ZN(n913) );
  NOR2_X1 U1012 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(n917), .ZN(G319) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1017 ( .A(G2084), .B(G34), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(n918), .B(KEYINPUT54), .ZN(n934) );
  XNOR2_X1 U1019 ( .A(G2090), .B(G35), .ZN(n931) );
  XNOR2_X1 U1020 ( .A(G1996), .B(G32), .ZN(n920) );
  XNOR2_X1 U1021 ( .A(G33), .B(G2072), .ZN(n919) );
  NOR2_X1 U1022 ( .A1(n920), .A2(n919), .ZN(n925) );
  XOR2_X1 U1023 ( .A(G1991), .B(G25), .Z(n921) );
  NAND2_X1 U1024 ( .A1(n921), .A2(G28), .ZN(n923) );
  XNOR2_X1 U1025 ( .A(G26), .B(G2067), .ZN(n922) );
  NOR2_X1 U1026 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1027 ( .A1(n925), .A2(n924), .ZN(n928) );
  XOR2_X1 U1028 ( .A(G27), .B(n926), .Z(n927) );
  NOR2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(KEYINPUT53), .B(n929), .ZN(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1032 ( .A(KEYINPUT118), .B(n932), .Z(n933) );
  NOR2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1034 ( .A(KEYINPUT55), .B(n935), .Z(n936) );
  NOR2_X1 U1035 ( .A1(G29), .A2(n936), .ZN(n937) );
  XOR2_X1 U1036 ( .A(KEYINPUT119), .B(n937), .Z(n995) );
  XNOR2_X1 U1037 ( .A(KEYINPUT121), .B(n938), .ZN(n940) );
  NAND2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n956) );
  XNOR2_X1 U1039 ( .A(G1348), .B(n941), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n954) );
  XNOR2_X1 U1041 ( .A(n944), .B(G1956), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(G301), .B(G1961), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(G303), .B(G1971), .ZN(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G1341), .B(n949), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(KEYINPUT122), .B(n950), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(KEYINPUT123), .B(n957), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(G1966), .B(G168), .ZN(n959) );
  NAND2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1054 ( .A(KEYINPUT57), .B(n960), .Z(n961) );
  NOR2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n965) );
  XOR2_X1 U1056 ( .A(G16), .B(KEYINPUT56), .Z(n963) );
  XNOR2_X1 U1057 ( .A(KEYINPUT120), .B(n963), .ZN(n964) );
  NOR2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n992) );
  XNOR2_X1 U1059 ( .A(G1966), .B(G21), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(G1961), .B(G5), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n979) );
  XOR2_X1 U1062 ( .A(G4), .B(KEYINPUT124), .Z(n969) );
  XNOR2_X1 U1063 ( .A(G1348), .B(KEYINPUT59), .ZN(n968) );
  XNOR2_X1 U1064 ( .A(n969), .B(n968), .ZN(n976) );
  XNOR2_X1 U1065 ( .A(G19), .B(n970), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(G1956), .B(G20), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(G6), .B(G1981), .ZN(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(n977), .B(KEYINPUT60), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n987) );
  XNOR2_X1 U1073 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n985) );
  XOR2_X1 U1074 ( .A(G1986), .B(G24), .Z(n983) );
  XNOR2_X1 U1075 ( .A(G1971), .B(G22), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(G23), .B(G1976), .ZN(n980) );
  NOR2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1079 ( .A(n985), .B(n984), .Z(n986) );
  NOR2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1081 ( .A(KEYINPUT61), .B(n988), .Z(n989) );
  NOR2_X1 U1082 ( .A1(G16), .A2(n989), .ZN(n990) );
  XNOR2_X1 U1083 ( .A(n990), .B(KEYINPUT126), .ZN(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(n993), .B(KEYINPUT127), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1087 ( .A1(G11), .A2(n996), .ZN(n1026) );
  INV_X1 U1088 ( .A(KEYINPUT55), .ZN(n1022) );
  XNOR2_X1 U1089 ( .A(KEYINPUT52), .B(KEYINPUT116), .ZN(n1020) );
  XNOR2_X1 U1090 ( .A(G160), .B(G2084), .ZN(n998) );
  NAND2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1014) );
  XNOR2_X1 U1094 ( .A(G164), .B(G2078), .ZN(n1003) );
  XNOR2_X1 U1095 ( .A(n1003), .B(KEYINPUT115), .ZN(n1006) );
  XOR2_X1 U1096 ( .A(G2072), .B(n1004), .Z(n1005) );
  NOR2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1098 ( .A(KEYINPUT50), .B(n1007), .ZN(n1012) );
  XOR2_X1 U1099 ( .A(G2090), .B(G162), .Z(n1008) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1101 ( .A(KEYINPUT51), .B(n1010), .Z(n1011) );
  NAND2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(n1020), .B(n1019), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(G29), .ZN(n1024) );
  XNOR2_X1 U1109 ( .A(n1024), .B(KEYINPUT117), .ZN(n1025) );
  NOR2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1111 ( .A(n1027), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

