//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n459), .B1(new_n449), .B2(new_n455), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT68), .Z(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  OAI21_X1  g037(.A(G2104), .B1(KEYINPUT71), .B2(KEYINPUT3), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT71), .A2(KEYINPUT3), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT69), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT70), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n467), .A2(new_n469), .A3(new_n472), .A4(KEYINPUT3), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n465), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n474), .A2(G137), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(KEYINPUT69), .B(G2104), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n481), .A2(G2105), .B1(G101), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n476), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  NAND2_X1  g061(.A1(new_n474), .A2(new_n475), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n474), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n475), .A2(G112), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n489), .B(new_n491), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  XOR2_X1   g069(.A(new_n494), .B(KEYINPUT72), .Z(G162));
  NAND2_X1  g070(.A1(new_n475), .A2(G138), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n479), .A2(KEYINPUT4), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n465), .ZN(new_n498));
  INV_X1    g073(.A(new_n496), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n472), .B1(new_n482), .B2(KEYINPUT3), .ZN(new_n500));
  AND4_X1   g075(.A1(new_n472), .A2(new_n467), .A3(new_n469), .A4(KEYINPUT3), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n498), .B(new_n499), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n497), .B1(new_n502), .B2(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(G126), .A2(G2105), .ZN(new_n504));
  AOI211_X1 g079(.A(new_n465), .B(new_n504), .C1(new_n471), .C2(new_n473), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(G114), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(G2105), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT73), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n504), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n498), .B(new_n510), .C1(new_n500), .C2(new_n501), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n512));
  INV_X1    g087(.A(new_n508), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n503), .B1(new_n509), .B2(new_n514), .ZN(G164));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT74), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT74), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT5), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n523), .B2(KEYINPUT75), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n525), .A2(KEYINPUT5), .A3(G543), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n521), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(G75), .A2(G543), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n520), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n524), .A2(new_n526), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT6), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n531), .B1(new_n517), .B2(new_n519), .ZN(new_n532));
  NOR2_X1   g107(.A1(KEYINPUT6), .A2(G651), .ZN(new_n533));
  OAI211_X1 g108(.A(G88), .B(new_n530), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  OAI211_X1 g109(.A(G50), .B(G543), .C1(new_n532), .C2(new_n533), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n529), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT76), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(G166));
  OAI21_X1  g115(.A(G543), .B1(new_n532), .B2(new_n533), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G51), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT77), .B(G89), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AND2_X1   g122(.A1(G63), .A2(G651), .ZN(new_n548));
  NAND3_X1  g123(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(KEYINPUT7), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(KEYINPUT7), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n530), .A2(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n543), .A2(new_n547), .A3(new_n552), .ZN(G286));
  INV_X1    g128(.A(G286), .ZN(G168));
  NAND2_X1  g129(.A1(new_n542), .A2(G52), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n545), .A2(G90), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n530), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n557));
  INV_X1    g132(.A(new_n520), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n555), .A2(new_n556), .A3(new_n559), .ZN(G301));
  INV_X1    g135(.A(G301), .ZN(G171));
  NAND2_X1  g136(.A1(new_n542), .A2(G43), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n545), .A2(G81), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n530), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n558), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  INV_X1    g147(.A(G53), .ZN(new_n573));
  OR3_X1    g148(.A1(new_n541), .A2(KEYINPUT9), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT9), .B1(new_n541), .B2(new_n573), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n524), .A2(new_n526), .ZN(new_n578));
  INV_X1    g153(.A(G65), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n545), .A2(G91), .B1(new_n580), .B2(G651), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n576), .A2(new_n581), .ZN(G299));
  INV_X1    g157(.A(G166), .ZN(G303));
  OAI21_X1  g158(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n584));
  INV_X1    g159(.A(G87), .ZN(new_n585));
  INV_X1    g160(.A(G49), .ZN(new_n586));
  OAI221_X1 g161(.A(new_n584), .B1(new_n544), .B2(new_n585), .C1(new_n586), .C2(new_n541), .ZN(G288));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n578), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n590), .A2(new_n591), .A3(new_n520), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n591), .B1(new_n590), .B2(new_n520), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G48), .ZN(new_n596));
  INV_X1    g171(.A(G86), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n596), .A2(new_n541), .B1(new_n544), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(G305));
  AOI22_X1  g175(.A1(G47), .A2(new_n542), .B1(new_n545), .B2(G85), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n530), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n558), .B2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT79), .Z(new_n605));
  NAND2_X1  g180(.A1(new_n545), .A2(G92), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XOR2_X1   g183(.A(KEYINPUT80), .B(G66), .Z(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(new_n530), .B1(G79), .B2(G543), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n610), .A2(KEYINPUT81), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n516), .B1(new_n610), .B2(KEYINPUT81), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n611), .A2(new_n612), .B1(G54), .B2(new_n542), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT82), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT83), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT82), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n614), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(KEYINPUT83), .ZN(new_n620));
  AND2_X1   g195(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n605), .B1(new_n621), .B2(G868), .ZN(G284));
  OAI21_X1  g197(.A(new_n605), .B1(new_n621), .B2(G868), .ZN(G321));
  NAND2_X1  g198(.A1(G286), .A2(G868), .ZN(new_n624));
  AND2_X1   g199(.A1(new_n576), .A2(new_n581), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G297));
  OAI21_X1  g201(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n621), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND3_X1  g204(.A1(new_n617), .A2(new_n620), .A3(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G868), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(G868), .B2(new_n567), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n483), .A2(new_n478), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2100), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n488), .A2(G135), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n490), .A2(G123), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT84), .ZN(new_n640));
  OR3_X1    g215(.A1(new_n640), .A2(new_n475), .A3(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n475), .B2(G111), .ZN(new_n642));
  OR2_X1    g217(.A1(G99), .A2(G2105), .ZN(new_n643));
  NAND4_X1  g218(.A1(new_n641), .A2(G2104), .A3(new_n642), .A4(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n638), .A2(new_n639), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT85), .B(G2096), .Z(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n637), .A2(new_n647), .A3(new_n648), .ZN(G156));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT87), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2427), .B(G2430), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G1341), .B(G1348), .Z(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2451), .B(G2454), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(G14), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n663), .B2(new_n660), .ZN(G401));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2100), .ZN(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n669), .B2(KEYINPUT18), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2096), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n680), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(KEYINPUT88), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n682), .A2(new_n683), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT20), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT89), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1981), .B(G1986), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  NAND2_X1  g272(.A1(G162), .A2(G29), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G29), .B2(G35), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(KEYINPUT29), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT29), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n698), .B(new_n701), .C1(G29), .C2(G35), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n700), .A2(G2090), .A3(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT101), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT90), .B(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G20), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT23), .Z(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G299), .B2(G16), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1956), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n700), .A2(KEYINPUT101), .A3(G2090), .A4(new_n702), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n705), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(KEYINPUT102), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n645), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT99), .Z(new_n716));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n717), .A2(G21), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G286), .B2(G16), .ZN(new_n719));
  INV_X1    g294(.A(G1966), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT30), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n722), .A2(G28), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n714), .B1(new_n722), .B2(G28), .ZN(new_n724));
  AND2_X1   g299(.A1(KEYINPUT31), .A2(G11), .ZN(new_n725));
  NOR2_X1   g300(.A1(KEYINPUT31), .A2(G11), .ZN(new_n726));
  OAI22_X1  g301(.A1(new_n723), .A2(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n721), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n717), .A2(G5), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G171), .B2(new_n717), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n730), .A2(G1961), .B1(new_n720), .B2(new_n719), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n716), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT100), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n714), .A2(G32), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n490), .A2(G129), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT98), .ZN(new_n736));
  NAND3_X1  g311(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT26), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n483), .A2(G105), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n738), .B(new_n739), .C1(new_n488), .C2(G141), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n734), .B1(new_n742), .B2(new_n714), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT27), .B(G1996), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n730), .A2(G1961), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n706), .A2(G19), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n567), .B2(new_n706), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n746), .B1(G1341), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G1341), .B2(new_n748), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n751));
  INV_X1    g326(.A(new_n497), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AND3_X1   g328(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n512), .B1(new_n511), .B2(new_n513), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G29), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n714), .A2(G27), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n750), .B1(G2078), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n733), .A2(new_n745), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n714), .A2(G33), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT25), .Z(new_n765));
  AOI22_X1  g340(.A1(new_n478), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n765), .B1(new_n766), .B2(new_n475), .ZN(new_n767));
  INV_X1    g342(.A(G139), .ZN(new_n768));
  OR3_X1    g343(.A1(new_n487), .A2(KEYINPUT94), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(KEYINPUT94), .B1(new_n487), .B2(new_n768), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n767), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n763), .B1(new_n771), .B2(new_n714), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT95), .ZN(new_n773));
  INV_X1    g348(.A(G2072), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT96), .Z(new_n776));
  NAND2_X1  g351(.A1(new_n714), .A2(G26), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT28), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n488), .A2(G140), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n490), .A2(G128), .ZN(new_n780));
  OR2_X1    g355(.A1(G104), .A2(G2105), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n781), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n779), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n778), .B1(new_n783), .B2(G29), .ZN(new_n784));
  INV_X1    g359(.A(G2067), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G2078), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(new_n759), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT24), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(G34), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(G34), .ZN(new_n791));
  AOI21_X1  g366(.A(G29), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n485), .B2(G29), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT97), .ZN(new_n794));
  INV_X1    g369(.A(G2084), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n788), .B(new_n796), .C1(new_n774), .C2(new_n773), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n762), .A2(new_n776), .A3(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT102), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n705), .A2(new_n799), .A3(new_n710), .A4(new_n711), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n700), .A2(new_n702), .ZN(new_n801));
  INV_X1    g376(.A(G2090), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(G1348), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n717), .A2(G4), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n804), .B(new_n805), .C1(new_n621), .C2(new_n717), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n621), .B2(new_n717), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(G1348), .ZN(new_n808));
  AND3_X1   g383(.A1(new_n803), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n713), .A2(new_n798), .A3(new_n800), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n717), .A2(G23), .ZN(new_n811));
  INV_X1    g386(.A(G288), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(new_n717), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT33), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G1976), .ZN(new_n815));
  INV_X1    g390(.A(new_n706), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(G22), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G166), .B2(new_n816), .ZN(new_n818));
  INV_X1    g393(.A(G1971), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n717), .A2(G6), .ZN(new_n821));
  INV_X1    g396(.A(G305), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n822), .B2(new_n717), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT32), .B(G1981), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT91), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n823), .B(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n815), .A2(new_n820), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(KEYINPUT34), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT34), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n815), .A2(new_n826), .A3(new_n829), .A4(new_n820), .ZN(new_n830));
  NOR2_X1   g405(.A1(G25), .A2(G29), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n488), .A2(G131), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n490), .A2(G119), .ZN(new_n833));
  OR2_X1    g408(.A1(G95), .A2(G2105), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n834), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n832), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n831), .B1(new_n836), .B2(G29), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT35), .B(G1991), .Z(new_n838));
  XOR2_X1   g413(.A(new_n837), .B(new_n838), .Z(new_n839));
  MUX2_X1   g414(.A(G24), .B(G290), .S(new_n816), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G1986), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n828), .A2(new_n830), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(KEYINPUT93), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT93), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n828), .A2(new_n845), .A3(new_n830), .A4(new_n842), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT92), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n847), .A2(new_n848), .A3(KEYINPUT36), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT36), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n844), .B(new_n846), .C1(KEYINPUT92), .C2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n810), .B1(new_n849), .B2(new_n851), .ZN(G311));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n851), .ZN(new_n853));
  AND3_X1   g428(.A1(new_n798), .A2(new_n800), .A3(new_n809), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n853), .A2(new_n713), .A3(new_n854), .ZN(G150));
  NAND2_X1  g430(.A1(new_n621), .A2(G559), .ZN(new_n856));
  XOR2_X1   g431(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n857), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n621), .A2(G559), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n542), .A2(G55), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n545), .A2(G93), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n862), .B(new_n863), .C1(new_n558), .C2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n566), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n567), .B(new_n865), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n858), .A2(new_n868), .A3(new_n860), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n871));
  AOI21_X1  g446(.A(G860), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n872), .B1(new_n871), .B2(new_n870), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n865), .A2(G860), .ZN(new_n874));
  XOR2_X1   g449(.A(KEYINPUT104), .B(KEYINPUT37), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n873), .A2(new_n876), .ZN(G145));
  XNOR2_X1  g452(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n645), .B(G160), .ZN(new_n880));
  XOR2_X1   g455(.A(G162), .B(new_n880), .Z(new_n881));
  INV_X1    g456(.A(new_n771), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n741), .A2(new_n783), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n741), .A2(new_n783), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n511), .A2(new_n513), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n503), .A2(new_n885), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n886), .B1(new_n883), .B2(new_n884), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n882), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n883), .A2(new_n884), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n503), .A2(new_n885), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(new_n771), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n488), .A2(G142), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n490), .A2(G130), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n475), .A2(G118), .ZN(new_n897));
  OAI21_X1  g472(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n895), .B(new_n896), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(new_n635), .ZN(new_n900));
  INV_X1    g475(.A(new_n836), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n900), .B(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n889), .A2(new_n894), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n889), .A2(new_n894), .ZN(new_n906));
  INV_X1    g481(.A(new_n902), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n906), .A2(new_n904), .A3(new_n907), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n881), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n908), .A2(new_n881), .A3(new_n903), .ZN(new_n912));
  INV_X1    g487(.A(G37), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n879), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n914), .ZN(new_n916));
  INV_X1    g491(.A(new_n881), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n902), .B1(new_n889), .B2(new_n894), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n918), .B1(new_n904), .B2(new_n903), .ZN(new_n919));
  INV_X1    g494(.A(new_n910), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n916), .A2(new_n921), .A3(new_n878), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n915), .A2(new_n922), .ZN(G395));
  XOR2_X1   g498(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n924));
  NAND2_X1  g499(.A1(new_n630), .A2(new_n868), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n614), .A2(G299), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n625), .A2(new_n608), .A3(new_n613), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n617), .A2(new_n620), .A3(new_n628), .A4(new_n866), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n925), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n928), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT41), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT41), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n928), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(new_n925), .B2(new_n929), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n924), .B1(new_n931), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n924), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n925), .A2(new_n929), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n939), .B(new_n930), .C1(new_n940), .C2(new_n936), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n822), .A2(G166), .ZN(new_n942));
  NAND2_X1  g517(.A1(G303), .A2(G305), .ZN(new_n943));
  XNOR2_X1  g518(.A(G290), .B(new_n812), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n942), .B(new_n943), .C1(new_n944), .C2(KEYINPUT107), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(KEYINPUT107), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n945), .B(new_n946), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n938), .A2(new_n941), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n947), .B1(new_n938), .B2(new_n941), .ZN(new_n949));
  OAI21_X1  g524(.A(G868), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G868), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n865), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(G295));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n952), .ZN(G331));
  NAND2_X1  g529(.A1(new_n866), .A2(G171), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n866), .A2(G171), .ZN(new_n957));
  OAI21_X1  g532(.A(G286), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n957), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(G168), .A3(new_n955), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n932), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n958), .A2(new_n960), .A3(new_n935), .A4(new_n933), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n947), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n962), .A2(new_n947), .A3(new_n963), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(new_n913), .A3(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n972));
  AOI21_X1  g547(.A(G37), .B1(new_n964), .B2(new_n965), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n973), .A2(new_n969), .A3(new_n967), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(KEYINPUT110), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n973), .A2(new_n977), .A3(new_n969), .A4(new_n967), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n975), .B1(KEYINPUT44), .B2(new_n980), .ZN(G397));
  INV_X1    g556(.A(G1384), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(new_n503), .B2(new_n885), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT45), .B1(new_n983), .B2(KEYINPUT111), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(KEYINPUT111), .B2(new_n983), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n476), .A2(G40), .A3(new_n484), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1996), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n741), .B(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n783), .B(new_n785), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n836), .B(new_n838), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n987), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(G290), .A2(G1986), .ZN(new_n994));
  AND2_X1   g569(.A1(G290), .A2(G1986), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n987), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n997), .B(KEYINPUT112), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n999));
  INV_X1    g574(.A(G8), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n999), .B1(G166), .B2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n538), .A2(KEYINPUT55), .A3(G8), .A4(new_n539), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT45), .B1(new_n756), .B2(new_n982), .ZN(new_n1005));
  INV_X1    g580(.A(new_n986), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT45), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1007), .A2(G1384), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1006), .B1(new_n891), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n819), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n756), .A2(new_n1012), .A3(new_n982), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n986), .B1(new_n983), .B2(KEYINPUT50), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1013), .A2(new_n1014), .A3(new_n802), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1004), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1016), .A2(new_n1000), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n1011), .A2(new_n1015), .A3(new_n1004), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1003), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n986), .B1(new_n886), .B2(new_n1008), .ZN(new_n1021));
  NOR2_X1   g596(.A1(G164), .A2(G1384), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1021), .B(new_n787), .C1(new_n1022), .C2(KEYINPUT45), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(G164), .B2(new_n1009), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n756), .A2(KEYINPUT116), .A3(new_n1008), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n986), .B1(new_n983), .B2(new_n1007), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1024), .A2(G2078), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1012), .B(new_n982), .C1(new_n503), .C2(new_n885), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1032), .A2(new_n1006), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1033), .B1(new_n1022), .B2(new_n1012), .ZN(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT124), .B(G1961), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1025), .A2(new_n1031), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(G171), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1033), .B(new_n802), .C1(new_n1022), .C2(new_n1012), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1000), .B1(new_n1039), .B2(new_n1011), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1001), .A2(new_n1041), .A3(new_n1002), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1041), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n886), .A2(new_n982), .A3(new_n1006), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n812), .A2(G1976), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1046), .A2(G8), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT52), .ZN(new_n1049));
  INV_X1    g624(.A(G1981), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n599), .B(new_n1050), .C1(new_n593), .C2(new_n594), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n590), .A2(new_n520), .ZN(new_n1052));
  OAI21_X1  g627(.A(G1981), .B1(new_n1052), .B2(new_n598), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT49), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1051), .A2(KEYINPUT49), .A3(new_n1053), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1056), .A2(G8), .A3(new_n1046), .A4(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G1976), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT52), .B1(G288), .B2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1046), .A2(G8), .A3(new_n1047), .A4(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1049), .A2(new_n1058), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1045), .A2(new_n1063), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1020), .A2(new_n1038), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT126), .ZN(new_n1066));
  NAND2_X1  g641(.A1(G286), .A2(G8), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n720), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1012), .B1(new_n756), .B2(new_n982), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1032), .A2(new_n1006), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n795), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1071), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1069), .B1(new_n1076), .B2(G8), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(G8), .ZN(new_n1078));
  XOR2_X1   g653(.A(new_n1067), .B(KEYINPUT123), .Z(new_n1079));
  AOI21_X1  g654(.A(new_n1068), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1076), .A2(G8), .A3(G286), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1077), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1065), .B(new_n1066), .C1(new_n1082), .C2(KEYINPUT62), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n720), .A2(new_n1070), .B1(new_n1074), .B2(new_n795), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1079), .B1(new_n1084), .B2(new_n1000), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1085), .A2(new_n1081), .A3(KEYINPUT51), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1077), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT62), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1062), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1023), .A2(new_n1024), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1090));
  AOI21_X1  g665(.A(G301), .B1(new_n1090), .B2(new_n1031), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1018), .A2(new_n1016), .A3(new_n1000), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1089), .B(new_n1091), .C1(new_n1092), .C2(new_n1003), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT126), .B1(new_n1088), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1082), .A2(KEYINPUT62), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1083), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1046), .A2(G8), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1097), .B(KEYINPUT114), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1058), .A2(new_n1059), .A3(new_n812), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1051), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1045), .B2(new_n1062), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1084), .A2(new_n1000), .A3(G286), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1089), .B(new_n1103), .C1(new_n1092), .C2(new_n1003), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT63), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1040), .A2(new_n1003), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1089), .A2(new_n1103), .A3(new_n1107), .A4(KEYINPUT63), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1102), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n886), .A2(KEYINPUT119), .A3(new_n982), .A4(new_n1006), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n983), .B2(new_n986), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1034), .A2(new_n804), .B1(new_n1113), .B2(new_n785), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1114), .A2(new_n619), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1116), .A2(KEYINPUT57), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(KEYINPUT57), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n625), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(G299), .A2(new_n1116), .A3(KEYINPUT57), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1122));
  INV_X1    g697(.A(G1956), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT56), .B(G2072), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1021), .B(new_n1125), .C1(new_n1022), .C2(KEYINPUT45), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1115), .A2(KEYINPUT120), .B1(new_n1121), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT120), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(new_n1114), .B2(new_n619), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1125), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1005), .A2(new_n1010), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(G1956), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1135));
  AOI21_X1  g710(.A(KEYINPUT118), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1124), .A2(new_n1135), .A3(new_n1126), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT118), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1128), .A2(new_n1130), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1121), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1143), .A2(new_n1138), .A3(KEYINPUT61), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1143), .A2(new_n1138), .A3(KEYINPUT121), .A4(KEYINPUT61), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1144), .A2(new_n1145), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g725(.A(KEYINPUT58), .B(G1341), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1113), .A2(new_n1151), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1005), .A2(G1996), .A3(new_n1010), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n567), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT59), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  OAI211_X1 g731(.A(KEYINPUT59), .B(new_n567), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1114), .A2(KEYINPUT60), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT122), .B1(new_n1114), .B2(KEYINPUT60), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1159), .B1(new_n1160), .B2(new_n619), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1113), .A2(new_n785), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1162), .B(KEYINPUT60), .C1(G1348), .C2(new_n1074), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT122), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1114), .A2(KEYINPUT122), .A3(KEYINPUT60), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1165), .A2(new_n615), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1158), .B1(new_n1161), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1142), .B1(new_n1150), .B2(new_n1168), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1010), .A2(new_n1024), .A3(G2078), .ZN(new_n1170));
  AOI21_X1  g745(.A(KEYINPUT125), .B1(new_n1170), .B2(new_n985), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1170), .A2(new_n985), .A3(KEYINPUT125), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1090), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(G171), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1090), .A2(G301), .A3(new_n1031), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1174), .A2(KEYINPUT54), .A3(new_n1175), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1090), .B(G301), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n1038), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT54), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1020), .A2(new_n1064), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1082), .A2(new_n1176), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1109), .B1(new_n1169), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n998), .B1(new_n1096), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n836), .A2(new_n838), .ZN(new_n1185));
  OAI22_X1  g760(.A1(new_n991), .A2(new_n1185), .B1(G2067), .B2(new_n783), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1186), .A2(new_n987), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n987), .A2(new_n988), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n1188), .B(KEYINPUT46), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n742), .A2(new_n990), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n987), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT47), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1192), .B(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n987), .A2(new_n994), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1195), .B(KEYINPUT48), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n993), .B(KEYINPUT127), .ZN(new_n1197));
  AOI211_X1 g772(.A(new_n1187), .B(new_n1194), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1184), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g774(.A1(new_n971), .A2(new_n974), .ZN(new_n1201));
  NOR4_X1   g775(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1202));
  OAI211_X1 g776(.A(new_n1201), .B(new_n1202), .C1(new_n911), .C2(new_n914), .ZN(G225));
  INV_X1    g777(.A(G225), .ZN(G308));
endmodule


