

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595;

  NOR2_X1 U326 ( .A1(n554), .A2(n536), .ZN(n539) );
  XNOR2_X1 U327 ( .A(n422), .B(KEYINPUT64), .ZN(n423) );
  INV_X1 U328 ( .A(KEYINPUT48), .ZN(n422) );
  XNOR2_X1 U329 ( .A(n491), .B(n490), .ZN(n492) );
  INV_X1 U330 ( .A(KEYINPUT107), .ZN(n490) );
  XNOR2_X1 U331 ( .A(n369), .B(n294), .ZN(n332) );
  XOR2_X1 U332 ( .A(KEYINPUT41), .B(n583), .Z(n571) );
  AND2_X1 U333 ( .A1(G226GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U334 ( .A(G176GAT), .B(G92GAT), .ZN(n331) );
  XNOR2_X1 U335 ( .A(KEYINPUT27), .B(KEYINPUT102), .ZN(n477) );
  XNOR2_X1 U336 ( .A(n331), .B(G64GAT), .ZN(n391) );
  XNOR2_X1 U337 ( .A(n529), .B(n477), .ZN(n484) );
  XNOR2_X1 U338 ( .A(n424), .B(n423), .ZN(n552) );
  XNOR2_X1 U339 ( .A(n493), .B(n492), .ZN(n525) );
  XNOR2_X1 U340 ( .A(n408), .B(n407), .ZN(n583) );
  XNOR2_X1 U341 ( .A(n470), .B(G190GAT), .ZN(n471) );
  XNOR2_X1 U342 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n496) );
  XNOR2_X1 U343 ( .A(n472), .B(n471), .ZN(G1351GAT) );
  XNOR2_X1 U344 ( .A(n497), .B(n496), .ZN(G1330GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n296) );
  XNOR2_X1 U346 ( .A(G106GAT), .B(KEYINPUT78), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n308) );
  XOR2_X1 U348 ( .A(G99GAT), .B(G85GAT), .Z(n398) );
  XOR2_X1 U349 ( .A(KEYINPUT10), .B(n398), .Z(n298) );
  XOR2_X1 U350 ( .A(G29GAT), .B(G134GAT), .Z(n434) );
  XNOR2_X1 U351 ( .A(G218GAT), .B(n434), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U353 ( .A(n299), .B(G92GAT), .Z(n306) );
  XNOR2_X1 U354 ( .A(G36GAT), .B(G190GAT), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n300), .B(KEYINPUT79), .ZN(n337) );
  INV_X1 U356 ( .A(KEYINPUT77), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n337), .B(n301), .ZN(n303) );
  NAND2_X1 U358 ( .A1(G232GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U360 ( .A(G162GAT), .B(n304), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U363 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n310) );
  XNOR2_X1 U364 ( .A(G50GAT), .B(G43GAT), .ZN(n309) );
  XNOR2_X1 U365 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U366 ( .A(KEYINPUT68), .B(n311), .ZN(n380) );
  XNOR2_X1 U367 ( .A(n312), .B(n380), .ZN(n469) );
  XOR2_X1 U368 ( .A(G113GAT), .B(KEYINPUT0), .Z(n446) );
  XOR2_X1 U369 ( .A(G190GAT), .B(G99GAT), .Z(n314) );
  XNOR2_X1 U370 ( .A(G43GAT), .B(G134GAT), .ZN(n313) );
  XNOR2_X1 U371 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U372 ( .A(n446), .B(n315), .Z(n317) );
  NAND2_X1 U373 ( .A1(G227GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U375 ( .A(n318), .B(G71GAT), .Z(n322) );
  XOR2_X1 U376 ( .A(G183GAT), .B(KEYINPUT17), .Z(n320) );
  XNOR2_X1 U377 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n338) );
  XNOR2_X1 U379 ( .A(G15GAT), .B(n338), .ZN(n321) );
  XNOR2_X1 U380 ( .A(n322), .B(n321), .ZN(n330) );
  XOR2_X1 U381 ( .A(G127GAT), .B(KEYINPUT88), .Z(n324) );
  XNOR2_X1 U382 ( .A(G169GAT), .B(G120GAT), .ZN(n323) );
  XNOR2_X1 U383 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U384 ( .A(G176GAT), .B(KEYINPUT65), .Z(n326) );
  XNOR2_X1 U385 ( .A(KEYINPUT87), .B(KEYINPUT20), .ZN(n325) );
  XNOR2_X1 U386 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U387 ( .A(n328), .B(n327), .Z(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n541) );
  XNOR2_X1 U389 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n426) );
  XOR2_X1 U390 ( .A(G169GAT), .B(G8GAT), .Z(n369) );
  XNOR2_X1 U391 ( .A(n332), .B(n391), .ZN(n336) );
  XOR2_X1 U392 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n334) );
  XNOR2_X1 U393 ( .A(G204GAT), .B(KEYINPUT99), .ZN(n333) );
  XNOR2_X1 U394 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U395 ( .A(n336), .B(n335), .Z(n340) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U397 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U398 ( .A(KEYINPUT89), .B(G218GAT), .Z(n342) );
  XNOR2_X1 U399 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n341) );
  XNOR2_X1 U400 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U401 ( .A(G197GAT), .B(n343), .ZN(n462) );
  XNOR2_X1 U402 ( .A(n344), .B(n462), .ZN(n529) );
  XOR2_X1 U403 ( .A(KEYINPUT115), .B(KEYINPUT47), .Z(n415) );
  XOR2_X1 U404 ( .A(G71GAT), .B(KEYINPUT13), .Z(n397) );
  XOR2_X1 U405 ( .A(G1GAT), .B(G127GAT), .Z(n430) );
  XOR2_X1 U406 ( .A(n397), .B(n430), .Z(n346) );
  XNOR2_X1 U407 ( .A(G211GAT), .B(G78GAT), .ZN(n345) );
  XNOR2_X1 U408 ( .A(n346), .B(n345), .ZN(n351) );
  XNOR2_X1 U409 ( .A(G15GAT), .B(G22GAT), .ZN(n347) );
  XNOR2_X1 U410 ( .A(n347), .B(KEYINPUT69), .ZN(n372) );
  XOR2_X1 U411 ( .A(n372), .B(KEYINPUT14), .Z(n349) );
  NAND2_X1 U412 ( .A1(G231GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U413 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U414 ( .A(n351), .B(n350), .Z(n353) );
  XNOR2_X1 U415 ( .A(G183GAT), .B(G155GAT), .ZN(n352) );
  XNOR2_X1 U416 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U417 ( .A(KEYINPUT12), .B(G64GAT), .Z(n355) );
  XNOR2_X1 U418 ( .A(G8GAT), .B(G57GAT), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U420 ( .A(n357), .B(n356), .Z(n365) );
  XOR2_X1 U421 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n359) );
  XNOR2_X1 U422 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n358) );
  XNOR2_X1 U423 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U424 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n361) );
  XNOR2_X1 U425 ( .A(KEYINPUT86), .B(KEYINPUT85), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U427 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n563) );
  INV_X1 U429 ( .A(n563), .ZN(n588) );
  XNOR2_X1 U430 ( .A(KEYINPUT46), .B(KEYINPUT114), .ZN(n410) );
  XOR2_X1 U431 ( .A(G1GAT), .B(G197GAT), .Z(n367) );
  XNOR2_X1 U432 ( .A(G113GAT), .B(G141GAT), .ZN(n366) );
  XNOR2_X1 U433 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U434 ( .A(n368), .B(G36GAT), .Z(n371) );
  XNOR2_X1 U435 ( .A(n369), .B(G29GAT), .ZN(n370) );
  XNOR2_X1 U436 ( .A(n371), .B(n370), .ZN(n376) );
  XOR2_X1 U437 ( .A(KEYINPUT29), .B(n372), .Z(n374) );
  NAND2_X1 U438 ( .A1(G229GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U439 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U440 ( .A(n376), .B(n375), .Z(n382) );
  XOR2_X1 U441 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n378) );
  XNOR2_X1 U442 ( .A(KEYINPUT30), .B(KEYINPUT70), .ZN(n377) );
  XNOR2_X1 U443 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U444 ( .A(n380), .B(n379), .Z(n381) );
  XNOR2_X1 U445 ( .A(n382), .B(n381), .ZN(n579) );
  INV_X1 U446 ( .A(n391), .ZN(n390) );
  INV_X1 U447 ( .A(KEYINPUT32), .ZN(n383) );
  NAND2_X1 U448 ( .A1(KEYINPUT31), .A2(n383), .ZN(n386) );
  INV_X1 U449 ( .A(KEYINPUT31), .ZN(n384) );
  NAND2_X1 U450 ( .A1(n384), .A2(KEYINPUT32), .ZN(n385) );
  NAND2_X1 U451 ( .A1(n386), .A2(n385), .ZN(n388) );
  XNOR2_X1 U452 ( .A(KEYINPUT74), .B(KEYINPUT33), .ZN(n387) );
  XNOR2_X1 U453 ( .A(n388), .B(n387), .ZN(n392) );
  INV_X1 U454 ( .A(n392), .ZN(n389) );
  NAND2_X1 U455 ( .A1(n390), .A2(n389), .ZN(n394) );
  NAND2_X1 U456 ( .A1(n392), .A2(n391), .ZN(n393) );
  NAND2_X1 U457 ( .A1(n394), .A2(n393), .ZN(n396) );
  XOR2_X1 U458 ( .A(KEYINPUT71), .B(KEYINPUT75), .Z(n395) );
  XNOR2_X1 U459 ( .A(n396), .B(n395), .ZN(n402) );
  XOR2_X1 U460 ( .A(n398), .B(n397), .Z(n400) );
  NAND2_X1 U461 ( .A1(G230GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U462 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U463 ( .A(n402), .B(n401), .Z(n408) );
  XNOR2_X1 U464 ( .A(G148GAT), .B(KEYINPUT72), .ZN(n403) );
  XNOR2_X1 U465 ( .A(n403), .B(KEYINPUT73), .ZN(n404) );
  XNOR2_X1 U466 ( .A(n404), .B(G204GAT), .ZN(n406) );
  XOR2_X1 U467 ( .A(G78GAT), .B(G106GAT), .Z(n405) );
  XNOR2_X1 U468 ( .A(n406), .B(n405), .ZN(n456) );
  XOR2_X1 U469 ( .A(G120GAT), .B(G57GAT), .Z(n433) );
  XNOR2_X1 U470 ( .A(n456), .B(n433), .ZN(n407) );
  NOR2_X1 U471 ( .A1(n579), .A2(n571), .ZN(n409) );
  XNOR2_X1 U472 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U473 ( .A(n411), .B(KEYINPUT113), .ZN(n412) );
  AND2_X1 U474 ( .A1(n588), .A2(n412), .ZN(n413) );
  NAND2_X1 U475 ( .A1(n413), .A2(n469), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n415), .B(n414), .ZN(n421) );
  INV_X1 U477 ( .A(n469), .ZN(n498) );
  XNOR2_X1 U478 ( .A(n498), .B(KEYINPUT36), .ZN(n591) );
  NAND2_X1 U479 ( .A1(n591), .A2(n563), .ZN(n416) );
  XNOR2_X1 U480 ( .A(n416), .B(KEYINPUT116), .ZN(n417) );
  XNOR2_X1 U481 ( .A(KEYINPUT45), .B(n417), .ZN(n419) );
  NAND2_X1 U482 ( .A1(n583), .A2(n579), .ZN(n418) );
  NOR2_X1 U483 ( .A1(n419), .A2(n418), .ZN(n420) );
  NOR2_X1 U484 ( .A1(n421), .A2(n420), .ZN(n424) );
  NAND2_X1 U485 ( .A1(n529), .A2(n552), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n426), .B(n425), .ZN(n575) );
  XOR2_X1 U487 ( .A(KEYINPUT6), .B(KEYINPUT95), .Z(n428) );
  XNOR2_X1 U488 ( .A(KEYINPUT94), .B(KEYINPUT4), .ZN(n427) );
  XNOR2_X1 U489 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U490 ( .A(n429), .B(G85GAT), .Z(n432) );
  XNOR2_X1 U491 ( .A(G148GAT), .B(n430), .ZN(n431) );
  XNOR2_X1 U492 ( .A(n432), .B(n431), .ZN(n450) );
  XOR2_X1 U493 ( .A(n434), .B(n433), .Z(n436) );
  NAND2_X1 U494 ( .A1(G225GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U496 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n438) );
  XNOR2_X1 U497 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n437) );
  XNOR2_X1 U498 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U499 ( .A(n440), .B(n439), .Z(n448) );
  XOR2_X1 U500 ( .A(KEYINPUT91), .B(KEYINPUT2), .Z(n442) );
  XNOR2_X1 U501 ( .A(G162GAT), .B(KEYINPUT90), .ZN(n441) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U503 ( .A(n443), .B(KEYINPUT3), .Z(n445) );
  XNOR2_X1 U504 ( .A(G141GAT), .B(G155GAT), .ZN(n444) );
  XNOR2_X1 U505 ( .A(n445), .B(n444), .ZN(n461) );
  XNOR2_X1 U506 ( .A(n446), .B(n461), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n450), .B(n449), .ZN(n481) );
  XNOR2_X1 U509 ( .A(KEYINPUT98), .B(n481), .ZN(n527) );
  INV_X1 U510 ( .A(n527), .ZN(n576) );
  XOR2_X1 U511 ( .A(KEYINPUT23), .B(KEYINPUT93), .Z(n452) );
  XNOR2_X1 U512 ( .A(KEYINPUT92), .B(KEYINPUT24), .ZN(n451) );
  XNOR2_X1 U513 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U514 ( .A(KEYINPUT22), .B(n453), .Z(n455) );
  NAND2_X1 U515 ( .A1(G228GAT), .A2(G233GAT), .ZN(n454) );
  XNOR2_X1 U516 ( .A(n455), .B(n454), .ZN(n457) );
  XOR2_X1 U517 ( .A(n457), .B(n456), .Z(n459) );
  XNOR2_X1 U518 ( .A(G50GAT), .B(G22GAT), .ZN(n458) );
  XNOR2_X1 U519 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n461), .B(n460), .ZN(n463) );
  XNOR2_X1 U521 ( .A(n463), .B(n462), .ZN(n486) );
  AND2_X1 U522 ( .A1(n576), .A2(n486), .ZN(n464) );
  NAND2_X1 U523 ( .A1(n575), .A2(n464), .ZN(n466) );
  XOR2_X1 U524 ( .A(KEYINPUT122), .B(KEYINPUT55), .Z(n465) );
  XNOR2_X1 U525 ( .A(n466), .B(n465), .ZN(n467) );
  NOR2_X1 U526 ( .A1(n541), .A2(n467), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n468), .B(KEYINPUT123), .ZN(n567) );
  NOR2_X1 U528 ( .A1(n469), .A2(n567), .ZN(n472) );
  INV_X1 U529 ( .A(KEYINPUT58), .ZN(n470) );
  INV_X1 U530 ( .A(n579), .ZN(n555) );
  NAND2_X1 U531 ( .A1(n555), .A2(n583), .ZN(n473) );
  XNOR2_X1 U532 ( .A(KEYINPUT76), .B(n473), .ZN(n502) );
  INV_X1 U533 ( .A(n541), .ZN(n532) );
  NAND2_X1 U534 ( .A1(n532), .A2(n529), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n474), .B(KEYINPUT104), .ZN(n475) );
  NAND2_X1 U536 ( .A1(n475), .A2(n486), .ZN(n476) );
  XNOR2_X1 U537 ( .A(n476), .B(KEYINPUT25), .ZN(n480) );
  NOR2_X1 U538 ( .A1(n532), .A2(n486), .ZN(n478) );
  XNOR2_X1 U539 ( .A(KEYINPUT26), .B(n478), .ZN(n577) );
  AND2_X1 U540 ( .A1(n484), .A2(n577), .ZN(n479) );
  NOR2_X1 U541 ( .A1(n480), .A2(n479), .ZN(n482) );
  NOR2_X1 U542 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n483), .B(KEYINPUT105), .ZN(n488) );
  NAND2_X1 U544 ( .A1(n484), .A2(n527), .ZN(n485) );
  XOR2_X1 U545 ( .A(KEYINPUT103), .B(n485), .Z(n554) );
  XOR2_X1 U546 ( .A(KEYINPUT28), .B(n486), .Z(n536) );
  NAND2_X1 U547 ( .A1(n539), .A2(n541), .ZN(n487) );
  NAND2_X1 U548 ( .A1(n488), .A2(n487), .ZN(n500) );
  NAND2_X1 U549 ( .A1(n591), .A2(n500), .ZN(n489) );
  NOR2_X1 U550 ( .A1(n563), .A2(n489), .ZN(n493) );
  XNOR2_X1 U551 ( .A(KEYINPUT108), .B(KEYINPUT37), .ZN(n491) );
  OR2_X1 U552 ( .A1(n502), .A2(n525), .ZN(n494) );
  XNOR2_X1 U553 ( .A(n494), .B(KEYINPUT38), .ZN(n495) );
  XNOR2_X1 U554 ( .A(KEYINPUT109), .B(n495), .ZN(n514) );
  NAND2_X1 U555 ( .A1(n514), .A2(n532), .ZN(n497) );
  NOR2_X1 U556 ( .A1(n498), .A2(n588), .ZN(n499) );
  XNOR2_X1 U557 ( .A(n499), .B(KEYINPUT16), .ZN(n501) );
  NAND2_X1 U558 ( .A1(n501), .A2(n500), .ZN(n516) );
  NOR2_X1 U559 ( .A1(n502), .A2(n516), .ZN(n509) );
  NAND2_X1 U560 ( .A1(n509), .A2(n527), .ZN(n503) );
  XNOR2_X1 U561 ( .A(n503), .B(KEYINPUT34), .ZN(n504) );
  XNOR2_X1 U562 ( .A(G1GAT), .B(n504), .ZN(G1324GAT) );
  NAND2_X1 U563 ( .A1(n509), .A2(n529), .ZN(n505) );
  XNOR2_X1 U564 ( .A(n505), .B(KEYINPUT106), .ZN(n506) );
  XNOR2_X1 U565 ( .A(G8GAT), .B(n506), .ZN(G1325GAT) );
  XOR2_X1 U566 ( .A(G15GAT), .B(KEYINPUT35), .Z(n508) );
  NAND2_X1 U567 ( .A1(n509), .A2(n532), .ZN(n507) );
  XNOR2_X1 U568 ( .A(n508), .B(n507), .ZN(G1326GAT) );
  NAND2_X1 U569 ( .A1(n536), .A2(n509), .ZN(n510) );
  XNOR2_X1 U570 ( .A(n510), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U571 ( .A1(n527), .A2(n514), .ZN(n512) );
  XOR2_X1 U572 ( .A(G29GAT), .B(KEYINPUT39), .Z(n511) );
  XNOR2_X1 U573 ( .A(n512), .B(n511), .ZN(G1328GAT) );
  NAND2_X1 U574 ( .A1(n514), .A2(n529), .ZN(n513) );
  XNOR2_X1 U575 ( .A(n513), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U576 ( .A1(n514), .A2(n536), .ZN(n515) );
  XNOR2_X1 U577 ( .A(n515), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U578 ( .A(n571), .ZN(n558) );
  NAND2_X1 U579 ( .A1(n558), .A2(n579), .ZN(n526) );
  NOR2_X1 U580 ( .A1(n526), .A2(n516), .ZN(n521) );
  NAND2_X1 U581 ( .A1(n527), .A2(n521), .ZN(n517) );
  XNOR2_X1 U582 ( .A(KEYINPUT42), .B(n517), .ZN(n518) );
  XNOR2_X1 U583 ( .A(G57GAT), .B(n518), .ZN(G1332GAT) );
  NAND2_X1 U584 ( .A1(n521), .A2(n529), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U586 ( .A1(n521), .A2(n532), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n520), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT43), .B(KEYINPUT110), .Z(n523) );
  NAND2_X1 U589 ( .A1(n521), .A2(n536), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U591 ( .A(G78GAT), .B(n524), .ZN(G1335GAT) );
  NOR2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n527), .A2(n535), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G85GAT), .B(n528), .ZN(G1336GAT) );
  XOR2_X1 U595 ( .A(G92GAT), .B(KEYINPUT111), .Z(n531) );
  NAND2_X1 U596 ( .A1(n535), .A2(n529), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(G1337GAT) );
  NAND2_X1 U598 ( .A1(n535), .A2(n532), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n533), .B(KEYINPUT112), .ZN(n534) );
  XNOR2_X1 U600 ( .A(G99GAT), .B(n534), .ZN(G1338GAT) );
  NAND2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n537), .B(KEYINPUT44), .ZN(n538) );
  XNOR2_X1 U603 ( .A(G106GAT), .B(n538), .ZN(G1339GAT) );
  NAND2_X1 U604 ( .A1(n539), .A2(n552), .ZN(n540) );
  NOR2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n555), .A2(n549), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n542), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n544) );
  NAND2_X1 U609 ( .A1(n549), .A2(n558), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U611 ( .A(G120GAT), .B(n545), .Z(G1341GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n547) );
  NAND2_X1 U613 ( .A1(n549), .A2(n563), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U615 ( .A(G127GAT), .B(n548), .Z(G1342GAT) );
  XOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U617 ( .A1(n549), .A2(n498), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(G1343GAT) );
  XOR2_X1 U619 ( .A(G141GAT), .B(KEYINPUT119), .Z(n557) );
  NAND2_X1 U620 ( .A1(n552), .A2(n577), .ZN(n553) );
  NOR2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n565) );
  NAND2_X1 U622 ( .A1(n565), .A2(n555), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1344GAT) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n562) );
  XOR2_X1 U625 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n560) );
  NAND2_X1 U626 ( .A1(n565), .A2(n558), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1345GAT) );
  NAND2_X1 U629 ( .A1(n565), .A2(n563), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n498), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U633 ( .A1(n579), .A2(n567), .ZN(n568) );
  XOR2_X1 U634 ( .A(G169GAT), .B(n568), .Z(G1348GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT56), .B(KEYINPUT124), .Z(n570) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n573) );
  NOR2_X1 U638 ( .A1(n571), .A2(n567), .ZN(n572) );
  XOR2_X1 U639 ( .A(n573), .B(n572), .Z(G1349GAT) );
  NOR2_X1 U640 ( .A1(n588), .A2(n567), .ZN(n574) );
  XOR2_X1 U641 ( .A(G183GAT), .B(n574), .Z(G1350GAT) );
  AND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n590) );
  NOR2_X1 U644 ( .A1(n579), .A2(n590), .ZN(n581) );
  XNOR2_X1 U645 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(G197GAT), .B(n582), .ZN(G1352GAT) );
  NOR2_X1 U648 ( .A1(n590), .A2(n583), .ZN(n587) );
  XOR2_X1 U649 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n585) );
  XNOR2_X1 U650 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1353GAT) );
  NOR2_X1 U653 ( .A1(n588), .A2(n590), .ZN(n589) );
  XOR2_X1 U654 ( .A(G211GAT), .B(n589), .Z(G1354GAT) );
  XOR2_X1 U655 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n594) );
  INV_X1 U656 ( .A(n590), .ZN(n592) );
  NAND2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U658 ( .A(n594), .B(n593), .ZN(n595) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(n595), .ZN(G1355GAT) );
endmodule

