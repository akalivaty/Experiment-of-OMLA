//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967;
  INV_X1    g000(.A(KEYINPUT80), .ZN(new_n202));
  XOR2_X1   g001(.A(G1gat), .B(G29gat), .Z(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT76), .ZN(new_n209));
  INV_X1    g008(.A(G113gat), .ZN(new_n210));
  INV_X1    g009(.A(G120gat), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT1), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G127gat), .B(G134gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G113gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n212), .B(new_n213), .C1(new_n214), .C2(new_n211), .ZN(new_n215));
  INV_X1    g014(.A(G134gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G127gat), .ZN(new_n217));
  INV_X1    g016(.A(G127gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G134gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G113gat), .B2(G120gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n210), .A2(new_n211), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n220), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n215), .A2(new_n224), .ZN(new_n225));
  AND2_X1   g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G141gat), .B(G148gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT2), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n230), .B1(G155gat), .B2(G162gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n228), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G141gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G148gat), .ZN(new_n234));
  INV_X1    g033(.A(G148gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G141gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G155gat), .B(G162gat), .ZN(new_n238));
  INV_X1    g037(.A(G155gat), .ZN(new_n239));
  INV_X1    g038(.A(G162gat), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT2), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n237), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n232), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n243), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n215), .A2(new_n232), .A3(new_n224), .A4(new_n242), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G225gat), .A2(G233gat), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n209), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  AOI211_X1 g048(.A(KEYINPUT76), .B(new_n247), .C1(new_n244), .C2(new_n245), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT5), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n243), .A2(KEYINPUT3), .B1(new_n224), .B2(new_n215), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n232), .A2(new_n242), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n248), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT75), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n232), .A2(new_n242), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n220), .A2(new_n222), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n210), .A2(KEYINPUT65), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT65), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G113gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G120gat), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n212), .B1(new_n210), .B2(new_n211), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n258), .A2(new_n263), .B1(new_n264), .B2(new_n220), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n257), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT74), .B(KEYINPUT4), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n245), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n255), .A2(new_n256), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n256), .B1(new_n255), .B2(new_n270), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n251), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n255), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n257), .A2(new_n265), .A3(new_n268), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n245), .A2(new_n266), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR3_X1   g076(.A1(new_n274), .A2(new_n277), .A3(KEYINPUT5), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n208), .B1(new_n273), .B2(new_n278), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n249), .A2(new_n250), .ZN(new_n280));
  INV_X1    g079(.A(new_n272), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n255), .A2(new_n256), .A3(new_n270), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT5), .A4(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n278), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n207), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n279), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G226gat), .A2(G233gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT64), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT25), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT24), .ZN(new_n293));
  INV_X1    g092(.A(G183gat), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n293), .B1(new_n294), .B2(G190gat), .ZN(new_n295));
  INV_X1    g094(.A(G190gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G183gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n295), .A2(new_n297), .B1(new_n293), .B2(new_n298), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n289), .A2(new_n290), .B1(G169gat), .B2(G176gat), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NOR3_X1   g101(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n292), .B1(new_n299), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(KEYINPUT64), .B2(KEYINPUT25), .ZN(new_n307));
  NOR2_X1   g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT23), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n307), .B1(new_n301), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n298), .A2(new_n293), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT24), .B1(new_n296), .B2(G183gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n294), .A2(G190gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n311), .A2(new_n291), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n294), .A2(KEYINPUT27), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT27), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G183gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n319), .A3(new_n296), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT27), .B(G183gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n323), .A2(KEYINPUT28), .A3(new_n296), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n306), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n326), .A2(new_n308), .A3(KEYINPUT26), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n308), .A2(KEYINPUT26), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n298), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n305), .A2(new_n316), .B1(new_n325), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n288), .B1(new_n331), .B2(KEYINPUT29), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n325), .A2(new_n330), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n299), .A2(new_n304), .A3(new_n292), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n291), .B1(new_n311), .B2(new_n315), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n288), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT72), .B1(new_n332), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT72), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n340), .B1(new_n342), .B2(new_n288), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT71), .ZN(new_n344));
  XNOR2_X1  g143(.A(G211gat), .B(G218gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(G197gat), .B(G204gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT22), .ZN(new_n347));
  INV_X1    g146(.A(G211gat), .ZN(new_n348));
  INV_X1    g147(.A(G218gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n345), .A2(new_n346), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n345), .B1(new_n350), .B2(new_n346), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n344), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n346), .A2(new_n350), .ZN(new_n355));
  INV_X1    g154(.A(new_n345), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(KEYINPUT71), .A3(new_n351), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  NOR3_X1   g158(.A1(new_n339), .A2(new_n343), .A3(new_n359), .ZN(new_n360));
  AOI211_X1 g159(.A(new_n353), .B(new_n352), .C1(new_n332), .C2(new_n338), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT37), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT38), .ZN(new_n363));
  XNOR2_X1  g162(.A(G8gat), .B(G36gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(KEYINPUT73), .ZN(new_n365));
  XNOR2_X1  g164(.A(G64gat), .B(G92gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n359), .B1(new_n339), .B2(new_n343), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n337), .B1(new_n336), .B2(new_n341), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n331), .A2(new_n288), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n352), .A2(new_n353), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT79), .B(KEYINPUT37), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n369), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n362), .A2(new_n363), .A3(new_n368), .A4(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(KEYINPUT6), .B(new_n208), .C1(new_n273), .C2(new_n278), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n369), .A2(new_n367), .A3(new_n374), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n287), .A2(new_n377), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n376), .A2(new_n368), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n340), .B1(new_n370), .B2(new_n371), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n332), .A2(KEYINPUT72), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n382), .A2(new_n383), .B1(new_n358), .B2(new_n354), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT37), .B1(new_n384), .B2(new_n373), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n363), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G78gat), .B(G106gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(G22gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G228gat), .ZN(new_n391));
  INV_X1    g190(.A(G233gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n354), .A2(new_n358), .B1(new_n341), .B2(new_n254), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n341), .B1(new_n352), .B2(new_n353), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n257), .B1(new_n395), .B2(new_n253), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n393), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT29), .B1(new_n357), .B2(new_n351), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n243), .B1(new_n398), .B2(KEYINPUT3), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n254), .A2(new_n341), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n372), .ZN(new_n401));
  INV_X1    g200(.A(new_n393), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT31), .B(G50gat), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n397), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n405), .B1(new_n397), .B2(new_n403), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n390), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n408), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n410), .A2(new_n389), .A3(new_n406), .ZN(new_n411));
  AND2_X1   g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT30), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n379), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n368), .B1(new_n384), .B2(new_n373), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n369), .A2(new_n374), .A3(KEYINPUT30), .A4(new_n367), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n254), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n253), .B1(new_n232), .B2(new_n242), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n418), .A2(new_n419), .A3(new_n265), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n248), .B1(new_n277), .B2(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n421), .B(KEYINPUT39), .C1(new_n248), .C2(new_n246), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT39), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n423), .B(new_n248), .C1(new_n277), .C2(new_n420), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n424), .A2(KEYINPUT78), .A3(new_n207), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT78), .B1(new_n424), .B2(new_n207), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n422), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT40), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI211_X1 g228(.A(KEYINPUT40), .B(new_n422), .C1(new_n425), .C2(new_n426), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n279), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n412), .B1(new_n417), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n202), .B1(new_n387), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n409), .A2(new_n411), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n429), .A2(new_n279), .A3(new_n430), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n437), .B(KEYINPUT80), .C1(new_n386), .C2(new_n380), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n436), .B1(new_n378), .B2(new_n287), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n440), .A2(new_n412), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n336), .A2(new_n265), .ZN(new_n442));
  NAND2_X1  g241(.A1(G227gat), .A2(G233gat), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n305), .A2(new_n316), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n445), .A2(new_n225), .A3(new_n333), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n442), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G15gat), .B(G43gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(G71gat), .B(G99gat), .ZN(new_n449));
  XOR2_X1   g248(.A(new_n448), .B(new_n449), .Z(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT33), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n447), .A2(KEYINPUT32), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT66), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n447), .A2(KEYINPUT66), .A3(KEYINPUT32), .A4(new_n451), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n447), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n450), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n458), .B1(new_n447), .B2(KEYINPUT32), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n454), .A2(new_n455), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n446), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT34), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n462), .A3(new_n443), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT68), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT68), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n461), .A2(new_n465), .A3(new_n462), .A4(new_n443), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n461), .A2(new_n443), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT34), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n464), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n460), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n464), .A2(new_n466), .A3(new_n468), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT67), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n471), .B1(new_n460), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n454), .A2(new_n455), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n457), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n474), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  OAI211_X1 g275(.A(KEYINPUT36), .B(new_n470), .C1(new_n473), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT69), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n474), .A2(new_n475), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT67), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n460), .A2(new_n472), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(new_n471), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT69), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT36), .A4(new_n470), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n479), .A2(new_n471), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n470), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT70), .B(KEYINPUT36), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n441), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n439), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n434), .B1(new_n460), .B2(new_n469), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n287), .A2(new_n378), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n482), .A2(new_n492), .A3(new_n493), .A4(new_n417), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT35), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT82), .ZN(new_n496));
  XOR2_X1   g295(.A(KEYINPUT81), .B(KEYINPUT35), .Z(new_n497));
  NAND4_X1  g296(.A1(new_n486), .A2(new_n412), .A3(new_n470), .A4(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n496), .B1(new_n499), .B2(new_n440), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n493), .A2(new_n417), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n501), .A2(KEYINPUT82), .A3(new_n498), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n495), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n491), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT15), .ZN(new_n505));
  OR2_X1    g304(.A1(G43gat), .A2(G50gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(G43gat), .A2(G50gat), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(KEYINPUT83), .B(G43gat), .Z(new_n509));
  INV_X1    g308(.A(G50gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n511), .A2(new_n505), .A3(new_n507), .ZN(new_n512));
  INV_X1    g311(.A(G36gat), .ZN(new_n513));
  AND2_X1   g312(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(G29gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n508), .B1(new_n512), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n519), .A2(new_n508), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT17), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT84), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525));
  INV_X1    g324(.A(G1gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(KEYINPUT16), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(new_n526), .B2(new_n525), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n524), .B1(new_n528), .B2(KEYINPUT85), .ZN(new_n529));
  INV_X1    g328(.A(G8gat), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n530), .B1(new_n528), .B2(new_n524), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(G8gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT86), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n532), .A2(KEYINPUT86), .A3(new_n533), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n523), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G229gat), .A2(G233gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n534), .A2(new_n522), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT18), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n534), .B(new_n522), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n539), .B(KEYINPUT13), .Z(new_n544));
  AOI22_X1  g343(.A1(new_n541), .A2(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n538), .A2(KEYINPUT18), .A3(new_n539), .A4(new_n540), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n546), .A2(KEYINPUT87), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(KEYINPUT87), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G113gat), .B(G141gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(G197gat), .ZN(new_n551));
  XOR2_X1   g350(.A(KEYINPUT11), .B(G169gat), .Z(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(KEYINPUT12), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n554), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n556), .B(new_n545), .C1(new_n547), .C2(new_n548), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n504), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT88), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT88), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n562), .B1(new_n504), .B2(new_n559), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n493), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT95), .ZN(new_n566));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT91), .ZN(new_n568));
  XOR2_X1   g367(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n569));
  XOR2_X1   g368(.A(new_n568), .B(new_n569), .Z(new_n570));
  AND2_X1   g369(.A1(G71gat), .A2(G78gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(G57gat), .B(G64gat), .Z(new_n574));
  AOI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(KEYINPUT89), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n574), .B1(KEYINPUT9), .B2(new_n571), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI221_X1 g376(.A(new_n574), .B1(KEYINPUT9), .B2(new_n571), .C1(new_n573), .C2(KEYINPUT89), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT90), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n578), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT90), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT92), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n580), .A2(KEYINPUT92), .A3(new_n583), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(KEYINPUT21), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT93), .ZN(new_n589));
  INV_X1    g388(.A(new_n534), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n589), .B1(new_n588), .B2(new_n590), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n570), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  INV_X1    g394(.A(new_n570), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(new_n591), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT21), .B1(new_n580), .B2(new_n583), .ZN(new_n599));
  XNOR2_X1  g398(.A(G127gat), .B(G155gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G183gat), .B(G211gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n598), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n594), .A2(new_n597), .A3(new_n603), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(G232gat), .A2(G233gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(KEYINPUT41), .ZN(new_n609));
  XNOR2_X1  g408(.A(G134gat), .B(G162gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT94), .B(KEYINPUT7), .ZN(new_n613));
  INV_X1    g412(.A(G85gat), .ZN(new_n614));
  INV_X1    g413(.A(G92gat), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g417(.A1(G99gat), .A2(G106gat), .ZN(new_n619));
  AOI22_X1  g418(.A1(KEYINPUT8), .A2(new_n619), .B1(new_n614), .B2(new_n615), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G99gat), .B(G106gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n621), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n523), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n621), .B(new_n622), .ZN(new_n626));
  AOI22_X1  g425(.A1(new_n626), .A2(new_n522), .B1(KEYINPUT41), .B2(new_n608), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(G190gat), .B(G218gat), .Z(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n628), .A2(new_n629), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n612), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n632), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(new_n611), .A3(new_n630), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n566), .B1(new_n607), .B2(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n605), .A2(new_n636), .A3(KEYINPUT95), .A4(new_n606), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n586), .A2(KEYINPUT10), .A3(new_n587), .A4(new_n626), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT96), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n624), .A2(new_n580), .A3(new_n583), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n579), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AOI211_X1 g446(.A(KEYINPUT96), .B(KEYINPUT10), .C1(new_n643), .C2(new_n644), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n641), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(G230gat), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(new_n392), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n645), .A2(new_n652), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT97), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n657), .B(new_n658), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n656), .B(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n640), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n564), .A2(new_n565), .A3(new_n662), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n663), .A2(KEYINPUT99), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(KEYINPUT99), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT98), .B(G1gat), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n664), .A2(new_n665), .A3(new_n667), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(G1324gat));
  NAND2_X1  g470(.A1(new_n564), .A2(new_n662), .ZN(new_n672));
  OAI21_X1  g471(.A(G8gat), .B1(new_n672), .B2(new_n417), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT42), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT16), .B(G8gat), .Z(new_n675));
  NAND4_X1  g474(.A1(new_n564), .A2(new_n436), .A3(new_n662), .A4(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT100), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n676), .A2(new_n677), .A3(new_n674), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n677), .B1(new_n676), .B2(new_n674), .ZN(new_n679));
  OAI221_X1 g478(.A(new_n673), .B1(new_n674), .B2(new_n676), .C1(new_n678), .C2(new_n679), .ZN(G1325gat));
  OR3_X1    g479(.A1(new_n672), .A2(G15gat), .A3(new_n487), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n485), .A2(new_n489), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(G15gat), .B1(new_n672), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n684), .ZN(G1326gat));
  NAND3_X1  g484(.A1(new_n564), .A2(new_n434), .A3(new_n662), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n686), .A2(KEYINPUT101), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(KEYINPUT101), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT43), .B(G22gat), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n687), .A2(new_n688), .A3(new_n690), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(G1327gat));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT82), .B1(new_n501), .B2(new_n498), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n499), .A2(new_n440), .A3(new_n496), .ZN(new_n697));
  AOI221_X4 g496(.A(new_n695), .B1(new_n494), .B2(KEYINPUT35), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT103), .B1(new_n699), .B2(new_n495), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n491), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT104), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n491), .B(new_n703), .C1(new_n698), .C2(new_n700), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n636), .A2(KEYINPUT44), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n702), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT44), .B1(new_n504), .B2(new_n636), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n607), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n559), .A2(new_n661), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(G29gat), .B1(new_n711), .B2(new_n493), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n661), .A2(new_n709), .A3(new_n636), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n493), .A2(G29gat), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n564), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT102), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT102), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n564), .A2(new_n718), .A3(new_n713), .A4(new_n714), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n717), .B1(new_n716), .B2(new_n719), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n712), .B1(new_n720), .B2(new_n721), .ZN(G1328gat));
  NAND2_X1  g521(.A1(new_n564), .A2(new_n713), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n436), .A2(new_n513), .ZN(new_n724));
  OR3_X1    g523(.A1(new_n723), .A2(KEYINPUT46), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G36gat), .B1(new_n711), .B2(new_n417), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT46), .B1(new_n723), .B2(new_n724), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(G1329gat));
  OR3_X1    g527(.A1(new_n711), .A2(new_n683), .A3(new_n509), .ZN(new_n729));
  OR2_X1    g528(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n730));
  INV_X1    g529(.A(new_n487), .ZN(new_n731));
  INV_X1    g530(.A(new_n563), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n504), .A2(new_n562), .A3(new_n559), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n731), .B(new_n713), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n734), .A2(new_n509), .B1(KEYINPUT105), .B2(KEYINPUT47), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n729), .A2(new_n730), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n730), .B1(new_n729), .B2(new_n735), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(G1330gat));
  OAI21_X1  g537(.A(G50gat), .B1(new_n711), .B2(new_n412), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n564), .A2(new_n510), .A3(new_n434), .A4(new_n713), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT48), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1331gat));
  NOR3_X1   g542(.A1(new_n640), .A2(new_n558), .A3(new_n660), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n702), .A2(new_n704), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(new_n493), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT106), .B(G57gat), .Z(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1332gat));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n745), .A2(new_n749), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n417), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT108), .ZN(new_n754));
  NOR2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n750), .A2(new_n756), .A3(new_n751), .A4(new_n752), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n755), .B1(new_n754), .B2(new_n757), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(G1333gat));
  NAND4_X1  g559(.A1(new_n750), .A2(G71gat), .A3(new_n682), .A4(new_n751), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n487), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(G71gat), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT50), .ZN(G1334gat));
  NAND3_X1  g563(.A1(new_n750), .A2(new_n434), .A3(new_n751), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g565(.A1(new_n709), .A2(new_n558), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n661), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n708), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G85gat), .B1(new_n770), .B2(new_n493), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n503), .A2(new_n695), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n699), .A2(KEYINPUT103), .A3(new_n495), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n772), .A2(new_n773), .B1(new_n439), .B2(new_n490), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n767), .A2(new_n637), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT51), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n775), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n701), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n661), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n565), .A2(new_n614), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n771), .B1(new_n781), .B2(new_n782), .ZN(G1336gat));
  NOR3_X1   g582(.A1(new_n660), .A2(G92gat), .A3(new_n417), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT52), .B1(new_n780), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n770), .A2(new_n417), .ZN(new_n786));
  OAI21_X1  g585(.A(G92gat), .B1(new_n786), .B2(KEYINPUT111), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n770), .A2(new_n788), .A3(new_n417), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n785), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n786), .A2(new_n615), .ZN(new_n791));
  XOR2_X1   g590(.A(new_n784), .B(KEYINPUT109), .Z(new_n792));
  OAI211_X1 g591(.A(KEYINPUT110), .B(new_n778), .C1(new_n774), .C2(new_n775), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT110), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n701), .A2(new_n777), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n792), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT52), .B1(new_n791), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n790), .A2(new_n797), .ZN(G1337gat));
  INV_X1    g597(.A(G99gat), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n780), .A2(new_n799), .A3(new_n731), .A4(new_n661), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n770), .A2(new_n683), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n801), .B2(new_n799), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT112), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n804), .B(new_n800), .C1(new_n801), .C2(new_n799), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(G1338gat));
  NOR2_X1   g605(.A1(new_n412), .A2(G106gat), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n776), .A2(new_n661), .A3(new_n779), .A4(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI211_X1 g609(.A(new_n412), .B(new_n768), .C1(new_n706), .C2(new_n707), .ZN(new_n811));
  XNOR2_X1  g610(.A(KEYINPUT113), .B(G106gat), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n661), .A2(new_n807), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n793), .B2(new_n795), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n708), .A2(new_n434), .A3(new_n769), .ZN(new_n816));
  INV_X1    g615(.A(new_n812), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n813), .B1(new_n818), .B2(new_n809), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n813), .B(KEYINPUT114), .C1(new_n818), .C2(new_n809), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(G1339gat));
  AND4_X1   g622(.A1(new_n559), .A2(new_n638), .A3(new_n639), .A4(new_n660), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n539), .B1(new_n538), .B2(new_n540), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n543), .A2(new_n544), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n553), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n557), .A2(new_n827), .ZN(new_n828));
  OR3_X1    g627(.A1(new_n660), .A2(new_n828), .A3(new_n637), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n637), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n555), .A2(new_n557), .A3(new_n636), .ZN(new_n831));
  INV_X1    g630(.A(new_n659), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n656), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n651), .B(new_n641), .C1(new_n647), .C2(new_n648), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n653), .A2(KEYINPUT54), .A3(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n649), .A2(new_n836), .A3(new_n652), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n835), .A2(new_n832), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n833), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n830), .A2(new_n831), .A3(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n835), .A2(KEYINPUT55), .A3(new_n832), .A4(new_n837), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT115), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n829), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n824), .B1(new_n844), .B2(new_n607), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n493), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n482), .A2(new_n492), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(new_n417), .A3(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n214), .A3(new_n558), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n845), .A2(new_n434), .A3(new_n487), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n493), .A2(new_n436), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT116), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n855), .A2(new_n558), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n851), .B1(new_n856), .B2(new_n210), .ZN(G1340gat));
  AOI21_X1  g656(.A(G120gat), .B1(new_n850), .B2(new_n661), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n660), .A2(new_n211), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n858), .B1(new_n855), .B2(new_n859), .ZN(G1341gat));
  NAND3_X1  g659(.A1(new_n850), .A2(new_n218), .A3(new_n709), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n855), .A2(new_n709), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n861), .B1(new_n862), .B2(new_n218), .ZN(G1342gat));
  NOR2_X1   g662(.A1(new_n636), .A2(new_n436), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT117), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT56), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n865), .B(new_n216), .C1(KEYINPUT118), .C2(new_n866), .ZN(new_n867));
  NOR4_X1   g666(.A1(new_n845), .A2(new_n493), .A3(new_n847), .A4(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(KEYINPUT118), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n868), .B(new_n869), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n855), .A2(new_n637), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n216), .ZN(G1343gat));
  NAND2_X1  g671(.A1(new_n683), .A2(new_n853), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n844), .A2(new_n607), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(KEYINPUT119), .ZN(new_n875));
  INV_X1    g674(.A(new_n824), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n844), .A2(new_n607), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI211_X1 g678(.A(KEYINPUT57), .B(new_n434), .C1(new_n875), .C2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n881), .B1(new_n845), .B2(new_n412), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n873), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(G141gat), .A3(new_n558), .ZN(new_n884));
  NAND2_X1  g683(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n885));
  NOR2_X1   g684(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n682), .A2(new_n412), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n846), .A2(new_n417), .A3(new_n558), .A4(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n886), .B1(new_n888), .B2(new_n233), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n884), .A2(new_n885), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n885), .B1(new_n884), .B2(new_n889), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n890), .A2(new_n891), .ZN(G1344gat));
  NAND2_X1  g691(.A1(new_n846), .A2(new_n887), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n436), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n235), .A3(new_n661), .ZN(new_n895));
  AOI211_X1 g694(.A(KEYINPUT59), .B(new_n235), .C1(new_n883), .C2(new_n661), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n873), .A2(new_n660), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n877), .A2(new_n876), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT57), .B1(new_n899), .B2(new_n434), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n845), .A2(new_n881), .A3(new_n412), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n897), .B1(new_n902), .B2(G148gat), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n895), .B1(new_n896), .B2(new_n903), .ZN(G1345gat));
  INV_X1    g703(.A(new_n883), .ZN(new_n905));
  OAI21_X1  g704(.A(G155gat), .B1(new_n905), .B2(new_n607), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n894), .A2(new_n239), .A3(new_n709), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1346gat));
  OAI21_X1  g707(.A(G162gat), .B1(new_n905), .B2(new_n636), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n865), .A2(new_n240), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n893), .B2(new_n910), .ZN(G1347gat));
  NOR2_X1   g710(.A1(new_n565), .A2(new_n417), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n852), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(G169gat), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n913), .A2(new_n914), .A3(new_n559), .ZN(new_n915));
  NOR4_X1   g714(.A1(new_n845), .A2(new_n565), .A3(new_n417), .A4(new_n847), .ZN(new_n916));
  AOI21_X1  g715(.A(G169gat), .B1(new_n916), .B2(new_n558), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n915), .A2(new_n917), .ZN(G1348gat));
  OAI21_X1  g717(.A(G176gat), .B1(new_n913), .B2(new_n660), .ZN(new_n919));
  INV_X1    g718(.A(G176gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n916), .A2(new_n920), .A3(new_n661), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1349gat));
  OAI21_X1  g721(.A(G183gat), .B1(new_n913), .B2(new_n607), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n916), .A2(new_n323), .A3(new_n709), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT60), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n926), .A2(KEYINPUT121), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n925), .B(new_n927), .ZN(G1350gat));
  OAI21_X1  g727(.A(G190gat), .B1(new_n913), .B2(new_n636), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT61), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n916), .A2(new_n296), .A3(new_n637), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT122), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(G1351gat));
  NAND2_X1  g732(.A1(new_n887), .A2(new_n436), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT123), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n845), .A2(new_n565), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  XOR2_X1   g737(.A(KEYINPUT124), .B(G197gat), .Z(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n558), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n683), .A2(new_n912), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n899), .A2(KEYINPUT57), .A3(new_n434), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(new_n882), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n944), .A2(new_n559), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n940), .B1(new_n945), .B2(new_n939), .ZN(G1352gat));
  NOR3_X1   g745(.A1(new_n937), .A2(G204gat), .A3(new_n660), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT62), .ZN(new_n948));
  OAI21_X1  g747(.A(G204gat), .B1(new_n944), .B2(new_n660), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1353gat));
  AOI21_X1  g749(.A(new_n348), .B1(new_n943), .B2(new_n709), .ZN(new_n951));
  OAI21_X1  g750(.A(KEYINPUT126), .B1(new_n951), .B2(KEYINPUT63), .ZN(new_n952));
  INV_X1    g751(.A(new_n941), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n709), .B(new_n953), .C1(new_n900), .C2(new_n901), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n954), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(KEYINPUT125), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT63), .ZN(new_n958));
  AOI211_X1 g757(.A(new_n607), .B(new_n941), .C1(new_n942), .C2(new_n882), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n957), .B(new_n958), .C1(new_n959), .C2(new_n348), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n954), .A2(new_n961), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n952), .A2(new_n956), .A3(new_n960), .A4(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n938), .A2(new_n348), .A3(new_n709), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1354gat));
  OAI21_X1  g764(.A(G218gat), .B1(new_n944), .B2(new_n636), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n938), .A2(new_n349), .A3(new_n637), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(G1355gat));
endmodule


