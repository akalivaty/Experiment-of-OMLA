//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n808, new_n810, new_n811, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939;
  INV_X1    g000(.A(G64gat), .ZN(new_n202));
  AND2_X1   g001(.A1(new_n202), .A2(G57gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(G57gat), .ZN(new_n204));
  INV_X1    g003(.A(G71gat), .ZN(new_n205));
  INV_X1    g004(.A(G78gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI22_X1  g006(.A1(new_n203), .A2(new_n204), .B1(new_n207), .B2(KEYINPUT9), .ZN(new_n208));
  XOR2_X1   g007(.A(G71gat), .B(G78gat), .Z(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n211), .A2(KEYINPUT21), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n213));
  XOR2_X1   g012(.A(new_n212), .B(new_n213), .Z(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n210), .B(KEYINPUT97), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT21), .ZN(new_n217));
  INV_X1    g016(.A(G183gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(G15gat), .B(G22gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT16), .ZN(new_n220));
  AOI21_X1  g019(.A(G1gat), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(G8gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(KEYINPUT95), .ZN(new_n223));
  XOR2_X1   g022(.A(new_n222), .B(new_n223), .Z(new_n224));
  AND3_X1   g023(.A1(new_n217), .A2(new_n218), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n218), .B1(new_n217), .B2(new_n224), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(G231gat), .A3(G233gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(G231gat), .A2(G233gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(new_n225), .B2(new_n226), .ZN(new_n230));
  XNOR2_X1  g029(.A(G127gat), .B(G155gat), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n231), .B(G211gat), .Z(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n228), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n233), .B1(new_n228), .B2(new_n230), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n215), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n236), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(new_n214), .A3(new_n234), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G99gat), .A2(G106gat), .ZN(new_n241));
  INV_X1    g040(.A(G85gat), .ZN(new_n242));
  INV_X1    g041(.A(G92gat), .ZN(new_n243));
  AOI22_X1  g042(.A1(KEYINPUT8), .A2(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(new_n242), .B2(new_n243), .ZN(new_n246));
  NAND4_X1  g045(.A1(KEYINPUT98), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n244), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(G99gat), .B(G106gat), .Z(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G43gat), .B(G50gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT93), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT15), .ZN(new_n254));
  OR2_X1    g053(.A1(new_n252), .A2(KEYINPUT15), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT14), .ZN(new_n257));
  OR3_X1    g056(.A1(new_n257), .A2(G29gat), .A3(G36gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n257), .B1(G29gat), .B2(G36gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(G29gat), .A2(G36gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(KEYINPUT94), .A2(KEYINPUT17), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n262), .B1(new_n253), .B2(KEYINPUT15), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT94), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT17), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n263), .A2(new_n264), .A3(new_n266), .A4(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n261), .B1(new_n254), .B2(new_n255), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n267), .B(new_n268), .C1(new_n271), .C2(new_n265), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n251), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G232gat), .A2(G233gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT41), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n263), .A2(new_n266), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n277), .A2(new_n250), .ZN(new_n278));
  OR3_X1    g077(.A1(new_n273), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(G190gat), .B(G218gat), .Z(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT99), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n274), .A2(new_n275), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n279), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NOR3_X1   g085(.A1(new_n273), .A2(new_n276), .A3(new_n278), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n275), .B(new_n274), .C1(new_n287), .C2(new_n283), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n281), .A2(new_n282), .ZN(new_n290));
  XOR2_X1   g089(.A(G134gat), .B(G162gat), .Z(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n286), .A2(new_n288), .A3(new_n292), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n240), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n270), .A2(new_n272), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n224), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n224), .A2(new_n277), .ZN(new_n300));
  NAND2_X1  g099(.A1(G229gat), .A2(G233gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT18), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n224), .B(new_n277), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n301), .B(KEYINPUT13), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n299), .A2(new_n300), .A3(KEYINPUT18), .A4(new_n301), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n304), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n311), .B(G197gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(G113gat), .B(G141gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT92), .B(G169gat), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n314), .B(new_n315), .Z(new_n316));
  INV_X1    g115(.A(KEYINPUT12), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n310), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n304), .A2(new_n308), .A3(new_n309), .A4(new_n318), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(KEYINPUT96), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT96), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n310), .A2(new_n323), .A3(new_n319), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G176gat), .B(G204gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT103), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(G120gat), .ZN(new_n329));
  INV_X1    g128(.A(G148gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n250), .A2(KEYINPUT100), .ZN(new_n332));
  OR2_X1    g131(.A1(new_n248), .A2(new_n249), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT100), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n248), .A2(new_n249), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n332), .A2(new_n210), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n211), .A2(KEYINPUT100), .A3(new_n250), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(KEYINPUT101), .A2(KEYINPUT10), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT101), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT10), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n339), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n216), .A2(KEYINPUT10), .A3(new_n251), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G230gat), .ZN(new_n347));
  INV_X1    g146(.A(G233gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n339), .A2(new_n350), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n331), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT104), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT102), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n356), .B1(new_n346), .B2(new_n350), .ZN(new_n357));
  AOI211_X1 g156(.A(KEYINPUT102), .B(new_n349), .C1(new_n344), .C2(new_n345), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n331), .B(new_n353), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n326), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT27), .B(G183gat), .ZN(new_n363));
  INV_X1    g162(.A(G190gat), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(KEYINPUT28), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT67), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT27), .B1(new_n366), .B2(new_n218), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT27), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n368), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n367), .A2(new_n364), .A3(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n365), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G169gat), .ZN(new_n373));
  INV_X1    g172(.A(G176gat), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT69), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT69), .A4(KEYINPUT26), .ZN(new_n378));
  NAND2_X1  g177(.A1(G183gat), .A2(G190gat), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n372), .A2(new_n377), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT24), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n218), .A2(new_n364), .A3(KEYINPUT65), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT65), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n384), .B1(G183gat), .B2(G190gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n382), .A2(new_n383), .A3(new_n385), .A4(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT23), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n388), .A2(new_n373), .A3(new_n374), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n389), .A2(new_n390), .B1(G169gat), .B2(G176gat), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT25), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n387), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT66), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n386), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n218), .A2(new_n364), .ZN(new_n396));
  NAND4_X1  g195(.A1(KEYINPUT66), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n395), .A2(new_n396), .A3(new_n382), .A4(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n392), .B1(new_n398), .B2(new_n391), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n380), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT71), .ZN(new_n402));
  INV_X1    g201(.A(G120gat), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n402), .B1(new_n403), .B2(G113gat), .ZN(new_n404));
  INV_X1    g203(.A(G113gat), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT70), .B1(new_n405), .B2(G120gat), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT70), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(new_n403), .A3(G113gat), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n405), .A2(KEYINPUT71), .A3(G120gat), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n404), .A2(new_n406), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  OR2_X1    g209(.A1(G127gat), .A2(G134gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(G127gat), .A2(G134gat), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT1), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT72), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n410), .A2(KEYINPUT72), .A3(new_n413), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G113gat), .B(G120gat), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n419), .A2(KEYINPUT1), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n411), .A2(new_n412), .ZN(new_n421));
  OR2_X1    g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n401), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n420), .A2(new_n421), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n425), .B1(new_n416), .B2(new_n417), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n426), .A2(new_n380), .A3(new_n400), .ZN(new_n427));
  NAND2_X1  g226(.A1(G227gat), .A2(G233gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT34), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n424), .A2(new_n427), .ZN(new_n431));
  XOR2_X1   g230(.A(new_n428), .B(KEYINPUT64), .Z(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(KEYINPUT34), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n430), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n432), .B1(new_n424), .B2(new_n427), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT32), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  OAI221_X1 g239(.A(new_n430), .B1(new_n431), .B2(new_n435), .C1(new_n438), .C2(new_n437), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n437), .A2(KEYINPUT33), .ZN(new_n442));
  XNOR2_X1  g241(.A(G71gat), .B(G99gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(KEYINPUT73), .ZN(new_n444));
  XNOR2_X1  g243(.A(G15gat), .B(G43gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n440), .A2(new_n441), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n447), .B1(new_n440), .B2(new_n441), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT31), .B(G50gat), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(G228gat), .A2(G233gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n453), .B(KEYINPUT81), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT83), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n330), .A2(G141gat), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(KEYINPUT76), .B(G148gat), .ZN(new_n458));
  INV_X1    g257(.A(G141gat), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(KEYINPUT77), .A2(G155gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT2), .ZN(new_n462));
  INV_X1    g261(.A(G162gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(G155gat), .ZN(new_n464));
  INV_X1    g263(.A(G155gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(G162gat), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n462), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT2), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n459), .A2(G148gat), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n468), .B1(new_n456), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n464), .A2(new_n466), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n460), .A2(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(G211gat), .B(G218gat), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  XOR2_X1   g273(.A(G197gat), .B(G204gat), .Z(new_n475));
  AOI21_X1  g274(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OR2_X1    g276(.A1(G197gat), .A2(G204gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(G197gat), .A2(G204gat), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n473), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n477), .A2(KEYINPUT75), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT29), .ZN(new_n483));
  OR3_X1    g282(.A1(new_n480), .A2(KEYINPUT75), .A3(new_n473), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT3), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n472), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n455), .B1(new_n487), .B2(new_n453), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n486), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n483), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n482), .A2(new_n484), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT83), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n490), .A2(new_n494), .A3(new_n491), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n470), .A2(new_n471), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n462), .A2(new_n464), .A3(new_n466), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n330), .A2(KEYINPUT76), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n330), .A2(KEYINPUT76), .ZN(new_n500));
  OAI21_X1  g299(.A(G141gat), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n498), .B1(new_n501), .B2(new_n457), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT78), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT78), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n472), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT82), .B1(new_n480), .B2(new_n473), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT29), .B1(new_n507), .B2(new_n477), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n474), .B(KEYINPUT82), .C1(new_n475), .C2(new_n476), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT3), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n454), .B1(new_n495), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n493), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT84), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT84), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n493), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G78gat), .B(G106gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(G22gat), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n514), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n519), .B1(new_n514), .B2(new_n516), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n452), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n514), .A2(new_n516), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n518), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n514), .A2(new_n516), .A3(new_n519), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n525), .A3(new_n451), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n450), .A2(new_n522), .A3(new_n526), .ZN(new_n527));
  AND2_X1   g326(.A1(G226gat), .A2(G233gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n401), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT29), .B1(new_n380), .B2(new_n400), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n491), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n529), .B(new_n491), .C1(new_n528), .C2(new_n530), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G8gat), .B(G36gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(new_n202), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(new_n243), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n533), .A2(new_n538), .A3(new_n534), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(KEYINPUT30), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n535), .A2(new_n543), .A3(new_n539), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G225gat), .A2(G233gat), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n472), .B1(new_n418), .B2(new_n422), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n410), .A2(KEYINPUT72), .A3(new_n413), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT72), .B1(new_n410), .B2(new_n413), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n472), .B(new_n422), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n547), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT79), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n506), .A2(KEYINPUT4), .A3(new_n426), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT3), .B1(new_n502), .B2(new_n497), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n423), .A2(new_n489), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT4), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n547), .B1(new_n551), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n555), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT79), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n561), .B(new_n547), .C1(new_n548), .C2(new_n552), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n554), .A2(KEYINPUT5), .A3(new_n560), .A4(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT0), .B(G57gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(G85gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(G1gat), .B(G29gat), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n565), .B(new_n566), .Z(new_n567));
  NOR2_X1   g366(.A1(new_n551), .A2(new_n558), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n547), .A2(KEYINPUT5), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n556), .A2(new_n489), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n558), .B1(new_n571), .B2(new_n423), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n506), .A2(new_n426), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n569), .B(new_n570), .C1(new_n572), .C2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n563), .A2(new_n567), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT6), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n567), .B1(new_n563), .B2(new_n575), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n575), .ZN(new_n581));
  INV_X1    g380(.A(new_n567), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(KEYINPUT6), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n545), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT80), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n581), .A2(new_n582), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(new_n577), .A3(new_n576), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n583), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n590), .A2(KEYINPUT80), .A3(new_n545), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n527), .B1(new_n587), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT35), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT90), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n450), .A2(new_n522), .A3(new_n526), .ZN(new_n595));
  AOI221_X4 g394(.A(new_n586), .B1(new_n542), .B2(new_n544), .C1(new_n589), .C2(new_n583), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT80), .B1(new_n590), .B2(new_n545), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT90), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(new_n599), .A3(KEYINPUT35), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT88), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(KEYINPUT89), .B(KEYINPUT35), .Z(new_n603));
  NAND3_X1  g402(.A1(new_n590), .A2(KEYINPUT88), .A3(new_n545), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n595), .A2(new_n602), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n594), .A2(new_n600), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n533), .A2(KEYINPUT37), .A3(new_n534), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT86), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT86), .A4(KEYINPUT37), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n539), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT38), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT37), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n535), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n611), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n615), .A2(new_n583), .A3(new_n589), .A4(new_n540), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT87), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n580), .A2(new_n584), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT87), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n618), .A2(new_n619), .A3(new_n540), .A4(new_n615), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n614), .A2(new_n538), .A3(new_n607), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT38), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n569), .B1(new_n572), .B2(new_n574), .ZN(new_n624));
  XOR2_X1   g423(.A(KEYINPUT85), .B(KEYINPUT39), .Z(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n547), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n557), .A2(KEYINPUT4), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n568), .B1(new_n627), .B2(new_n573), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT39), .B1(new_n628), .B2(new_n546), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n548), .A2(new_n552), .A3(new_n547), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n567), .B(new_n626), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT40), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NOR4_X1   g433(.A1(new_n633), .A2(new_n634), .A3(new_n545), .A4(new_n579), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n522), .A2(new_n526), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n623), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n587), .A2(new_n591), .A3(new_n636), .ZN(new_n639));
  INV_X1    g438(.A(new_n450), .ZN(new_n640));
  NAND2_X1  g439(.A1(KEYINPUT74), .A2(KEYINPUT36), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n643));
  OAI21_X1  g442(.A(new_n642), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n638), .A2(new_n639), .A3(new_n644), .ZN(new_n645));
  AOI211_X1 g444(.A(new_n297), .B(new_n362), .C1(new_n606), .C2(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n646), .A2(KEYINPUT105), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(KEYINPUT105), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n618), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(G1gat), .ZN(G1324gat));
  INV_X1    g451(.A(KEYINPUT106), .ZN(new_n653));
  INV_X1    g452(.A(new_n545), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n654), .B1(new_n647), .B2(new_n648), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT16), .B(G8gat), .Z(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n653), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT42), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT42), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n653), .B(new_n660), .C1(new_n655), .C2(new_n657), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT107), .B1(new_n655), .B2(G8gat), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n655), .A2(KEYINPUT107), .A3(G8gat), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n659), .B(new_n661), .C1(new_n662), .C2(new_n663), .ZN(G1325gat));
  AOI21_X1  g463(.A(G15gat), .B1(new_n650), .B2(new_n450), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n649), .A2(new_n644), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n665), .B1(G15gat), .B2(new_n666), .ZN(G1326gat));
  INV_X1    g466(.A(new_n636), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n649), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT43), .B(G22gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  AOI21_X1  g470(.A(new_n296), .B1(new_n606), .B2(new_n645), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n362), .A2(new_n240), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n674), .A2(G29gat), .A3(new_n590), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(KEYINPUT45), .Z(new_n676));
  NAND2_X1  g475(.A1(new_n606), .A2(new_n645), .ZN(new_n677));
  INV_X1    g476(.A(new_n296), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n680), .B1(new_n681), .B2(new_n672), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n618), .A3(new_n673), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(G29gat), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n676), .A2(new_n684), .ZN(G1328gat));
  NAND3_X1  g484(.A1(new_n682), .A2(new_n654), .A3(new_n673), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT109), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(G36gat), .A3(new_n689), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n674), .A2(G36gat), .A3(new_n545), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT46), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(G1329gat));
  NOR3_X1   g492(.A1(new_n674), .A2(G43gat), .A3(new_n640), .ZN(new_n694));
  INV_X1    g493(.A(new_n644), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n682), .A2(new_n695), .A3(new_n673), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n694), .B1(new_n696), .B2(G43gat), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT47), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n698), .A2(KEYINPUT110), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(KEYINPUT110), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n697), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n699), .B1(new_n697), .B2(new_n700), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(G1330gat));
  NAND4_X1  g502(.A1(new_n682), .A2(G50gat), .A3(new_n636), .A4(new_n673), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n674), .A2(new_n668), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(G50gat), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g506(.A(new_n360), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n297), .A2(new_n325), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n677), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n590), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT111), .B(G57gat), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1332gat));
  AOI211_X1 g512(.A(new_n545), .B(new_n710), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT112), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  OR2_X1    g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  OR3_X1    g517(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n716), .B2(new_n717), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(G1333gat));
  OAI21_X1  g520(.A(G71gat), .B1(new_n710), .B2(new_n644), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n677), .A2(new_n205), .A3(new_n709), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n640), .B2(new_n723), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n668), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(new_n206), .ZN(G1335gat));
  NAND2_X1  g526(.A1(new_n677), .A2(new_n678), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n325), .A2(new_n240), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  OR3_X1    g529(.A1(new_n728), .A2(KEYINPUT51), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT51), .B1(new_n728), .B2(new_n730), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n731), .A2(new_n618), .A3(new_n360), .A4(new_n732), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n733), .A2(new_n242), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n730), .A2(new_n708), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT113), .B1(new_n682), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n672), .A2(new_n681), .ZN(new_n738));
  INV_X1    g537(.A(new_n679), .ZN(new_n739));
  AOI211_X1 g538(.A(new_n296), .B(new_n739), .C1(new_n606), .C2(new_n645), .ZN(new_n740));
  OAI211_X1 g539(.A(KEYINPUT113), .B(new_n735), .C1(new_n738), .C2(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n590), .B1(new_n737), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n734), .B1(G85gat), .B2(new_n742), .ZN(G1336gat));
  NAND2_X1  g542(.A1(new_n682), .A2(new_n735), .ZN(new_n744));
  OAI21_X1  g543(.A(G92gat), .B1(new_n744), .B2(new_n545), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n545), .A2(G92gat), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n731), .A2(new_n360), .A3(new_n732), .A4(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n748), .ZN(new_n750));
  INV_X1    g549(.A(new_n741), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n654), .B1(new_n751), .B2(new_n736), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n750), .B1(new_n752), .B2(G92gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n749), .B1(new_n753), .B2(new_n746), .ZN(G1337gat));
  AND2_X1   g553(.A1(new_n731), .A2(new_n732), .ZN(new_n755));
  INV_X1    g554(.A(G99gat), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n755), .A2(new_n756), .A3(new_n450), .A4(new_n360), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n644), .B1(new_n737), .B2(new_n741), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n758), .B2(new_n756), .ZN(G1338gat));
  XOR2_X1   g558(.A(KEYINPUT114), .B(G106gat), .Z(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n744), .B2(new_n668), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n668), .A2(G106gat), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n731), .A2(new_n360), .A3(new_n732), .A4(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n761), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n764), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n636), .B1(new_n751), .B2(new_n736), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n766), .B1(new_n767), .B2(new_n760), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n765), .B1(new_n768), .B2(new_n762), .ZN(G1339gat));
  NOR3_X1   g568(.A1(new_n297), .A2(new_n325), .A3(new_n360), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n344), .A2(new_n349), .A3(new_n345), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n771), .B(KEYINPUT54), .C1(new_n357), .C2(new_n358), .ZN(new_n772));
  INV_X1    g571(.A(new_n351), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT54), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n331), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n772), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n776), .B1(new_n772), .B2(new_n775), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n359), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n299), .A2(new_n300), .ZN(new_n781));
  OAI22_X1  g580(.A1(new_n781), .A2(new_n301), .B1(new_n305), .B2(new_n307), .ZN(new_n782));
  INV_X1    g581(.A(new_n316), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n784), .A2(new_n321), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n785), .A2(new_n295), .A3(new_n294), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT115), .B1(new_n780), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n359), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n775), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT55), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n788), .B1(new_n790), .B2(new_n777), .ZN(new_n791));
  AND4_X1   g590(.A1(new_n295), .A2(new_n294), .A3(new_n321), .A4(new_n784), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n325), .A2(new_n791), .B1(new_n360), .B2(new_n785), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n787), .B(new_n794), .C1(new_n795), .C2(new_n678), .ZN(new_n796));
  INV_X1    g595(.A(new_n240), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n770), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n798), .A2(new_n590), .A3(new_n527), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n545), .ZN(new_n800));
  OAI21_X1  g599(.A(G113gat), .B1(new_n800), .B2(new_n326), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n325), .A2(new_n405), .ZN(new_n802));
  XOR2_X1   g601(.A(new_n802), .B(KEYINPUT116), .Z(new_n803));
  OAI21_X1  g602(.A(new_n801), .B1(new_n800), .B2(new_n803), .ZN(G1340gat));
  NOR2_X1   g603(.A1(new_n708), .A2(new_n654), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n799), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n360), .A2(new_n403), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT117), .ZN(new_n808));
  OAI22_X1  g607(.A1(new_n806), .A2(new_n403), .B1(new_n800), .B2(new_n808), .ZN(G1341gat));
  INV_X1    g608(.A(new_n800), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n240), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n678), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n814));
  XOR2_X1   g613(.A(KEYINPUT56), .B(G134gat), .Z(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n813), .B2(new_n815), .ZN(G1343gat));
  NAND2_X1  g615(.A1(new_n325), .A2(new_n791), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n360), .A2(new_n785), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n678), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n787), .A2(new_n794), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n797), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n770), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n668), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n823), .A2(new_n618), .A3(new_n545), .A4(new_n644), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n824), .A2(G141gat), .A3(new_n326), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT58), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(KEYINPUT57), .B1(new_n798), .B2(new_n668), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n644), .A2(new_n618), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n654), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n829), .A2(new_n830), .A3(new_n325), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(G141gat), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n827), .B(new_n834), .C1(new_n826), .C2(new_n825), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n833), .A2(new_n836), .A3(G141gat), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n833), .B2(G141gat), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n837), .A2(new_n838), .A3(new_n825), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT58), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n835), .B1(new_n839), .B2(new_n840), .ZN(G1344gat));
  INV_X1    g640(.A(new_n458), .ZN(new_n842));
  INV_X1    g641(.A(new_n831), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n823), .A2(new_n842), .A3(new_n805), .A4(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845));
  INV_X1    g644(.A(new_n819), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n791), .A2(new_n792), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n240), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n828), .B(new_n636), .C1(new_n848), .C2(new_n770), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n830), .A3(new_n360), .ZN(new_n850));
  INV_X1    g649(.A(new_n832), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n845), .B1(new_n852), .B2(G148gat), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n829), .A2(new_n830), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n854), .A2(new_n708), .A3(new_n851), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n855), .A2(KEYINPUT59), .A3(new_n842), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n844), .B1(new_n853), .B2(new_n856), .ZN(G1345gat));
  XNOR2_X1  g656(.A(KEYINPUT77), .B(G155gat), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n860), .B1(new_n824), .B2(new_n797), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n824), .A2(new_n860), .A3(new_n797), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR4_X1   g663(.A1(new_n854), .A2(new_n859), .A3(new_n797), .A4(new_n851), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(KEYINPUT121), .A3(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n868));
  INV_X1    g667(.A(new_n824), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(KEYINPUT120), .A3(new_n240), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n858), .B1(new_n870), .B2(new_n861), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n868), .B1(new_n871), .B2(new_n865), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n867), .A2(new_n872), .ZN(G1346gat));
  INV_X1    g672(.A(new_n854), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n678), .A3(new_n832), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT122), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n874), .A2(KEYINPUT122), .A3(new_n678), .A4(new_n832), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n877), .A2(G162gat), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n869), .A2(new_n463), .A3(new_n678), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1347gat));
  NAND2_X1  g680(.A1(new_n821), .A2(new_n822), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n618), .A2(new_n545), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(new_n595), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(G169gat), .B1(new_n884), .B2(new_n326), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n595), .A2(new_n654), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n886), .B(KEYINPUT123), .Z(new_n887));
  AOI211_X1 g686(.A(new_n618), .B(new_n887), .C1(new_n821), .C2(new_n822), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n373), .A3(new_n325), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n885), .A2(new_n889), .ZN(G1348gat));
  NOR3_X1   g689(.A1(new_n884), .A2(new_n374), .A3(new_n708), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n891), .A2(KEYINPUT124), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n891), .A2(KEYINPUT124), .ZN(new_n893));
  AOI21_X1  g692(.A(G176gat), .B1(new_n888), .B2(new_n360), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(G1349gat));
  NAND3_X1  g694(.A1(new_n888), .A2(new_n363), .A3(new_n240), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n884), .A2(new_n797), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(new_n218), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n296), .ZN(new_n900));
  OR3_X1    g699(.A1(new_n900), .A2(KEYINPUT125), .A3(new_n364), .ZN(new_n901));
  OAI21_X1  g700(.A(KEYINPUT125), .B1(new_n900), .B2(new_n364), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(KEYINPUT61), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n888), .A2(new_n364), .A3(new_n678), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n905));
  OAI211_X1 g704(.A(KEYINPUT125), .B(new_n905), .C1(new_n900), .C2(new_n364), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(G1351gat));
  NAND2_X1  g706(.A1(new_n644), .A2(new_n883), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n849), .A2(new_n830), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(G197gat), .B1(new_n910), .B2(new_n326), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n798), .A2(new_n668), .A3(new_n908), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n326), .A2(G197gat), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(G1352gat));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT126), .ZN(new_n917));
  NOR4_X1   g716(.A1(new_n798), .A2(G204gat), .A3(new_n668), .A4(new_n908), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(new_n360), .ZN(new_n919));
  INV_X1    g718(.A(G204gat), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n882), .A2(new_n920), .A3(new_n636), .A4(new_n909), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n921), .A2(KEYINPUT126), .A3(new_n708), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n916), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(G204gat), .B1(new_n850), .B2(new_n908), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n918), .A2(new_n917), .A3(new_n360), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT126), .B1(new_n921), .B2(new_n708), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n926), .A3(KEYINPUT62), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n923), .A2(new_n924), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT127), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n923), .A2(new_n930), .A3(new_n924), .A4(new_n927), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1353gat));
  OR3_X1    g731(.A1(new_n913), .A2(G211gat), .A3(new_n797), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n910), .A2(new_n797), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n934), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT63), .B1(new_n934), .B2(G211gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(G1354gat));
  OAI21_X1  g736(.A(G218gat), .B1(new_n910), .B2(new_n296), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n296), .A2(G218gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n913), .B2(new_n939), .ZN(G1355gat));
endmodule


