//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n553, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n573, new_n574, new_n575,
    new_n576, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT67), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  NAND3_X1  g033(.A1(new_n458), .A2(G101), .A3(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(G125), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n459), .B1(new_n463), .B2(new_n458), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n466), .A2(new_n468), .A3(G137), .A4(new_n458), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT68), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n462), .A2(new_n471), .A3(G137), .A4(new_n458), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n464), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n474), .B(new_n475), .ZN(G160));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n458), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n466), .A2(new_n468), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(new_n458), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n479), .A2(G2105), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n483), .A2(KEYINPUT70), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n483), .A2(KEYINPUT70), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n478), .B(new_n481), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND2_X1  g062(.A1(G102), .A2(G2104), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .A3(G138), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n488), .B1(new_n479), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(new_n458), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n466), .A2(new_n468), .A3(G126), .ZN(new_n493));
  NAND2_X1  g068(.A1(G114), .A2(G2104), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n462), .A2(G138), .A3(new_n458), .ZN(new_n497));
  XNOR2_X1  g072(.A(KEYINPUT71), .B(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n492), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(KEYINPUT72), .A2(KEYINPUT6), .A3(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n507), .A2(G50), .ZN(new_n508));
  AND2_X1   g083(.A1(G75), .A2(G651), .ZN(new_n509));
  OAI21_X1  g084(.A(G543), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G543), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n507), .A2(G88), .ZN(new_n516));
  AND2_X1   g091(.A1(G62), .A2(G651), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n510), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT73), .ZN(new_n522));
  XOR2_X1   g097(.A(new_n522), .B(KEYINPUT7), .Z(new_n523));
  AOI22_X1  g098(.A1(new_n507), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n512), .A2(new_n514), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n507), .A2(G543), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n524), .A2(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n523), .A2(new_n528), .ZN(G168));
  INV_X1    g104(.A(new_n527), .ZN(new_n530));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G64), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n525), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n530), .A2(G52), .B1(G651), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n507), .A2(new_n515), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G90), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n534), .A2(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  NAND2_X1  g114(.A1(new_n536), .A2(G81), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n530), .A2(G43), .ZN(new_n541));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n525), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G651), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n540), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT74), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n530), .A2(G43), .B1(G651), .B2(new_n544), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT74), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n548), .A2(new_n549), .A3(new_n540), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n553), .A2(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n525), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G651), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n560), .A2(KEYINPUT75), .A3(G651), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n536), .A2(G91), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT9), .B1(new_n527), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n507), .A2(new_n569), .A3(G53), .A4(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n565), .A2(new_n566), .A3(new_n571), .ZN(G299));
  OAI21_X1  g147(.A(KEYINPUT76), .B1(new_n523), .B2(new_n528), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NOR3_X1   g149(.A1(new_n523), .A2(new_n528), .A3(KEYINPUT76), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G286));
  AOI22_X1  g152(.A1(G87), .A2(new_n536), .B1(new_n530), .B2(G49), .ZN(new_n578));
  INV_X1    g153(.A(G74), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n504), .B1(new_n525), .B2(new_n579), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT77), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n578), .A2(new_n581), .ZN(G288));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  INV_X1    g158(.A(G48), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n583), .A2(new_n535), .B1(new_n527), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n515), .A2(G61), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT78), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n504), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n585), .A2(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(new_n536), .A2(G85), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n530), .A2(G47), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n591), .B(new_n592), .C1(new_n504), .C2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n535), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n507), .A2(new_n515), .A3(KEYINPUT10), .A4(G92), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n530), .A2(G54), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n525), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G651), .ZN(new_n605));
  AND3_X1   g180(.A1(new_n600), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n595), .B1(new_n606), .B2(G868), .ZN(G284));
  XNOR2_X1  g182(.A(G284), .B(KEYINPUT79), .ZN(G321));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(G299), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n576), .B2(new_n609), .ZN(G297));
  OAI21_X1  g186(.A(new_n610), .B1(new_n576), .B2(new_n609), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n606), .A2(new_n613), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n616), .A2(new_n609), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n551), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(KEYINPUT80), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(KEYINPUT80), .B2(new_n617), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n480), .A2(G123), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT82), .Z(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n626), .B(new_n627), .C1(G111), .C2(new_n458), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n482), .A2(G135), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n623), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(G2096), .Z(new_n631));
  NAND2_X1  g206(.A1(new_n458), .A2(G2104), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n479), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT13), .B(G2100), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n631), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XOR2_X1   g215(.A(KEYINPUT15), .B(G2435), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G1341), .B(G1348), .Z(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2443), .B(G2446), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT85), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n648), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n645), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(G14), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n655));
  XOR2_X1   g230(.A(G2067), .B(G2678), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  OAI21_X1  g233(.A(KEYINPUT17), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n658), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n660), .A2(new_n656), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n655), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2072), .B(G2078), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n662), .B(new_n663), .C1(new_n661), .C2(new_n655), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n663), .B2(new_n662), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2096), .B(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n670), .A2(KEYINPUT87), .ZN(new_n671));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(KEYINPUT87), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n671), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT20), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n668), .A2(new_n669), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  OR3_X1    g254(.A1(new_n673), .A2(new_n670), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n676), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n673), .A2(new_n679), .ZN(new_n682));
  NAND4_X1  g257(.A1(new_n677), .A2(new_n680), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT89), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1996), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT88), .B(G1986), .Z(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1991), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n685), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(G229));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n693), .A2(G33), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT25), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n482), .A2(G139), .ZN(new_n697));
  AOI22_X1  g272(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n696), .B(new_n697), .C1(new_n458), .C2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT94), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT95), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n694), .B1(new_n702), .B2(G29), .ZN(new_n703));
  INV_X1    g278(.A(G2072), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  NAND2_X1  g281(.A1(G168), .A2(G16), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G16), .B2(G21), .ZN(new_n708));
  INV_X1    g283(.A(G1966), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT100), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n705), .A2(new_n706), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(G160), .A2(G29), .ZN(new_n713));
  INV_X1    g288(.A(G34), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(KEYINPUT24), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(KEYINPUT24), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n715), .A2(new_n716), .A3(new_n693), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT96), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G2084), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT31), .B(G11), .ZN(new_n723));
  INV_X1    g298(.A(G28), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(KEYINPUT30), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(KEYINPUT30), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n725), .A2(new_n726), .A3(new_n693), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n723), .B(new_n727), .C1(new_n630), .C2(new_n693), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(KEYINPUT101), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(KEYINPUT101), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n729), .A2(new_n730), .B1(new_n709), .B2(new_n708), .ZN(new_n731));
  NOR2_X1   g306(.A1(G164), .A2(new_n693), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G27), .B2(new_n693), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(G2078), .Z(new_n734));
  INV_X1    g309(.A(G16), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G5), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G171), .B2(new_n735), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1961), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n722), .A2(new_n731), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n712), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n693), .A2(G32), .ZN(new_n742));
  AOI22_X1  g317(.A1(G129), .A2(new_n480), .B1(new_n482), .B2(G141), .ZN(new_n743));
  NAND3_X1  g318(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT26), .Z(new_n745));
  INV_X1    g320(.A(G105), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n743), .B(new_n745), .C1(new_n746), .C2(new_n632), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n747), .A2(KEYINPUT98), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(KEYINPUT98), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n742), .B1(new_n751), .B2(new_n693), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT27), .B(G1996), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT99), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n752), .B(new_n754), .ZN(new_n755));
  OR3_X1    g330(.A1(new_n720), .A2(KEYINPUT97), .A3(new_n721), .ZN(new_n756));
  OAI21_X1  g331(.A(KEYINPUT97), .B1(new_n720), .B2(new_n721), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n741), .A2(KEYINPUT102), .A3(new_n755), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT90), .B(G16), .ZN(new_n760));
  INV_X1    g335(.A(G19), .ZN(new_n761));
  OAI21_X1  g336(.A(KEYINPUT93), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OR3_X1    g337(.A1(new_n760), .A2(KEYINPUT93), .A3(new_n761), .ZN(new_n763));
  INV_X1    g338(.A(new_n760), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n762), .B(new_n763), .C1(new_n551), .C2(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1341), .ZN(new_n766));
  NAND2_X1  g341(.A1(G299), .A2(G16), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n764), .A2(KEYINPUT23), .A3(G20), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT23), .ZN(new_n769));
  INV_X1    g344(.A(G20), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n760), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n767), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1956), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n693), .A2(G26), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n480), .A2(G128), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n482), .A2(G140), .ZN(new_n776));
  NOR2_X1   g351(.A1(G104), .A2(G2105), .ZN(new_n777));
  OAI21_X1  g352(.A(G2104), .B1(new_n458), .B2(G116), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n775), .B(new_n776), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n774), .B1(new_n779), .B2(G29), .ZN(new_n780));
  MUX2_X1   g355(.A(new_n774), .B(new_n780), .S(KEYINPUT28), .Z(new_n781));
  INV_X1    g356(.A(G2067), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(KEYINPUT92), .B1(G4), .B2(G16), .ZN(new_n784));
  OR3_X1    g359(.A1(KEYINPUT92), .A2(G4), .A3(G16), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n598), .A2(new_n599), .B1(G651), .B2(new_n604), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(new_n601), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n784), .B(new_n785), .C1(new_n787), .C2(new_n735), .ZN(new_n788));
  INV_X1    g363(.A(G1348), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR4_X1   g365(.A1(new_n766), .A2(new_n773), .A3(new_n783), .A4(new_n790), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n759), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n735), .A2(G23), .ZN(new_n793));
  INV_X1    g368(.A(G288), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n735), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(KEYINPUT33), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(KEYINPUT33), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n796), .A2(G1976), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n764), .A2(G22), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G166), .B2(new_n764), .ZN(new_n800));
  INV_X1    g375(.A(G1971), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n735), .A2(G6), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n585), .A2(new_n589), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n735), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT32), .B(G1981), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n796), .A2(new_n797), .ZN(new_n809));
  INV_X1    g384(.A(G1976), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n803), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT34), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n764), .A2(G24), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G290), .B2(new_n760), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(G1986), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT34), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n803), .A2(new_n818), .A3(new_n808), .A4(new_n811), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n693), .A2(G25), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n480), .A2(G119), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n482), .A2(G131), .ZN(new_n822));
  OR2_X1    g397(.A1(G95), .A2(G2105), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n823), .B(G2104), .C1(G107), .C2(new_n458), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n820), .B1(new_n826), .B2(new_n693), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT35), .B(G1991), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G1986), .B2(new_n816), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n813), .A2(new_n817), .A3(new_n819), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n830), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n812), .B2(KEYINPUT34), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n836), .A2(new_n832), .A3(new_n817), .A4(new_n819), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n693), .A2(G35), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(G162), .B2(new_n693), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT29), .B(G2090), .Z(new_n841));
  XOR2_X1   g416(.A(new_n840), .B(new_n841), .Z(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n741), .A2(new_n755), .A3(new_n758), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT102), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n792), .A2(new_n838), .A3(new_n843), .A4(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(G311));
  NAND2_X1  g423(.A1(new_n847), .A2(KEYINPUT103), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n846), .A2(new_n759), .A3(new_n791), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT103), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n850), .A2(new_n851), .A3(new_n843), .A4(new_n838), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n852), .ZN(G150));
  AOI22_X1  g428(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n854), .A2(new_n504), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n507), .A2(new_n515), .A3(G93), .ZN(new_n856));
  XOR2_X1   g431(.A(KEYINPUT105), .B(G55), .Z(new_n857));
  NOR2_X1   g432(.A1(new_n527), .A2(new_n857), .ZN(new_n858));
  NOR3_X1   g433(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(G860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT37), .Z(new_n862));
  AOI21_X1  g437(.A(new_n859), .B1(new_n547), .B2(new_n550), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n859), .A2(new_n546), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT106), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n866), .B(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n787), .A2(new_n613), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT39), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n869), .B(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n862), .B1(new_n872), .B2(G860), .ZN(G145));
  XNOR2_X1  g448(.A(new_n750), .B(new_n779), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n500), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n875), .A2(new_n701), .ZN(new_n876));
  INV_X1    g451(.A(new_n702), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n480), .A2(G130), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n482), .A2(G142), .ZN(new_n881));
  OR2_X1    g456(.A1(G106), .A2(G2105), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n882), .B(G2104), .C1(G118), .C2(new_n458), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n825), .B(new_n884), .Z(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n635), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n630), .ZN(new_n887));
  XNOR2_X1  g462(.A(G162), .B(G160), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n879), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n887), .B(new_n888), .Z(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(new_n876), .B2(new_n878), .ZN(new_n892));
  INV_X1    g467(.A(G37), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n890), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g470(.A(new_n616), .B1(new_n863), .B2(new_n865), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n551), .A2(new_n860), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(new_n615), .A3(new_n864), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  AOI22_X1  g474(.A1(new_n563), .A2(new_n564), .B1(G91), .B2(new_n536), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n606), .A2(new_n900), .A3(new_n571), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n787), .A2(G299), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT107), .B1(new_n903), .B2(KEYINPUT41), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n787), .A2(G299), .ZN(new_n906));
  AOI22_X1  g481(.A1(new_n900), .A2(new_n571), .B1(new_n786), .B2(new_n601), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT41), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n901), .A2(new_n909), .A3(new_n902), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT107), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n899), .B1(new_n905), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT108), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n899), .A2(new_n903), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n899), .B(new_n915), .C1(new_n905), .C2(new_n911), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(G290), .B(KEYINPUT109), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(G288), .ZN(new_n921));
  XNOR2_X1  g496(.A(G303), .B(new_n805), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n922), .A2(KEYINPUT110), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n922), .A2(KEYINPUT110), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n921), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n913), .A2(KEYINPUT42), .A3(new_n914), .A4(new_n916), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n919), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n927), .B1(new_n919), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g505(.A(G868), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT111), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n860), .A2(new_n609), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n931), .B2(new_n933), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(G295));
  NAND2_X1  g511(.A1(new_n931), .A2(new_n933), .ZN(G331));
  NAND2_X1  g512(.A1(new_n908), .A2(new_n910), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n904), .ZN(new_n941));
  INV_X1    g516(.A(new_n575), .ZN(new_n942));
  AOI21_X1  g517(.A(G301), .B1(new_n942), .B2(new_n573), .ZN(new_n943));
  NAND2_X1  g518(.A1(G168), .A2(G301), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n866), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(G171), .B1(new_n574), .B2(new_n575), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n947), .B(new_n944), .C1(new_n865), .C2(new_n863), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n941), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT112), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n949), .A2(new_n903), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n924), .A2(new_n926), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n941), .A2(new_n949), .A3(KEYINPUT112), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n952), .A2(new_n954), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n949), .A2(new_n938), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n927), .B1(new_n953), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n957), .A2(new_n959), .A3(new_n960), .A4(new_n893), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n961), .A2(KEYINPUT113), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n952), .A2(new_n954), .A3(new_n956), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n927), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n957), .A2(new_n893), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT43), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n961), .A2(KEYINPUT113), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n962), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n966), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n972), .A2(KEYINPUT43), .A3(new_n959), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT43), .B1(new_n972), .B2(new_n964), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT44), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n971), .A2(new_n975), .ZN(G397));
  INV_X1    g551(.A(new_n459), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n460), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n977), .B1(new_n979), .B2(G2105), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n980), .A2(G40), .A3(new_n470), .A4(new_n472), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n473), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n984), .A2(KEYINPUT114), .A3(new_n980), .A4(G40), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1384), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT45), .B1(new_n500), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n825), .A2(new_n828), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n779), .B(new_n782), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n751), .A2(G1996), .ZN(new_n995));
  INV_X1    g570(.A(G1996), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n750), .A2(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n993), .B(new_n994), .C1(new_n995), .C2(new_n997), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n779), .A2(G2067), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n992), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n992), .B1(new_n751), .B2(new_n994), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n991), .A2(KEYINPUT46), .A3(new_n996), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT46), .B1(new_n991), .B2(new_n996), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1004), .B(KEYINPUT47), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n994), .B1(new_n995), .B2(new_n997), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n825), .A2(new_n828), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1006), .A2(new_n1007), .A3(new_n993), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n991), .ZN(new_n1010));
  NOR2_X1   g585(.A1(G290), .A2(G1986), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n991), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1012), .B(KEYINPUT48), .ZN(new_n1013));
  AOI211_X1 g588(.A(new_n1000), .B(new_n1005), .C1(new_n1010), .C2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G8), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n500), .A2(new_n988), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT50), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n500), .A2(new_n1018), .A3(new_n988), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n986), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n1020), .A2(G2090), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n988), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n986), .A2(new_n990), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n801), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1015), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G303), .A2(G8), .ZN(new_n1026));
  XOR2_X1   g601(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n1027));
  XNOR2_X1  g602(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1025), .B(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(G305), .A2(G1981), .ZN(new_n1030));
  OR3_X1    g605(.A1(new_n585), .A2(G1981), .A3(new_n589), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(KEYINPUT49), .A3(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1032), .B(KEYINPUT116), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1016), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT114), .B1(new_n474), .B2(G40), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n981), .A2(new_n982), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(new_n1015), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1033), .B(new_n1039), .C1(KEYINPUT49), .C2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1037), .B(G8), .C1(new_n810), .C2(G288), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT52), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n794), .A2(G1976), .ZN(new_n1044));
  OR3_X1    g619(.A1(new_n1042), .A2(KEYINPUT52), .A3(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1041), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1029), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1023), .A2(new_n709), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n986), .A2(new_n721), .A3(new_n1017), .A4(new_n1019), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1015), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1047), .A2(new_n576), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(KEYINPUT63), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1046), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(new_n1025), .A3(new_n1028), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1047), .A2(new_n576), .A3(new_n1050), .A4(new_n1053), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1041), .A2(new_n810), .A3(new_n794), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n1031), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n1039), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1055), .A2(new_n1057), .A3(new_n1058), .A4(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1038), .A2(new_n782), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1020), .A2(new_n789), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1063), .A2(new_n787), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n787), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT60), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT61), .ZN(new_n1068));
  INV_X1    g643(.A(G1956), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1020), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n1071));
  XNOR2_X1  g646(.A(G299), .B(new_n1071), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n988), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(new_n989), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT56), .B(G2072), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(new_n986), .A3(new_n1075), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1070), .A2(new_n1072), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1072), .B1(new_n1070), .B2(new_n1076), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1068), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1070), .A2(new_n1076), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1072), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1070), .A2(new_n1072), .A3(new_n1076), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(KEYINPUT61), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT60), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1063), .A2(new_n1085), .A3(new_n606), .A4(new_n1064), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1079), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT118), .B(G1996), .ZN(new_n1090));
  AND4_X1   g665(.A1(new_n986), .A2(new_n990), .A3(new_n1022), .A4(new_n1090), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT58), .B(G1341), .Z(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1093), .B1(new_n986), .B2(new_n1034), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1089), .B(new_n551), .C1(new_n1091), .C2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT119), .ZN(new_n1096));
  INV_X1    g671(.A(new_n551), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1037), .A2(new_n1092), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1074), .A2(new_n986), .A3(new_n1090), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1096), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT59), .B1(new_n1100), .B2(new_n1089), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1088), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1095), .A2(KEYINPUT119), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1107), .A2(KEYINPUT121), .A3(new_n1104), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1067), .B(new_n1087), .C1(new_n1106), .C2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1078), .B1(new_n1066), .B2(new_n1083), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n981), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(G2078), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n990), .A2(new_n1112), .A3(new_n1022), .A4(new_n1114), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1115), .A2(KEYINPUT125), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1113), .B1(new_n1023), .B2(G2078), .ZN(new_n1117));
  INV_X1    g692(.A(G1961), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1020), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1115), .A2(KEYINPUT125), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1116), .A2(new_n1117), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT126), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1121), .B(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1123), .A2(G301), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1117), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1114), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1119), .B1(new_n1023), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT124), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1119), .B(new_n1129), .C1(new_n1023), .C2(new_n1126), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1125), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT54), .B1(new_n1131), .B2(G171), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1131), .A2(G301), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n1121), .B2(G171), .ZN(new_n1135));
  OAI22_X1  g710(.A1(new_n1124), .A2(new_n1132), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1049), .ZN(new_n1139));
  AOI21_X1  g714(.A(G1966), .B1(new_n1074), .B2(new_n986), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1048), .A2(KEYINPUT122), .A3(new_n1049), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1141), .A2(G168), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT51), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1144), .A2(new_n1015), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1137), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1143), .A2(new_n1137), .A3(new_n1145), .ZN(new_n1148));
  NOR2_X1   g723(.A1(G168), .A2(new_n1015), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1050), .A2(KEYINPUT51), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1147), .A2(new_n1148), .A3(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1149), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1111), .A2(new_n1136), .A3(new_n1157), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1143), .A2(new_n1137), .A3(new_n1145), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1159), .A2(new_n1146), .A3(new_n1150), .ZN(new_n1160));
  OAI21_X1  g735(.A(KEYINPUT62), .B1(new_n1160), .B2(new_n1155), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1152), .A2(new_n1162), .A3(new_n1156), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1161), .A2(new_n1133), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1158), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1062), .B1(new_n1165), .B2(new_n1047), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1009), .B1(G1986), .B2(G290), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1011), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n992), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1014), .B1(new_n1166), .B2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g745(.A1(new_n894), .A2(new_n653), .ZN(new_n1172));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n1173));
  INV_X1    g747(.A(G319), .ZN(new_n1174));
  OR2_X1    g748(.A1(G227), .A2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g749(.A(new_n691), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g750(.A(new_n1176), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1177));
  AND3_X1   g751(.A1(new_n969), .A2(new_n1172), .A3(new_n1177), .ZN(G308));
  NAND3_X1  g752(.A1(new_n969), .A2(new_n1172), .A3(new_n1177), .ZN(G225));
endmodule


