

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U556 ( .A1(G2104), .A2(n541), .ZN(n883) );
  AND2_X2 U557 ( .A1(n541), .A2(G2104), .ZN(n886) );
  AND2_X1 U558 ( .A1(G160), .A2(G40), .ZN(n609) );
  OR2_X1 U559 ( .A1(n645), .A2(n644), .ZN(n655) );
  NOR2_X1 U560 ( .A1(n695), .A2(KEYINPUT33), .ZN(n696) );
  OR2_X1 U561 ( .A1(n712), .A2(n711), .ZN(n523) );
  INV_X1 U562 ( .A(KEYINPUT30), .ZN(n666) );
  XNOR2_X1 U563 ( .A(n666), .B(KEYINPUT97), .ZN(n667) );
  XNOR2_X1 U564 ( .A(n668), .B(n667), .ZN(n669) );
  INV_X1 U565 ( .A(KEYINPUT29), .ZN(n656) );
  BUF_X1 U566 ( .A(n637), .Z(n664) );
  INV_X1 U567 ( .A(KEYINPUT99), .ZN(n678) );
  INV_X1 U568 ( .A(KEYINPUT17), .ZN(n535) );
  XNOR2_X1 U569 ( .A(n535), .B(KEYINPUT66), .ZN(n536) );
  INV_X1 U570 ( .A(G651), .ZN(n530) );
  XNOR2_X1 U571 ( .A(n537), .B(n536), .ZN(n716) );
  NOR2_X1 U572 ( .A1(G651), .A2(n592), .ZN(n795) );
  NAND2_X1 U573 ( .A1(n623), .A2(n622), .ZN(n984) );
  XOR2_X1 U574 ( .A(KEYINPUT0), .B(G543), .Z(n592) );
  NAND2_X1 U575 ( .A1(n795), .A2(G47), .ZN(n527) );
  NOR2_X1 U576 ( .A1(G543), .A2(n530), .ZN(n524) );
  XOR2_X1 U577 ( .A(KEYINPUT68), .B(n524), .Z(n525) );
  XNOR2_X2 U578 ( .A(KEYINPUT1), .B(n525), .ZN(n791) );
  NAND2_X1 U579 ( .A1(G60), .A2(n791), .ZN(n526) );
  NAND2_X1 U580 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U581 ( .A(KEYINPUT69), .B(n528), .ZN(n534) );
  NOR2_X1 U582 ( .A1(G543), .A2(G651), .ZN(n529) );
  XNOR2_X1 U583 ( .A(n529), .B(KEYINPUT64), .ZN(n792) );
  NAND2_X1 U584 ( .A1(n792), .A2(G85), .ZN(n532) );
  NOR2_X1 U585 ( .A1(n592), .A2(n530), .ZN(n796) );
  NAND2_X1 U586 ( .A1(n796), .A2(G72), .ZN(n531) );
  AND2_X1 U587 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U588 ( .A1(n534), .A2(n533), .ZN(G290) );
  NOR2_X1 U589 ( .A1(G2105), .A2(G2104), .ZN(n537) );
  NAND2_X1 U590 ( .A1(n716), .A2(G138), .ZN(n538) );
  XNOR2_X1 U591 ( .A(n538), .B(KEYINPUT88), .ZN(n540) );
  AND2_X1 U592 ( .A1(G2105), .A2(G2104), .ZN(n882) );
  NAND2_X1 U593 ( .A1(n882), .A2(G114), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n540), .A2(n539), .ZN(n545) );
  INV_X1 U595 ( .A(G2105), .ZN(n541) );
  NAND2_X1 U596 ( .A1(G102), .A2(n886), .ZN(n543) );
  NAND2_X1 U597 ( .A1(G126), .A2(n883), .ZN(n542) );
  NAND2_X1 U598 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U599 ( .A1(n545), .A2(n544), .ZN(G164) );
  NAND2_X1 U600 ( .A1(n716), .A2(G137), .ZN(n546) );
  XOR2_X1 U601 ( .A(KEYINPUT67), .B(n546), .Z(n550) );
  NAND2_X1 U602 ( .A1(G101), .A2(n886), .ZN(n547) );
  XNOR2_X1 U603 ( .A(n547), .B(KEYINPUT65), .ZN(n548) );
  XNOR2_X1 U604 ( .A(n548), .B(KEYINPUT23), .ZN(n549) );
  NAND2_X1 U605 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U606 ( .A1(G113), .A2(n882), .ZN(n552) );
  NAND2_X1 U607 ( .A1(G125), .A2(n883), .ZN(n551) );
  NAND2_X1 U608 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X4 U609 ( .A1(n554), .A2(n553), .ZN(G160) );
  NAND2_X1 U610 ( .A1(n795), .A2(G50), .ZN(n561) );
  NAND2_X1 U611 ( .A1(n796), .A2(G75), .ZN(n556) );
  NAND2_X1 U612 ( .A1(G88), .A2(n792), .ZN(n555) );
  NAND2_X1 U613 ( .A1(n556), .A2(n555), .ZN(n559) );
  NAND2_X1 U614 ( .A1(n791), .A2(G62), .ZN(n557) );
  XOR2_X1 U615 ( .A(KEYINPUT82), .B(n557), .Z(n558) );
  NOR2_X1 U616 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U618 ( .A(KEYINPUT83), .B(n562), .Z(G303) );
  NAND2_X1 U619 ( .A1(n795), .A2(G51), .ZN(n563) );
  XNOR2_X1 U620 ( .A(n563), .B(KEYINPUT76), .ZN(n565) );
  NAND2_X1 U621 ( .A1(G63), .A2(n791), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U623 ( .A(KEYINPUT6), .B(n566), .ZN(n573) );
  NAND2_X1 U624 ( .A1(G89), .A2(n792), .ZN(n567) );
  XNOR2_X1 U625 ( .A(n567), .B(KEYINPUT4), .ZN(n569) );
  NAND2_X1 U626 ( .A1(G76), .A2(n796), .ZN(n568) );
  NAND2_X1 U627 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U628 ( .A(KEYINPUT75), .B(n570), .ZN(n571) );
  XNOR2_X1 U629 ( .A(KEYINPUT5), .B(n571), .ZN(n572) );
  NOR2_X1 U630 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U631 ( .A(n574), .B(KEYINPUT7), .ZN(n575) );
  XNOR2_X1 U632 ( .A(n575), .B(KEYINPUT77), .ZN(G168) );
  XOR2_X1 U633 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U634 ( .A1(n791), .A2(G65), .ZN(n576) );
  XNOR2_X1 U635 ( .A(n576), .B(KEYINPUT72), .ZN(n583) );
  NAND2_X1 U636 ( .A1(G53), .A2(n795), .ZN(n578) );
  NAND2_X1 U637 ( .A1(G91), .A2(n792), .ZN(n577) );
  NAND2_X1 U638 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U639 ( .A1(G78), .A2(n796), .ZN(n579) );
  XNOR2_X1 U640 ( .A(KEYINPUT71), .B(n579), .ZN(n580) );
  NOR2_X1 U641 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U642 ( .A1(n583), .A2(n582), .ZN(G299) );
  NAND2_X1 U643 ( .A1(n796), .A2(G77), .ZN(n585) );
  NAND2_X1 U644 ( .A1(G90), .A2(n792), .ZN(n584) );
  NAND2_X1 U645 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U646 ( .A(n586), .B(KEYINPUT9), .ZN(n588) );
  NAND2_X1 U647 ( .A1(G64), .A2(n791), .ZN(n587) );
  NAND2_X1 U648 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U649 ( .A1(n795), .A2(G52), .ZN(n589) );
  XOR2_X1 U650 ( .A(KEYINPUT70), .B(n589), .Z(n590) );
  NOR2_X1 U651 ( .A1(n591), .A2(n590), .ZN(G171) );
  NAND2_X1 U652 ( .A1(n795), .A2(G49), .ZN(n597) );
  NAND2_X1 U653 ( .A1(G87), .A2(n592), .ZN(n594) );
  NAND2_X1 U654 ( .A1(G74), .A2(G651), .ZN(n593) );
  NAND2_X1 U655 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U656 ( .A1(n791), .A2(n595), .ZN(n596) );
  NAND2_X1 U657 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U658 ( .A(KEYINPUT81), .B(n598), .Z(G288) );
  NAND2_X1 U659 ( .A1(G61), .A2(n791), .ZN(n600) );
  NAND2_X1 U660 ( .A1(G86), .A2(n792), .ZN(n599) );
  NAND2_X1 U661 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U662 ( .A1(n796), .A2(G73), .ZN(n601) );
  XOR2_X1 U663 ( .A(KEYINPUT2), .B(n601), .Z(n602) );
  NOR2_X1 U664 ( .A1(n603), .A2(n602), .ZN(n605) );
  NAND2_X1 U665 ( .A1(n795), .A2(G48), .ZN(n604) );
  NAND2_X1 U666 ( .A1(n605), .A2(n604), .ZN(G305) );
  INV_X1 U667 ( .A(G303), .ZN(G166) );
  XOR2_X1 U668 ( .A(G1986), .B(KEYINPUT89), .Z(n606) );
  XNOR2_X1 U669 ( .A(G290), .B(n606), .ZN(n981) );
  NOR2_X1 U670 ( .A1(G164), .A2(G1384), .ZN(n608) );
  NAND2_X1 U671 ( .A1(G160), .A2(G40), .ZN(n607) );
  NOR2_X1 U672 ( .A1(n608), .A2(n607), .ZN(n761) );
  NAND2_X1 U673 ( .A1(n981), .A2(n761), .ZN(n748) );
  NAND2_X1 U674 ( .A1(n609), .A2(n608), .ZN(n637) );
  NAND2_X1 U675 ( .A1(G8), .A2(n637), .ZN(n704) );
  NOR2_X1 U676 ( .A1(G2090), .A2(n664), .ZN(n610) );
  XNOR2_X1 U677 ( .A(n610), .B(KEYINPUT98), .ZN(n612) );
  NOR2_X1 U678 ( .A1(n704), .A2(G1971), .ZN(n611) );
  NOR2_X1 U679 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U680 ( .A1(n613), .A2(G303), .ZN(n677) );
  NAND2_X1 U681 ( .A1(G56), .A2(n791), .ZN(n614) );
  XNOR2_X1 U682 ( .A(n614), .B(KEYINPUT14), .ZN(n620) );
  NAND2_X1 U683 ( .A1(G81), .A2(n792), .ZN(n615) );
  XNOR2_X1 U684 ( .A(n615), .B(KEYINPUT12), .ZN(n617) );
  NAND2_X1 U685 ( .A1(G68), .A2(n796), .ZN(n616) );
  NAND2_X1 U686 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U687 ( .A(KEYINPUT13), .B(n618), .ZN(n619) );
  NAND2_X1 U688 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U689 ( .A(n621), .B(KEYINPUT73), .ZN(n623) );
  NAND2_X1 U690 ( .A1(n795), .A2(G43), .ZN(n622) );
  INV_X1 U691 ( .A(n637), .ZN(n624) );
  NAND2_X1 U692 ( .A1(G1996), .A2(n624), .ZN(n625) );
  XOR2_X1 U693 ( .A(KEYINPUT26), .B(n625), .Z(n626) );
  NOR2_X1 U694 ( .A1(n984), .A2(n626), .ZN(n628) );
  NAND2_X1 U695 ( .A1(G1341), .A2(n664), .ZN(n627) );
  NAND2_X1 U696 ( .A1(n628), .A2(n627), .ZN(n647) );
  NAND2_X1 U697 ( .A1(G54), .A2(n795), .ZN(n630) );
  NAND2_X1 U698 ( .A1(G79), .A2(n796), .ZN(n629) );
  NAND2_X1 U699 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U700 ( .A1(G66), .A2(n791), .ZN(n632) );
  NAND2_X1 U701 ( .A1(G92), .A2(n792), .ZN(n631) );
  NAND2_X1 U702 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U703 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U704 ( .A(n635), .B(KEYINPUT15), .ZN(n974) );
  NOR2_X1 U705 ( .A1(n647), .A2(n974), .ZN(n636) );
  XNOR2_X1 U706 ( .A(KEYINPUT96), .B(n636), .ZN(n645) );
  INV_X1 U707 ( .A(n637), .ZN(n659) );
  NOR2_X1 U708 ( .A1(n659), .A2(G1348), .ZN(n639) );
  NOR2_X1 U709 ( .A1(G2067), .A2(n664), .ZN(n638) );
  NOR2_X1 U710 ( .A1(n639), .A2(n638), .ZN(n643) );
  INV_X1 U711 ( .A(G299), .ZN(n973) );
  NAND2_X1 U712 ( .A1(n659), .A2(G2072), .ZN(n640) );
  XNOR2_X1 U713 ( .A(n640), .B(KEYINPUT27), .ZN(n642) );
  INV_X1 U714 ( .A(G1956), .ZN(n1004) );
  NOR2_X1 U715 ( .A1(n1004), .A2(n659), .ZN(n641) );
  NOR2_X1 U716 ( .A1(n642), .A2(n641), .ZN(n650) );
  NAND2_X1 U717 ( .A1(n973), .A2(n650), .ZN(n646) );
  NAND2_X1 U718 ( .A1(n643), .A2(n646), .ZN(n644) );
  INV_X1 U719 ( .A(n646), .ZN(n649) );
  NAND2_X1 U720 ( .A1(n647), .A2(n974), .ZN(n648) );
  OR2_X1 U721 ( .A1(n649), .A2(n648), .ZN(n653) );
  NOR2_X1 U722 ( .A1(n973), .A2(n650), .ZN(n651) );
  XOR2_X1 U723 ( .A(n651), .B(KEYINPUT28), .Z(n652) );
  AND2_X1 U724 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U725 ( .A1(n655), .A2(n654), .ZN(n657) );
  XNOR2_X1 U726 ( .A(n657), .B(n656), .ZN(n663) );
  NOR2_X1 U727 ( .A1(n659), .A2(G1961), .ZN(n658) );
  XNOR2_X1 U728 ( .A(n658), .B(KEYINPUT95), .ZN(n661) );
  XNOR2_X1 U729 ( .A(G2078), .B(KEYINPUT25), .ZN(n956) );
  NAND2_X1 U730 ( .A1(n659), .A2(n956), .ZN(n660) );
  NAND2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n670) );
  NAND2_X1 U732 ( .A1(n670), .A2(G171), .ZN(n662) );
  NAND2_X1 U733 ( .A1(n663), .A2(n662), .ZN(n675) );
  NOR2_X1 U734 ( .A1(G1966), .A2(n704), .ZN(n683) );
  NOR2_X1 U735 ( .A1(G2084), .A2(n664), .ZN(n684) );
  NOR2_X1 U736 ( .A1(n683), .A2(n684), .ZN(n665) );
  NAND2_X1 U737 ( .A1(G8), .A2(n665), .ZN(n668) );
  NOR2_X1 U738 ( .A1(G168), .A2(n669), .ZN(n672) );
  NOR2_X1 U739 ( .A1(G171), .A2(n670), .ZN(n671) );
  NOR2_X1 U740 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U741 ( .A(KEYINPUT31), .B(n673), .Z(n674) );
  NAND2_X1 U742 ( .A1(n675), .A2(n674), .ZN(n686) );
  NAND2_X1 U743 ( .A1(G286), .A2(n686), .ZN(n676) );
  NAND2_X1 U744 ( .A1(n677), .A2(n676), .ZN(n679) );
  XNOR2_X1 U745 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U746 ( .A1(n680), .A2(G8), .ZN(n682) );
  INV_X1 U747 ( .A(KEYINPUT32), .ZN(n681) );
  XNOR2_X1 U748 ( .A(n682), .B(n681), .ZN(n707) );
  NAND2_X1 U749 ( .A1(G8), .A2(n684), .ZN(n685) );
  NAND2_X1 U750 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U751 ( .A1(n683), .A2(n687), .ZN(n706) );
  NAND2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n991) );
  INV_X1 U753 ( .A(n991), .ZN(n691) );
  OR2_X1 U754 ( .A1(n706), .A2(n691), .ZN(n688) );
  NOR2_X1 U755 ( .A1(n707), .A2(n688), .ZN(n693) );
  NOR2_X1 U756 ( .A1(G1976), .A2(G288), .ZN(n697) );
  NOR2_X1 U757 ( .A1(G1971), .A2(G303), .ZN(n689) );
  NOR2_X1 U758 ( .A1(n697), .A2(n689), .ZN(n992) );
  XNOR2_X1 U759 ( .A(KEYINPUT100), .B(n992), .ZN(n690) );
  NOR2_X1 U760 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U762 ( .A1(n704), .A2(n694), .ZN(n695) );
  XNOR2_X1 U763 ( .A(n696), .B(KEYINPUT101), .ZN(n701) );
  XNOR2_X1 U764 ( .A(G1981), .B(G305), .ZN(n988) );
  NAND2_X1 U765 ( .A1(n697), .A2(KEYINPUT33), .ZN(n698) );
  NOR2_X1 U766 ( .A1(n704), .A2(n698), .ZN(n699) );
  NOR2_X1 U767 ( .A1(n988), .A2(n699), .ZN(n700) );
  AND2_X1 U768 ( .A1(n701), .A2(n700), .ZN(n715) );
  NOR2_X1 U769 ( .A1(G1981), .A2(G305), .ZN(n702) );
  XNOR2_X1 U770 ( .A(n702), .B(KEYINPUT24), .ZN(n703) );
  XNOR2_X1 U771 ( .A(n703), .B(KEYINPUT94), .ZN(n705) );
  INV_X1 U772 ( .A(n704), .ZN(n711) );
  NAND2_X1 U773 ( .A1(n705), .A2(n711), .ZN(n713) );
  NOR2_X1 U774 ( .A1(n707), .A2(n706), .ZN(n710) );
  NAND2_X1 U775 ( .A1(G166), .A2(G8), .ZN(n708) );
  NOR2_X1 U776 ( .A1(G2090), .A2(n708), .ZN(n709) );
  NOR2_X1 U777 ( .A1(n710), .A2(n709), .ZN(n712) );
  NAND2_X1 U778 ( .A1(n713), .A2(n523), .ZN(n714) );
  NOR2_X1 U779 ( .A1(n715), .A2(n714), .ZN(n746) );
  NAND2_X1 U780 ( .A1(n886), .A2(G104), .ZN(n718) );
  BUF_X1 U781 ( .A(n716), .Z(n887) );
  NAND2_X1 U782 ( .A1(G140), .A2(n887), .ZN(n717) );
  NAND2_X1 U783 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U784 ( .A(KEYINPUT34), .B(n719), .ZN(n725) );
  NAND2_X1 U785 ( .A1(G116), .A2(n882), .ZN(n721) );
  NAND2_X1 U786 ( .A1(G128), .A2(n883), .ZN(n720) );
  NAND2_X1 U787 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U788 ( .A(KEYINPUT90), .B(n722), .Z(n723) );
  XNOR2_X1 U789 ( .A(KEYINPUT35), .B(n723), .ZN(n724) );
  NOR2_X1 U790 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U791 ( .A(KEYINPUT36), .B(n726), .ZN(n896) );
  XNOR2_X1 U792 ( .A(KEYINPUT37), .B(G2067), .ZN(n759) );
  NOR2_X1 U793 ( .A1(n896), .A2(n759), .ZN(n925) );
  NAND2_X1 U794 ( .A1(n761), .A2(n925), .ZN(n756) );
  NAND2_X1 U795 ( .A1(n887), .A2(G141), .ZN(n727) );
  XNOR2_X1 U796 ( .A(n727), .B(KEYINPUT92), .ZN(n734) );
  NAND2_X1 U797 ( .A1(G117), .A2(n882), .ZN(n729) );
  NAND2_X1 U798 ( .A1(G129), .A2(n883), .ZN(n728) );
  NAND2_X1 U799 ( .A1(n729), .A2(n728), .ZN(n732) );
  NAND2_X1 U800 ( .A1(n886), .A2(G105), .ZN(n730) );
  XOR2_X1 U801 ( .A(KEYINPUT38), .B(n730), .Z(n731) );
  NOR2_X1 U802 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U803 ( .A1(n734), .A2(n733), .ZN(n875) );
  NAND2_X1 U804 ( .A1(G1996), .A2(n875), .ZN(n735) );
  XNOR2_X1 U805 ( .A(n735), .B(KEYINPUT93), .ZN(n744) );
  INV_X1 U806 ( .A(G1991), .ZN(n953) );
  NAND2_X1 U807 ( .A1(G107), .A2(n882), .ZN(n737) );
  NAND2_X1 U808 ( .A1(G119), .A2(n883), .ZN(n736) );
  NAND2_X1 U809 ( .A1(n737), .A2(n736), .ZN(n742) );
  NAND2_X1 U810 ( .A1(n886), .A2(G95), .ZN(n739) );
  NAND2_X1 U811 ( .A1(G131), .A2(n887), .ZN(n738) );
  NAND2_X1 U812 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U813 ( .A(KEYINPUT91), .B(n740), .Z(n741) );
  NOR2_X1 U814 ( .A1(n742), .A2(n741), .ZN(n893) );
  NOR2_X1 U815 ( .A1(n953), .A2(n893), .ZN(n743) );
  OR2_X1 U816 ( .A1(n744), .A2(n743), .ZN(n924) );
  NAND2_X1 U817 ( .A1(n924), .A2(n761), .ZN(n749) );
  NAND2_X1 U818 ( .A1(n756), .A2(n749), .ZN(n745) );
  NOR2_X1 U819 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U820 ( .A1(n748), .A2(n747), .ZN(n764) );
  NOR2_X1 U821 ( .A1(G1996), .A2(n875), .ZN(n936) );
  INV_X1 U822 ( .A(n749), .ZN(n753) );
  AND2_X1 U823 ( .A1(n953), .A2(n893), .ZN(n930) );
  NOR2_X1 U824 ( .A1(G1986), .A2(G290), .ZN(n750) );
  NOR2_X1 U825 ( .A1(n930), .A2(n750), .ZN(n751) );
  XNOR2_X1 U826 ( .A(n751), .B(KEYINPUT102), .ZN(n752) );
  NOR2_X1 U827 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U828 ( .A1(n936), .A2(n754), .ZN(n755) );
  XNOR2_X1 U829 ( .A(KEYINPUT39), .B(n755), .ZN(n757) );
  NAND2_X1 U830 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U831 ( .A(KEYINPUT103), .B(n758), .Z(n760) );
  NAND2_X1 U832 ( .A1(n896), .A2(n759), .ZN(n922) );
  NAND2_X1 U833 ( .A1(n760), .A2(n922), .ZN(n762) );
  NAND2_X1 U834 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U835 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U836 ( .A(n765), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U837 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U838 ( .A(G57), .ZN(G237) );
  INV_X1 U839 ( .A(G132), .ZN(G219) );
  INV_X1 U840 ( .A(G82), .ZN(G220) );
  NAND2_X1 U841 ( .A1(G7), .A2(G661), .ZN(n766) );
  XNOR2_X1 U842 ( .A(n766), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U843 ( .A(G223), .ZN(n831) );
  NAND2_X1 U844 ( .A1(n831), .A2(G567), .ZN(n767) );
  XOR2_X1 U845 ( .A(KEYINPUT11), .B(n767), .Z(G234) );
  INV_X1 U846 ( .A(G860), .ZN(n772) );
  OR2_X1 U847 ( .A1(n984), .A2(n772), .ZN(G153) );
  XOR2_X1 U848 ( .A(G171), .B(KEYINPUT74), .Z(G301) );
  NAND2_X1 U849 ( .A1(G868), .A2(G301), .ZN(n769) );
  INV_X1 U850 ( .A(G868), .ZN(n811) );
  NAND2_X1 U851 ( .A1(n974), .A2(n811), .ZN(n768) );
  NAND2_X1 U852 ( .A1(n769), .A2(n768), .ZN(G284) );
  NOR2_X1 U853 ( .A1(G286), .A2(n811), .ZN(n771) );
  NOR2_X1 U854 ( .A1(G868), .A2(G299), .ZN(n770) );
  NOR2_X1 U855 ( .A1(n771), .A2(n770), .ZN(G297) );
  NAND2_X1 U856 ( .A1(n772), .A2(G559), .ZN(n773) );
  INV_X1 U857 ( .A(n974), .ZN(n789) );
  NAND2_X1 U858 ( .A1(n773), .A2(n789), .ZN(n774) );
  XNOR2_X1 U859 ( .A(n774), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U860 ( .A1(G868), .A2(n984), .ZN(n777) );
  NAND2_X1 U861 ( .A1(G868), .A2(n789), .ZN(n775) );
  NOR2_X1 U862 ( .A1(G559), .A2(n775), .ZN(n776) );
  NOR2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U864 ( .A(KEYINPUT78), .B(n778), .ZN(G282) );
  NAND2_X1 U865 ( .A1(G123), .A2(n883), .ZN(n779) );
  XOR2_X1 U866 ( .A(KEYINPUT18), .B(n779), .Z(n780) );
  XNOR2_X1 U867 ( .A(n780), .B(KEYINPUT79), .ZN(n782) );
  NAND2_X1 U868 ( .A1(G111), .A2(n882), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n786) );
  NAND2_X1 U870 ( .A1(n886), .A2(G99), .ZN(n784) );
  NAND2_X1 U871 ( .A1(G135), .A2(n887), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U873 ( .A1(n786), .A2(n785), .ZN(n931) );
  XNOR2_X1 U874 ( .A(G2096), .B(n931), .ZN(n788) );
  INV_X1 U875 ( .A(G2100), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n788), .A2(n787), .ZN(G156) );
  NAND2_X1 U877 ( .A1(n789), .A2(G559), .ZN(n809) );
  XNOR2_X1 U878 ( .A(n984), .B(n809), .ZN(n790) );
  NOR2_X1 U879 ( .A1(G860), .A2(n790), .ZN(n802) );
  NAND2_X1 U880 ( .A1(G67), .A2(n791), .ZN(n794) );
  NAND2_X1 U881 ( .A1(G93), .A2(n792), .ZN(n793) );
  NAND2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n800) );
  NAND2_X1 U883 ( .A1(G55), .A2(n795), .ZN(n798) );
  NAND2_X1 U884 ( .A1(G80), .A2(n796), .ZN(n797) );
  NAND2_X1 U885 ( .A1(n798), .A2(n797), .ZN(n799) );
  OR2_X1 U886 ( .A1(n800), .A2(n799), .ZN(n812) );
  XOR2_X1 U887 ( .A(n812), .B(KEYINPUT80), .Z(n801) );
  XNOR2_X1 U888 ( .A(n802), .B(n801), .ZN(G145) );
  XNOR2_X1 U889 ( .A(G305), .B(G288), .ZN(n807) );
  XNOR2_X1 U890 ( .A(n973), .B(KEYINPUT19), .ZN(n803) );
  XOR2_X1 U891 ( .A(n803), .B(n812), .Z(n804) );
  XNOR2_X1 U892 ( .A(G166), .B(n804), .ZN(n805) );
  XNOR2_X1 U893 ( .A(n805), .B(G290), .ZN(n806) );
  XNOR2_X1 U894 ( .A(n807), .B(n806), .ZN(n808) );
  XNOR2_X1 U895 ( .A(n984), .B(n808), .ZN(n900) );
  XNOR2_X1 U896 ( .A(n809), .B(n900), .ZN(n810) );
  NAND2_X1 U897 ( .A1(n810), .A2(G868), .ZN(n814) );
  NAND2_X1 U898 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U899 ( .A1(n814), .A2(n813), .ZN(G295) );
  XOR2_X1 U900 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n816) );
  NAND2_X1 U901 ( .A1(G2084), .A2(G2078), .ZN(n815) );
  XNOR2_X1 U902 ( .A(n816), .B(n815), .ZN(n817) );
  NAND2_X1 U903 ( .A1(n817), .A2(G2090), .ZN(n818) );
  XOR2_X1 U904 ( .A(KEYINPUT85), .B(n818), .Z(n819) );
  XNOR2_X1 U905 ( .A(KEYINPUT21), .B(n819), .ZN(n820) );
  NAND2_X1 U906 ( .A1(n820), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U907 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U908 ( .A1(G220), .A2(G219), .ZN(n821) );
  XOR2_X1 U909 ( .A(KEYINPUT22), .B(n821), .Z(n822) );
  NOR2_X1 U910 ( .A1(G218), .A2(n822), .ZN(n823) );
  NAND2_X1 U911 ( .A1(G96), .A2(n823), .ZN(n919) );
  NAND2_X1 U912 ( .A1(n919), .A2(G2106), .ZN(n827) );
  NAND2_X1 U913 ( .A1(G69), .A2(G120), .ZN(n824) );
  NOR2_X1 U914 ( .A1(G237), .A2(n824), .ZN(n825) );
  NAND2_X1 U915 ( .A1(G108), .A2(n825), .ZN(n920) );
  NAND2_X1 U916 ( .A1(n920), .A2(G567), .ZN(n826) );
  NAND2_X1 U917 ( .A1(n827), .A2(n826), .ZN(n837) );
  NAND2_X1 U918 ( .A1(G661), .A2(G483), .ZN(n828) );
  XNOR2_X1 U919 ( .A(KEYINPUT86), .B(n828), .ZN(n829) );
  NOR2_X1 U920 ( .A1(n837), .A2(n829), .ZN(n836) );
  NAND2_X1 U921 ( .A1(n836), .A2(G36), .ZN(n830) );
  XOR2_X1 U922 ( .A(KEYINPUT87), .B(n830), .Z(G176) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n831), .ZN(G217) );
  NAND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n832) );
  XNOR2_X1 U925 ( .A(KEYINPUT105), .B(n832), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n833), .A2(G661), .ZN(n834) );
  XNOR2_X1 U927 ( .A(KEYINPUT106), .B(n834), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U929 ( .A1(n836), .A2(n835), .ZN(G188) );
  INV_X1 U930 ( .A(n837), .ZN(G319) );
  XOR2_X1 U931 ( .A(KEYINPUT107), .B(G2090), .Z(n839) );
  XNOR2_X1 U932 ( .A(G2078), .B(G2072), .ZN(n838) );
  XNOR2_X1 U933 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U934 ( .A(n840), .B(G2096), .Z(n842) );
  XNOR2_X1 U935 ( .A(G2067), .B(G2084), .ZN(n841) );
  XNOR2_X1 U936 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U937 ( .A(G2678), .B(KEYINPUT43), .Z(n844) );
  XNOR2_X1 U938 ( .A(KEYINPUT42), .B(G2100), .ZN(n843) );
  XNOR2_X1 U939 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U940 ( .A(n846), .B(n845), .Z(G227) );
  XOR2_X1 U941 ( .A(KEYINPUT109), .B(G1971), .Z(n848) );
  XNOR2_X1 U942 ( .A(G1961), .B(G1956), .ZN(n847) );
  XNOR2_X1 U943 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U944 ( .A(n849), .B(KEYINPUT41), .Z(n851) );
  XNOR2_X1 U945 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U946 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U947 ( .A(G1976), .B(G1981), .Z(n853) );
  XNOR2_X1 U948 ( .A(G1986), .B(G1966), .ZN(n852) );
  XNOR2_X1 U949 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U950 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U951 ( .A(KEYINPUT108), .B(G2474), .ZN(n856) );
  XNOR2_X1 U952 ( .A(n857), .B(n856), .ZN(G229) );
  NAND2_X1 U953 ( .A1(n886), .A2(G100), .ZN(n864) );
  NAND2_X1 U954 ( .A1(n882), .A2(G112), .ZN(n859) );
  NAND2_X1 U955 ( .A1(G136), .A2(n887), .ZN(n858) );
  NAND2_X1 U956 ( .A1(n859), .A2(n858), .ZN(n862) );
  NAND2_X1 U957 ( .A1(n883), .A2(G124), .ZN(n860) );
  XOR2_X1 U958 ( .A(KEYINPUT44), .B(n860), .Z(n861) );
  NOR2_X1 U959 ( .A1(n862), .A2(n861), .ZN(n863) );
  NAND2_X1 U960 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U961 ( .A(KEYINPUT110), .B(n865), .Z(G162) );
  XOR2_X1 U962 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n867) );
  XNOR2_X1 U963 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n866) );
  XNOR2_X1 U964 ( .A(n867), .B(n866), .ZN(n879) );
  NAND2_X1 U965 ( .A1(n886), .A2(G103), .ZN(n869) );
  NAND2_X1 U966 ( .A1(G139), .A2(n887), .ZN(n868) );
  NAND2_X1 U967 ( .A1(n869), .A2(n868), .ZN(n874) );
  NAND2_X1 U968 ( .A1(G115), .A2(n882), .ZN(n871) );
  NAND2_X1 U969 ( .A1(G127), .A2(n883), .ZN(n870) );
  NAND2_X1 U970 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U971 ( .A(KEYINPUT47), .B(n872), .Z(n873) );
  NOR2_X1 U972 ( .A1(n874), .A2(n873), .ZN(n926) );
  XNOR2_X1 U973 ( .A(n875), .B(n926), .ZN(n877) );
  XNOR2_X1 U974 ( .A(G164), .B(G160), .ZN(n876) );
  XNOR2_X1 U975 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U976 ( .A(n879), .B(n878), .ZN(n881) );
  XNOR2_X1 U977 ( .A(G162), .B(n931), .ZN(n880) );
  XNOR2_X1 U978 ( .A(n881), .B(n880), .ZN(n898) );
  NAND2_X1 U979 ( .A1(G118), .A2(n882), .ZN(n885) );
  NAND2_X1 U980 ( .A1(G130), .A2(n883), .ZN(n884) );
  NAND2_X1 U981 ( .A1(n885), .A2(n884), .ZN(n892) );
  NAND2_X1 U982 ( .A1(n886), .A2(G106), .ZN(n889) );
  NAND2_X1 U983 ( .A1(G142), .A2(n887), .ZN(n888) );
  NAND2_X1 U984 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U985 ( .A(n890), .B(KEYINPUT45), .Z(n891) );
  NOR2_X1 U986 ( .A1(n892), .A2(n891), .ZN(n894) );
  XOR2_X1 U987 ( .A(n894), .B(n893), .Z(n895) );
  XNOR2_X1 U988 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U989 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U990 ( .A1(G37), .A2(n899), .ZN(G395) );
  XNOR2_X1 U991 ( .A(G286), .B(n974), .ZN(n901) );
  XNOR2_X1 U992 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U993 ( .A(n902), .B(G171), .ZN(n903) );
  NOR2_X1 U994 ( .A1(G37), .A2(n903), .ZN(G397) );
  XOR2_X1 U995 ( .A(G2443), .B(G2427), .Z(n905) );
  XNOR2_X1 U996 ( .A(G2438), .B(G2454), .ZN(n904) );
  XNOR2_X1 U997 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U998 ( .A(n906), .B(G2435), .Z(n908) );
  XNOR2_X1 U999 ( .A(G1341), .B(G1348), .ZN(n907) );
  XNOR2_X1 U1000 ( .A(n908), .B(n907), .ZN(n912) );
  XOR2_X1 U1001 ( .A(G2430), .B(G2446), .Z(n910) );
  XNOR2_X1 U1002 ( .A(KEYINPUT104), .B(G2451), .ZN(n909) );
  XNOR2_X1 U1003 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1004 ( .A(n912), .B(n911), .Z(n913) );
  NAND2_X1 U1005 ( .A1(G14), .A2(n913), .ZN(n921) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n921), .ZN(n916) );
  NOR2_X1 U1007 ( .A1(G227), .A2(G229), .ZN(n914) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1009 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1011 ( .A1(n918), .A2(n917), .ZN(G225) );
  XNOR2_X1 U1012 ( .A(KEYINPUT113), .B(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G120), .ZN(G236) );
  INV_X1 U1015 ( .A(G96), .ZN(G221) );
  INV_X1 U1016 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(G325) );
  INV_X1 U1018 ( .A(G325), .ZN(G261) );
  INV_X1 U1019 ( .A(G108), .ZN(G238) );
  INV_X1 U1020 ( .A(n921), .ZN(G401) );
  XNOR2_X1 U1021 ( .A(G2084), .B(G160), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n943) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n941) );
  XOR2_X1 U1024 ( .A(G2072), .B(n926), .Z(n928) );
  XOR2_X1 U1025 ( .A(G164), .B(G2078), .Z(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(n929), .B(KEYINPUT50), .ZN(n934) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(n932), .B(KEYINPUT114), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n939) );
  XOR2_X1 U1031 ( .A(G2090), .B(G162), .Z(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1033 ( .A(n937), .B(KEYINPUT51), .ZN(n938) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1036 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n944), .ZN(n946) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1040 ( .A1(n947), .A2(G29), .ZN(n948) );
  XOR2_X1 U1041 ( .A(KEYINPUT115), .B(n948), .Z(n1033) );
  XOR2_X1 U1042 ( .A(G1996), .B(G32), .Z(n949) );
  NAND2_X1 U1043 ( .A1(n949), .A2(G28), .ZN(n952) );
  XNOR2_X1 U1044 ( .A(KEYINPUT116), .B(G2072), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(G33), .B(n950), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n960) );
  XOR2_X1 U1047 ( .A(G2067), .B(G26), .Z(n955) );
  XNOR2_X1 U1048 ( .A(n953), .B(G25), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n958) );
  XOR2_X1 U1050 ( .A(G27), .B(n956), .Z(n957) );
  NOR2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1052 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(KEYINPUT53), .B(n961), .ZN(n966) );
  XOR2_X1 U1054 ( .A(KEYINPUT118), .B(KEYINPUT117), .Z(n963) );
  XNOR2_X1 U1055 ( .A(G2084), .B(G34), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(n963), .B(n962), .ZN(n964) );
  XOR2_X1 U1057 ( .A(KEYINPUT54), .B(n964), .Z(n965) );
  NAND2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n968) );
  XNOR2_X1 U1059 ( .A(G35), .B(G2090), .ZN(n967) );
  NOR2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(KEYINPUT55), .B(n969), .ZN(n971) );
  INV_X1 U1062 ( .A(G29), .ZN(n970) );
  NAND2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1064 ( .A1(n972), .A2(G11), .ZN(n1031) );
  XNOR2_X1 U1065 ( .A(G16), .B(KEYINPUT56), .ZN(n1001) );
  XNOR2_X1 U1066 ( .A(n973), .B(G1956), .ZN(n983) );
  XNOR2_X1 U1067 ( .A(G1348), .B(KEYINPUT120), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n975), .B(n974), .ZN(n978) );
  XNOR2_X1 U1069 ( .A(G171), .B(G1961), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(n976), .B(KEYINPUT121), .ZN(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1072 ( .A(KEYINPUT122), .B(n979), .Z(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(G1341), .B(n984), .ZN(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n999) );
  XOR2_X1 U1077 ( .A(G168), .B(G1966), .Z(n987) );
  NOR2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1079 ( .A(KEYINPUT119), .B(n989), .Z(n990) );
  XNOR2_X1 U1080 ( .A(KEYINPUT57), .B(n990), .ZN(n997) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n994) );
  AND2_X1 U1082 ( .A1(G303), .A2(G1971), .ZN(n993) );
  NOR2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(KEYINPUT123), .B(n995), .ZN(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1029) );
  INV_X1 U1088 ( .A(G16), .ZN(n1027) );
  XOR2_X1 U1089 ( .A(G1348), .B(KEYINPUT59), .Z(n1002) );
  XNOR2_X1 U1090 ( .A(G4), .B(n1002), .ZN(n1011) );
  XNOR2_X1 U1091 ( .A(G1981), .B(G6), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(n1003), .B(KEYINPUT124), .ZN(n1008) );
  XOR2_X1 U1093 ( .A(G1341), .B(G19), .Z(n1006) );
  XNOR2_X1 U1094 ( .A(n1004), .B(G20), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(n1009), .B(KEYINPUT125), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(KEYINPUT60), .B(n1012), .ZN(n1016) );
  XNOR2_X1 U1100 ( .A(G1966), .B(G21), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(G1961), .B(G5), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1024) );
  XNOR2_X1 U1104 ( .A(G1986), .B(G24), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(G23), .B(G1976), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1021) );
  XOR2_X1 U1107 ( .A(G1971), .B(KEYINPUT126), .Z(n1019) );
  XNOR2_X1 U1108 ( .A(G22), .B(n1019), .ZN(n1020) );
  NAND2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1110 ( .A(KEYINPUT58), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1112 ( .A(KEYINPUT61), .B(n1025), .ZN(n1026) );
  NAND2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1115 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1116 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1117 ( .A(n1034), .B(KEYINPUT62), .ZN(n1035) );
  XNOR2_X1 U1118 ( .A(KEYINPUT127), .B(n1035), .ZN(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

