//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT32), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT70), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT28), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT11), .ZN(new_n191));
  OR2_X1    g005(.A1(KEYINPUT65), .A2(G134), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT65), .A2(G134), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(G137), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G137), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n191), .B1(new_n194), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n192), .A2(new_n193), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  AOI21_X1  g014(.A(KEYINPUT11), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(G131), .B1(new_n198), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  AND2_X1   g017(.A1(KEYINPUT65), .A2(G134), .ZN(new_n204));
  NOR2_X1   g018(.A1(KEYINPUT65), .A2(G134), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n191), .B1(new_n206), .B2(G137), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n196), .B1(new_n206), .B2(G137), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n203), .B(new_n207), .C1(new_n208), .C2(new_n191), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n202), .A2(new_n209), .A3(KEYINPUT66), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n211), .B(G131), .C1(new_n198), .C2(new_n201), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  AND3_X1   g029(.A1(new_n215), .A2(KEYINPUT64), .A3(G146), .ZN(new_n216));
  AOI21_X1  g030(.A(KEYINPUT64), .B1(new_n215), .B2(G146), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n214), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(KEYINPUT0), .A2(G128), .ZN(new_n219));
  NOR2_X1   g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n215), .A2(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n214), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n218), .A2(new_n221), .B1(new_n224), .B2(new_n219), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n210), .A2(new_n212), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n206), .A2(G137), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n200), .A2(G134), .ZN(new_n228));
  OAI21_X1  g042(.A(G131), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n209), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  NOR3_X1   g045(.A1(new_n223), .A2(KEYINPUT1), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n215), .A2(G146), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT1), .ZN(new_n235));
  OAI21_X1  g049(.A(G128), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT67), .B1(new_n218), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT64), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n238), .B1(new_n213), .B2(G143), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n215), .A2(KEYINPUT64), .A3(G146), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n234), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n231), .B1(new_n214), .B2(KEYINPUT1), .ZN(new_n243));
  NOR3_X1   g057(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n233), .B1(new_n237), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n230), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n226), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G119), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G116), .ZN(new_n249));
  INV_X1    g063(.A(G116), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G119), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT2), .B(G113), .ZN(new_n253));
  XOR2_X1   g067(.A(new_n252), .B(new_n253), .Z(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n247), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n245), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n218), .A2(KEYINPUT67), .A3(new_n236), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n242), .B1(new_n241), .B2(new_n243), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n232), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT68), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n258), .A2(new_n230), .A3(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(new_n254), .A3(new_n226), .ZN(new_n264));
  AOI211_X1 g078(.A(new_n189), .B(new_n190), .C1(new_n256), .C2(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n190), .B1(new_n256), .B2(new_n264), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT70), .B1(new_n264), .B2(new_n190), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(G237), .A2(G953), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G210), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(KEYINPUT27), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT26), .B(G101), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT30), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n247), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n263), .A2(KEYINPUT30), .A3(new_n226), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(new_n278), .A3(new_n255), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n275), .A2(KEYINPUT31), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(KEYINPUT31), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n275), .A2(KEYINPUT69), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n279), .A2(new_n282), .A3(new_n264), .A4(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n279), .A2(new_n264), .A3(new_n283), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n281), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n269), .A2(new_n275), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(G472), .A2(G902), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n187), .B(new_n188), .C1(new_n287), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n286), .A2(new_n284), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n256), .A2(new_n264), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n264), .A2(new_n190), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n189), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n293), .B(new_n275), .C1(new_n266), .C2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n289), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT71), .B1(new_n297), .B2(KEYINPUT32), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n290), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n293), .B(new_n274), .C1(new_n266), .C2(new_n295), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n279), .A2(new_n275), .A3(new_n264), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT29), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G902), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n263), .A2(new_n226), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n304), .B(new_n254), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n294), .B1(new_n305), .B2(new_n190), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n274), .A2(KEYINPUT29), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n303), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G472), .B1(new_n302), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n291), .A2(new_n296), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(KEYINPUT32), .A3(new_n288), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT72), .B1(new_n299), .B2(new_n312), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n309), .A2(new_n311), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT72), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n314), .A2(new_n315), .A3(new_n298), .A4(new_n290), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT23), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n318), .B1(new_n248), .B2(G128), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n231), .A2(KEYINPUT23), .A3(G119), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n319), .B(new_n320), .C1(G119), .C2(new_n231), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G110), .ZN(new_n322));
  XOR2_X1   g136(.A(G119), .B(G128), .Z(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT24), .B(G110), .ZN(new_n324));
  XNOR2_X1  g138(.A(G125), .B(G140), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT16), .ZN(new_n326));
  INV_X1    g140(.A(G140), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G125), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n326), .B(KEYINPUT73), .C1(KEYINPUT16), .C2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n325), .A2(new_n330), .A3(KEYINPUT16), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n331), .A3(new_n213), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n213), .B1(new_n329), .B2(new_n331), .ZN(new_n334));
  OAI221_X1 g148(.A(new_n322), .B1(new_n323), .B2(new_n324), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n329), .A2(new_n331), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G146), .ZN(new_n337));
  INV_X1    g151(.A(G125), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G140), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n328), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT75), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n325), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n343), .A3(new_n213), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n344), .A2(KEYINPUT76), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(KEYINPUT76), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n323), .A2(new_n324), .ZN(new_n347));
  XOR2_X1   g161(.A(new_n347), .B(KEYINPUT74), .Z(new_n348));
  NOR2_X1   g162(.A1(new_n321), .A2(G110), .ZN(new_n349));
  OAI221_X1 g163(.A(new_n337), .B1(new_n345), .B2(new_n346), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n335), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT22), .B(G137), .ZN(new_n352));
  INV_X1    g166(.A(G953), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n353), .A2(G221), .A3(G234), .ZN(new_n354));
  XOR2_X1   g168(.A(new_n352), .B(new_n354), .Z(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n335), .A2(new_n350), .A3(new_n355), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n303), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT25), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n359), .B(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G217), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(G234), .B2(new_n303), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(G902), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n357), .A2(new_n358), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G221), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT9), .B(G234), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n369), .B1(new_n371), .B2(new_n303), .ZN(new_n372));
  INV_X1    g186(.A(G469), .ZN(new_n373));
  XNOR2_X1  g187(.A(G110), .B(G140), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n353), .A2(G227), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n378));
  INV_X1    g192(.A(G104), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT3), .B1(new_n379), .B2(G107), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT3), .ZN(new_n381));
  INV_X1    g195(.A(G107), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(G104), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n380), .B(new_n383), .C1(G104), .C2(new_n382), .ZN(new_n384));
  XOR2_X1   g198(.A(KEYINPUT77), .B(G101), .Z(new_n385));
  OR2_X1    g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(G101), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n378), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT4), .B1(new_n384), .B2(G101), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n225), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n379), .A2(G107), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n382), .A2(G104), .ZN(new_n393));
  OAI21_X1  g207(.A(G101), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n386), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n232), .B1(new_n223), .B2(new_n236), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI22_X1  g211(.A1(new_n390), .A2(new_n391), .B1(new_n397), .B2(KEYINPUT10), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n259), .A2(new_n260), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT68), .B1(new_n400), .B2(new_n233), .ZN(new_n401));
  AOI211_X1 g215(.A(new_n257), .B(new_n232), .C1(new_n259), .C2(new_n260), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT10), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n395), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT78), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n258), .A2(new_n262), .A3(new_n405), .A4(KEYINPUT78), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n399), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n210), .A2(new_n212), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(KEYINPUT79), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT79), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n258), .A2(new_n262), .A3(new_n405), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT78), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n398), .B1(new_n416), .B2(new_n407), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n413), .B1(new_n417), .B2(new_n410), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n410), .B(new_n399), .C1(new_n406), .C2(new_n408), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n377), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n377), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n261), .A2(new_n395), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n423), .B1(new_n395), .B2(new_n396), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n411), .A2(new_n424), .A3(KEYINPUT12), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT12), .ZN(new_n426));
  INV_X1    g240(.A(new_n424), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n426), .B1(new_n427), .B2(new_n410), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n422), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n373), .B(new_n303), .C1(new_n421), .C2(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n373), .A2(new_n303), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n428), .A2(new_n425), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n377), .B1(new_n420), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n422), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n433), .B1(new_n419), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n431), .B1(new_n435), .B2(G469), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n372), .B1(new_n430), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G214), .B1(G237), .B2(G902), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(G210), .B1(G237), .B2(G902), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(KEYINPUT82), .ZN(new_n441));
  XNOR2_X1  g255(.A(G110), .B(G122), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n255), .B1(new_n388), .B2(new_n389), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n252), .A2(new_n253), .ZN(new_n446));
  INV_X1    g260(.A(new_n252), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT5), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n449));
  INV_X1    g263(.A(G113), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n446), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n386), .A3(new_n394), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT80), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT80), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n452), .A2(new_n455), .A3(new_n386), .A4(new_n394), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n443), .B1(new_n445), .B2(new_n457), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n444), .A2(new_n454), .A3(new_n442), .A4(new_n456), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(KEYINPUT6), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n261), .A2(new_n338), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n391), .A2(G125), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G224), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(G953), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n463), .A2(new_n465), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT6), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n469), .B(new_n443), .C1(new_n445), .C2(new_n457), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n460), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n465), .A2(KEYINPUT7), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n472), .B1(new_n466), .B2(new_n467), .ZN(new_n473));
  XOR2_X1   g287(.A(new_n442), .B(KEYINPUT8), .Z(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(new_n395), .B2(new_n452), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT81), .ZN(new_n476));
  AOI211_X1 g290(.A(new_n450), .B(new_n449), .C1(new_n448), .C2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n447), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n446), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n475), .B1(new_n479), .B2(new_n395), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n463), .A2(new_n472), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n459), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n303), .B1(new_n473), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n441), .B1(new_n471), .B2(new_n483), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n473), .A2(new_n482), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n460), .A2(new_n468), .A3(new_n470), .ZN(new_n486));
  INV_X1    g300(.A(new_n441), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n485), .A2(new_n486), .A3(new_n303), .A4(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n439), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G478), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(KEYINPUT15), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n231), .A2(G143), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n215), .A2(G128), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n199), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n492), .ZN(new_n495));
  INV_X1    g309(.A(new_n493), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n206), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n250), .A2(KEYINPUT14), .A3(G122), .ZN(new_n499));
  XOR2_X1   g313(.A(G116), .B(G122), .Z(new_n500));
  OAI211_X1 g314(.A(G107), .B(new_n499), .C1(new_n500), .C2(KEYINPUT14), .ZN(new_n501));
  XNOR2_X1  g315(.A(G116), .B(G122), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n382), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n498), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT89), .ZN(new_n505));
  INV_X1    g319(.A(new_n503), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n502), .A2(new_n382), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n500), .A2(G107), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n503), .A3(KEYINPUT89), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n497), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT13), .B1(new_n215), .B2(G128), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT90), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n493), .B1(KEYINPUT13), .B2(new_n492), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n195), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n504), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n370), .A2(new_n362), .A3(G953), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n504), .B(new_n517), .C1(new_n511), .C2(new_n515), .ZN(new_n520));
  AOI21_X1  g334(.A(G902), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT92), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT91), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n519), .A2(new_n520), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n525), .A2(KEYINPUT91), .A3(G902), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n491), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n523), .B1(KEYINPUT15), .B2(new_n490), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n333), .A2(new_n334), .ZN(new_n531));
  INV_X1    g345(.A(G237), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(new_n353), .A3(G214), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(KEYINPUT83), .A3(new_n215), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n215), .A2(KEYINPUT83), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(G214), .A3(new_n270), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT84), .B1(new_n537), .B2(G131), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT84), .ZN(new_n539));
  AOI211_X1 g353(.A(new_n539), .B(new_n203), .C1(new_n534), .C2(new_n536), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT17), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n538), .A2(new_n540), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n534), .A2(new_n203), .A3(new_n536), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n531), .B(new_n541), .C1(KEYINPUT17), .C2(new_n544), .ZN(new_n545));
  OAI22_X1  g359(.A1(new_n345), .A2(new_n346), .B1(new_n213), .B2(new_n325), .ZN(new_n546));
  NAND2_X1  g360(.A1(KEYINPUT18), .A2(G131), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n537), .B(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(G113), .B(G122), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT87), .B(G104), .ZN(new_n552));
  XOR2_X1   g366(.A(new_n551), .B(new_n552), .Z(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT88), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n545), .A2(new_n549), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n555), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(new_n303), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G475), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n334), .B1(new_n542), .B2(new_n543), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT19), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n341), .A2(new_n343), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n340), .A2(KEYINPUT19), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT85), .B1(new_n566), .B2(G146), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT85), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n564), .A2(new_n568), .A3(new_n213), .A4(new_n565), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n562), .A2(new_n570), .B1(new_n546), .B2(new_n548), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT86), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n554), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n562), .A2(new_n570), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n574), .A2(new_n572), .A3(new_n549), .ZN(new_n575));
  OAI22_X1  g389(.A1(new_n573), .A2(new_n575), .B1(new_n558), .B2(new_n554), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT20), .ZN(new_n577));
  NOR2_X1   g391(.A1(G475), .A2(G902), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n577), .B1(new_n576), .B2(new_n578), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n561), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(G234), .A2(G237), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(G952), .A3(new_n353), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT93), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n582), .A2(G902), .A3(G953), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT21), .B(G898), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(KEYINPUT94), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n581), .A2(new_n590), .ZN(new_n591));
  AND4_X1   g405(.A1(new_n437), .A2(new_n489), .A3(new_n530), .A4(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n317), .A2(new_n368), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(new_n385), .ZN(G3));
  NAND2_X1  g408(.A1(new_n437), .A2(new_n368), .ZN(new_n595));
  OAI211_X1 g409(.A(KEYINPUT95), .B(G472), .C1(new_n287), .C2(G902), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT95), .ZN(new_n597));
  AOI21_X1  g411(.A(G902), .B1(new_n291), .B2(new_n296), .ZN(new_n598));
  INV_X1    g412(.A(G472), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n297), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n596), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT96), .B1(new_n595), .B2(new_n602), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n596), .A2(new_n600), .A3(new_n601), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT96), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n604), .A2(new_n605), .A3(new_n368), .A4(new_n437), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n521), .A2(new_n490), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n490), .B2(new_n303), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n516), .B2(KEYINPUT97), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n525), .B(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n609), .B1(new_n612), .B2(G478), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n489), .A2(new_n581), .A3(new_n589), .A4(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n607), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT34), .B(G104), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  NAND2_X1  g431(.A1(new_n576), .A2(new_n578), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(KEYINPUT20), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n619), .A2(new_n620), .B1(G475), .B2(new_n560), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n621), .A2(new_n489), .A3(new_n529), .A4(new_n589), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n607), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT35), .B(G107), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G9));
  OAI21_X1  g439(.A(new_n351), .B1(KEYINPUT36), .B2(new_n356), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n356), .A2(KEYINPUT36), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n335), .A2(new_n350), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n626), .A2(new_n365), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT98), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n364), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n529), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n591), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n635), .A2(new_n437), .A3(new_n489), .A4(new_n604), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT37), .B(G110), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT99), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n636), .B(new_n638), .ZN(G12));
  NAND2_X1  g453(.A1(new_n621), .A2(new_n529), .ZN(new_n640));
  INV_X1    g454(.A(G900), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n585), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n584), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n644), .A2(new_n437), .A3(new_n489), .A4(new_n631), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n313), .B2(new_n316), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(new_n231), .ZN(G30));
  NAND2_X1  g461(.A1(new_n430), .A2(new_n436), .ZN(new_n648));
  INV_X1    g462(.A(new_n372), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n643), .B(KEYINPUT39), .Z(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(KEYINPUT40), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n530), .A2(new_n621), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n654), .A2(new_n632), .A3(new_n438), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n484), .A2(new_n488), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT38), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT40), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n437), .A2(new_n660), .A3(new_n651), .ZN(new_n661));
  AOI21_X1  g475(.A(G902), .B1(new_n305), .B2(new_n275), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n279), .A2(new_n264), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n274), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G472), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n290), .A2(new_n298), .A3(new_n311), .A4(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n653), .A2(new_n659), .A3(new_n661), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G143), .ZN(G45));
  INV_X1    g483(.A(new_n643), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n581), .A2(new_n613), .A3(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n437), .A2(new_n489), .A3(new_n631), .A4(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n313), .B2(new_n316), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT100), .B(G146), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G48));
  AOI21_X1  g489(.A(new_n367), .B1(new_n313), .B2(new_n316), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n373), .A2(KEYINPUT101), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n421), .A2(new_n429), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n677), .B1(new_n678), .B2(G902), .ZN(new_n679));
  OAI221_X1 g493(.A(new_n303), .B1(KEYINPUT101), .B2(new_n373), .C1(new_n421), .C2(new_n429), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(new_n649), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n614), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT41), .B(G113), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G15));
  NOR2_X1   g499(.A1(new_n681), .A2(new_n622), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n676), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G116), .ZN(G18));
  NAND4_X1  g502(.A1(new_n679), .A2(new_n649), .A3(new_n489), .A4(new_n680), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n317), .A2(new_n635), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G119), .ZN(G21));
  OAI21_X1  g506(.A(G472), .B1(new_n287), .B2(G902), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n306), .A2(new_n275), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n291), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n288), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n368), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n681), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n654), .A2(KEYINPUT102), .A3(new_n489), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n489), .A2(new_n529), .A3(new_n581), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n698), .A2(new_n589), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT103), .B(G122), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G24));
  NAND4_X1  g520(.A1(new_n671), .A2(new_n693), .A3(new_n631), .A4(new_n696), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n689), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n338), .ZN(G27));
  AND3_X1   g523(.A1(new_n484), .A2(new_n438), .A3(new_n488), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n710), .B1(new_n437), .B2(new_n711), .ZN(new_n712));
  AOI211_X1 g526(.A(KEYINPUT104), .B(new_n372), .C1(new_n430), .C2(new_n436), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n601), .A2(new_n188), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n367), .B1(new_n314), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n671), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT42), .ZN(new_n718));
  INV_X1    g532(.A(new_n671), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(KEYINPUT42), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n676), .A2(new_n714), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n203), .ZN(G33));
  NAND3_X1  g537(.A1(new_n676), .A2(new_n644), .A3(new_n714), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT105), .B(G134), .Z(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G36));
  INV_X1    g540(.A(new_n710), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n561), .B(new_n613), .C1(new_n579), .C2(new_n580), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT107), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n728), .A2(new_n729), .A3(KEYINPUT43), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT43), .B1(new_n728), .B2(new_n729), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n602), .A3(new_n631), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n727), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n730), .A2(new_n731), .A3(new_n632), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n736), .A2(KEYINPUT108), .A3(KEYINPUT44), .A4(new_n602), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n732), .A2(KEYINPUT44), .A3(new_n602), .A4(new_n631), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n735), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n419), .A2(new_n434), .ZN(new_n742));
  INV_X1    g556(.A(new_n433), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(KEYINPUT45), .A3(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n422), .B1(new_n418), .B2(new_n412), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n745), .B1(new_n746), .B2(new_n433), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n744), .A2(new_n747), .A3(G469), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT106), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT106), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n744), .A2(new_n747), .A3(new_n750), .A4(G469), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n431), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n430), .B1(new_n752), .B2(KEYINPUT46), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT46), .ZN(new_n754));
  AOI211_X1 g568(.A(new_n754), .B(new_n431), .C1(new_n749), .C2(new_n751), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n649), .B(new_n651), .C1(new_n753), .C2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n741), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n200), .ZN(G39));
  INV_X1    g572(.A(KEYINPUT47), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n759), .B(new_n649), .C1(new_n753), .C2(new_n755), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n431), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n742), .A2(new_n743), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n373), .B1(new_n764), .B2(new_n745), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n750), .B1(new_n765), .B2(new_n744), .ZN(new_n766));
  INV_X1    g580(.A(new_n751), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n763), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n754), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n752), .A2(KEYINPUT46), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n430), .A3(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(KEYINPUT109), .A3(new_n759), .A4(new_n649), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n762), .A2(new_n772), .ZN(new_n773));
  NOR4_X1   g587(.A1(new_n317), .A2(new_n368), .A3(new_n719), .A4(new_n727), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n649), .B1(new_n753), .B2(new_n755), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT110), .B1(new_n775), .B2(KEYINPUT47), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n775), .A2(KEYINPUT110), .A3(KEYINPUT47), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n773), .B(new_n774), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G140), .ZN(G42));
  AND4_X1   g593(.A1(new_n317), .A2(new_n714), .A3(new_n368), .A4(new_n644), .ZN(new_n780));
  AND4_X1   g594(.A1(new_n530), .A2(new_n631), .A3(new_n621), .A4(new_n710), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n781), .A2(new_n437), .A3(new_n670), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n317), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n727), .B1(new_n650), .B2(KEYINPUT104), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n693), .A2(new_n631), .A3(new_n696), .ZN(new_n785));
  INV_X1    g599(.A(new_n713), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n784), .A2(new_n785), .A3(new_n671), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT113), .B1(new_n780), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n724), .A2(new_n790), .A3(new_n787), .A4(new_n783), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n722), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n683), .A2(new_n687), .A3(new_n691), .A4(new_n704), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n614), .A2(KEYINPUT111), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n614), .A2(KEYINPUT111), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n622), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n603), .A2(new_n606), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n593), .A2(new_n797), .A3(new_n636), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n593), .A2(new_n797), .A3(KEYINPUT112), .A4(new_n636), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n793), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n646), .A2(new_n673), .A3(new_n708), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n650), .A2(new_n643), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n804), .A2(new_n703), .A3(new_n632), .A4(new_n667), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n803), .A2(KEYINPUT52), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n645), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n708), .B1(new_n317), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n673), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n809), .A3(new_n805), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n806), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n792), .A2(new_n802), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n817));
  NOR2_X1   g631(.A1(KEYINPUT114), .A2(KEYINPUT52), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(KEYINPUT114), .A2(KEYINPUT52), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n820), .B1(new_n803), .B2(new_n805), .ZN(new_n821));
  AND4_X1   g635(.A1(new_n809), .A2(new_n808), .A3(new_n805), .A4(new_n820), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n819), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n823), .A2(KEYINPUT53), .A3(new_n792), .A4(new_n802), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n816), .A2(new_n817), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n823), .A2(new_n802), .A3(new_n792), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n826), .A2(new_n827), .A3(new_n815), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n827), .B1(new_n826), .B2(new_n815), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n814), .A2(new_n815), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n825), .B1(new_n831), .B2(new_n817), .ZN(new_n832));
  OR3_X1    g646(.A1(new_n730), .A2(new_n731), .A3(new_n584), .ZN(new_n833));
  INV_X1    g647(.A(new_n658), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n833), .A2(new_n438), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n698), .ZN(new_n836));
  XOR2_X1   g650(.A(new_n836), .B(KEYINPUT50), .Z(new_n837));
  OR2_X1    g651(.A1(new_n681), .A2(new_n727), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n838), .A2(new_n367), .A3(new_n584), .A4(new_n667), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n581), .A2(new_n613), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n838), .A2(new_n833), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n785), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n837), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT51), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n777), .A2(new_n776), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n762), .A2(new_n772), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n679), .A2(new_n680), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n850), .A2(new_n649), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT117), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n833), .A2(new_n697), .A3(new_n727), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n849), .A2(KEYINPUT117), .A3(new_n851), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n846), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n842), .A2(new_n716), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n857), .B(KEYINPUT48), .Z(new_n858));
  NOR3_X1   g672(.A1(new_n833), .A2(new_n689), .A3(new_n697), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n859), .B(KEYINPUT118), .Z(new_n860));
  NAND2_X1  g674(.A1(new_n581), .A2(new_n613), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n839), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(G952), .A3(new_n353), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n858), .A2(new_n860), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n849), .A2(KEYINPUT116), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT116), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(new_n847), .B2(new_n848), .ZN(new_n868));
  INV_X1    g682(.A(new_n851), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n844), .B1(new_n870), .B2(new_n853), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n856), .B(new_n865), .C1(new_n871), .C2(KEYINPUT51), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n832), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(G952), .A2(G953), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n368), .A2(new_n649), .A3(new_n438), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n834), .A2(new_n875), .A3(new_n728), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n850), .A2(KEYINPUT49), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n850), .A2(KEYINPUT49), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  OAI22_X1  g693(.A1(new_n873), .A2(new_n874), .B1(new_n667), .B2(new_n879), .ZN(G75));
  NOR2_X1   g694(.A1(new_n353), .A2(G952), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT119), .Z(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n303), .B1(new_n816), .B2(new_n824), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT56), .B1(new_n884), .B2(new_n441), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n460), .A2(new_n470), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n886), .A2(new_n468), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(new_n471), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(KEYINPUT55), .Z(new_n889));
  OR2_X1    g703(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n885), .A2(new_n889), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n883), .B1(new_n890), .B2(new_n891), .ZN(G51));
  AND3_X1   g706(.A1(new_n816), .A2(new_n817), .A3(new_n824), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n817), .B1(new_n816), .B2(new_n824), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n431), .B(KEYINPUT57), .Z(new_n896));
  OAI22_X1  g710(.A1(new_n895), .A2(new_n896), .B1(new_n421), .B2(new_n429), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n884), .A2(new_n751), .A3(new_n749), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n881), .B1(new_n897), .B2(new_n898), .ZN(G54));
  AND2_X1   g713(.A1(KEYINPUT58), .A2(G475), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n884), .A2(new_n576), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n576), .B1(new_n884), .B2(new_n900), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n901), .A2(new_n902), .A3(new_n881), .ZN(G60));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n612), .B(KEYINPUT120), .Z(new_n905));
  XNOR2_X1  g719(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n490), .A2(new_n303), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n906), .B(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n816), .A2(new_n824), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT54), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n909), .B1(new_n911), .B2(new_n825), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n904), .B1(new_n912), .B2(new_n883), .ZN(new_n913));
  OAI211_X1 g727(.A(KEYINPUT122), .B(new_n882), .C1(new_n895), .C2(new_n909), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n905), .B1(new_n832), .B2(new_n908), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n915), .A2(new_n916), .ZN(G63));
  NAND2_X1  g731(.A1(G217), .A2(G902), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT60), .Z(new_n919));
  NAND2_X1  g733(.A1(new_n910), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n357), .A2(new_n358), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n626), .A2(new_n628), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n922), .B(new_n882), .C1(new_n923), .C2(new_n920), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n924), .B(new_n925), .ZN(G66));
  OAI21_X1  g740(.A(G953), .B1(new_n586), .B2(new_n464), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(new_n802), .B2(G953), .ZN(new_n928));
  INV_X1    g742(.A(new_n886), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(G898), .B2(new_n353), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n928), .B(new_n930), .ZN(G69));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n353), .B1(G227), .B2(G900), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n277), .A2(new_n278), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n566), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n437), .A2(new_n651), .ZN(new_n937));
  AOI211_X1 g751(.A(new_n727), .B(new_n937), .C1(new_n861), .C2(new_n640), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n676), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n741), .B2(new_n756), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n808), .A2(new_n809), .A3(new_n668), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n940), .B1(KEYINPUT62), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT62), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n803), .A2(new_n943), .A3(new_n944), .A4(new_n668), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT123), .B1(new_n941), .B2(KEYINPUT62), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n778), .A2(new_n942), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  AOI211_X1 g761(.A(KEYINPUT124), .B(new_n936), .C1(new_n947), .C2(new_n353), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT110), .ZN(new_n950));
  INV_X1    g764(.A(new_n430), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n768), .B2(new_n754), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n372), .B1(new_n952), .B2(new_n770), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n950), .B1(new_n953), .B2(new_n759), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n775), .A2(KEYINPUT110), .A3(KEYINPUT47), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n956), .A2(new_n773), .A3(new_n774), .ZN(new_n957));
  INV_X1    g771(.A(new_n940), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n941), .A2(KEYINPUT62), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n958), .A2(new_n946), .A3(new_n945), .A4(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n353), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n936), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n949), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n948), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n703), .A2(new_n716), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n756), .B1(new_n741), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n803), .A2(new_n724), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n966), .A2(new_n967), .A3(new_n722), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n778), .A2(new_n968), .A3(new_n353), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n962), .B1(G900), .B2(G953), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(KEYINPUT125), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n969), .A2(new_n973), .A3(new_n970), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n934), .B1(new_n964), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n961), .A2(new_n962), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(KEYINPUT124), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n961), .A2(new_n949), .A3(new_n962), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n933), .B1(new_n969), .B2(new_n970), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n932), .B1(new_n976), .B2(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n978), .A2(new_n979), .A3(new_n972), .A4(new_n974), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n933), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n964), .A2(new_n980), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n984), .A2(KEYINPUT126), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n982), .A2(new_n986), .ZN(G72));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT63), .Z(new_n989));
  NAND3_X1  g803(.A1(new_n664), .A2(new_n301), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n831), .A2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n802), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n947), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n664), .B1(new_n993), .B2(new_n989), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n301), .B(KEYINPUT127), .Z(new_n995));
  NAND3_X1  g809(.A1(new_n778), .A2(new_n968), .A3(new_n802), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n995), .B1(new_n996), .B2(new_n989), .ZN(new_n997));
  NOR4_X1   g811(.A1(new_n991), .A2(new_n881), .A3(new_n994), .A4(new_n997), .ZN(G57));
endmodule


