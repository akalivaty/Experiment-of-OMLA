//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n549, new_n550, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1240, new_n1241, new_n1242, new_n1243;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT66), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  XOR2_X1   g026(.A(KEYINPUT67), .B(KEYINPUT68), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n451), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT69), .ZN(G319));
  OR2_X1    g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  AOI21_X1  g035(.A(G2105), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G137), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n463), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT70), .ZN(G160));
  NAND2_X1  g048(.A1(new_n461), .A2(G136), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n463), .B1(new_n459), .B2(new_n460), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  INV_X1    g055(.A(G138), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n482), .B1(new_n467), .B2(new_n468), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT4), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n482), .B(new_n485), .C1(new_n468), .C2(new_n467), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT71), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G114), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT71), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n489), .A2(new_n491), .A3(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n475), .A2(G126), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n487), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT72), .B1(new_n499), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT73), .B1(new_n502), .B2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(new_n499), .A3(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n504), .A2(new_n508), .A3(G62), .ZN(new_n509));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n498), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n504), .A2(new_n508), .A3(G88), .A4(new_n514), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n502), .B1(new_n512), .B2(new_n513), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n511), .A2(new_n518), .ZN(G166));
  AOI22_X1  g094(.A1(new_n500), .A2(new_n503), .B1(new_n505), .B2(new_n507), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(G89), .A3(new_n514), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n525));
  AOI22_X1  g100(.A1(G51), .A2(new_n516), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n521), .A2(new_n522), .A3(new_n526), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  NAND2_X1  g103(.A1(G77), .A2(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n504), .A2(new_n508), .ZN(new_n530));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G651), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n504), .A2(new_n508), .A3(new_n514), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT74), .B(G90), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n534), .A2(new_n535), .B1(G52), .B2(new_n516), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n533), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  NAND4_X1  g113(.A1(new_n504), .A2(new_n508), .A3(G81), .A4(new_n514), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT75), .B(G43), .Z(new_n540));
  NAND2_X1  g115(.A1(new_n516), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n504), .A2(new_n508), .A3(G56), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n542), .B1(G651), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(G188));
  NAND2_X1  g126(.A1(new_n534), .A2(G91), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n520), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n553), .B2(new_n498), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n555), .B1(new_n516), .B2(G53), .ZN(new_n556));
  AND2_X1   g131(.A1(KEYINPUT6), .A2(G651), .ZN(new_n557));
  NOR2_X1   g132(.A1(KEYINPUT6), .A2(G651), .ZN(new_n558));
  OAI211_X1 g133(.A(G53), .B(G543), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT76), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n514), .A2(new_n555), .A3(G53), .A4(G543), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NOR3_X1   g141(.A1(new_n554), .A2(new_n566), .A3(KEYINPUT77), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n568));
  AND3_X1   g143(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n564), .B1(new_n562), .B2(new_n563), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n530), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(G651), .B1(G91), .B2(new_n534), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n568), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n567), .A2(new_n576), .ZN(G299));
  INV_X1    g152(.A(new_n518), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n509), .A2(new_n510), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G651), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(KEYINPUT78), .B1(new_n511), .B2(new_n518), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(G303));
  OAI21_X1  g159(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n504), .A2(new_n508), .A3(G87), .A4(new_n514), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n516), .A2(G49), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(new_n516), .A2(G48), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n530), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n590), .B1(new_n593), .B2(G651), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n504), .A2(new_n508), .A3(G86), .A4(new_n514), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(KEYINPUT79), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n520), .A2(new_n597), .A3(G86), .A4(new_n514), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n594), .A2(new_n596), .A3(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n534), .A2(G85), .B1(G47), .B2(new_n516), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  OAI21_X1  g176(.A(G651), .B1(new_n601), .B2(KEYINPUT80), .ZN(new_n602));
  NAND2_X1  g177(.A1(G72), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G60), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n530), .B2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT80), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n602), .B2(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n520), .A2(new_n514), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n534), .A2(KEYINPUT10), .A3(G92), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n613), .A2(new_n614), .B1(G54), .B2(new_n516), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  INV_X1    g191(.A(G79), .ZN(new_n617));
  OAI22_X1  g192(.A1(new_n530), .A2(new_n616), .B1(new_n617), .B2(new_n502), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT81), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI221_X1 g195(.A(KEYINPUT81), .B1(new_n617), .B2(new_n502), .C1(new_n530), .C2(new_n616), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n620), .A2(G651), .A3(new_n621), .ZN(new_n622));
  AND2_X1   g197(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n609), .B1(new_n623), .B2(G868), .ZN(G284));
  OAI21_X1  g199(.A(new_n609), .B1(new_n623), .B2(G868), .ZN(G321));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NAND2_X1  g201(.A1(G299), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n626), .B2(G168), .ZN(G297));
  OAI21_X1  g203(.A(new_n627), .B1(new_n626), .B2(G168), .ZN(G280));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n623), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n623), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g210(.A(KEYINPUT3), .B(G2104), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(new_n464), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT13), .ZN(new_n639));
  INV_X1    g214(.A(G2100), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n461), .A2(G135), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n475), .A2(G123), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n463), .A2(G111), .ZN(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n643), .B(new_n644), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(G2096), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n641), .A2(new_n642), .A3(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(KEYINPUT14), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  AND3_X1   g237(.A1(new_n662), .A2(KEYINPUT82), .A3(new_n651), .ZN(new_n663));
  AOI21_X1  g238(.A(KEYINPUT82), .B1(new_n662), .B2(new_n651), .ZN(new_n664));
  OAI221_X1 g239(.A(G14), .B1(new_n651), .B2(new_n662), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT83), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(G401));
  INV_X1    g244(.A(KEYINPUT18), .ZN(new_n670));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(KEYINPUT17), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n671), .A2(new_n672), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n670), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G2100), .ZN(new_n677));
  XOR2_X1   g252(.A(G2072), .B(G2078), .Z(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n673), .B2(KEYINPUT18), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(new_n648), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n677), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(G227));
  XOR2_X1   g257(.A(G1991), .B(G1996), .Z(new_n683));
  XNOR2_X1  g258(.A(G1956), .B(G2474), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT85), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1961), .B(G1966), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n692), .B(new_n693), .Z(new_n694));
  OR2_X1    g269(.A1(new_n685), .A2(new_n687), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n695), .A2(new_n691), .ZN(new_n696));
  AND3_X1   g271(.A1(new_n695), .A2(new_n688), .A3(new_n691), .ZN(new_n697));
  NOR3_X1   g272(.A1(new_n694), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n683), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n698), .A2(new_n699), .ZN(new_n703));
  INV_X1    g278(.A(new_n683), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n698), .A2(new_n699), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1981), .B(G1986), .ZN(new_n707));
  AND3_X1   g282(.A1(new_n702), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n707), .B1(new_n702), .B2(new_n706), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(G229));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n711), .A2(G32), .ZN(new_n712));
  NAND3_X1  g287(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT93), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT26), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n461), .A2(G141), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n475), .A2(G129), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n464), .A2(G105), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n720), .A2(KEYINPUT94), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(KEYINPUT94), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n712), .B1(new_n723), .B2(G29), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT27), .B(G1996), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NOR2_X1   g302(.A1(G168), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n727), .B2(G21), .ZN(new_n729));
  INV_X1    g304(.A(G1966), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n711), .A2(G27), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G164), .B2(new_n711), .ZN(new_n733));
  INV_X1    g308(.A(G2078), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(G29), .A2(G33), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT92), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n636), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(new_n463), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT25), .ZN(new_n740));
  NAND2_X1  g315(.A1(G103), .A2(G2104), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(G2105), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n463), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n461), .A2(G139), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n737), .B1(new_n745), .B2(new_n711), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(G2072), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n711), .A2(G26), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT28), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n461), .A2(G140), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n475), .A2(G128), .ZN(new_n751));
  OR2_X1    g326(.A1(G104), .A2(G2105), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n752), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n750), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n749), .B1(new_n755), .B2(new_n711), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2067), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n747), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n726), .A2(new_n731), .A3(new_n735), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(G160), .A2(G29), .ZN(new_n760));
  INV_X1    g335(.A(G34), .ZN(new_n761));
  AOI21_X1  g336(.A(G29), .B1(new_n761), .B2(KEYINPUT24), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(KEYINPUT24), .B2(new_n761), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G2084), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n711), .A2(G35), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G162), .B2(new_n711), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT29), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n765), .B1(G2090), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT30), .B(G28), .ZN(new_n770));
  OR2_X1    g345(.A1(KEYINPUT31), .A2(G11), .ZN(new_n771));
  NAND2_X1  g346(.A1(KEYINPUT31), .A2(G11), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n770), .A2(new_n711), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n647), .B2(new_n711), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n729), .B2(new_n730), .ZN(new_n775));
  NOR2_X1   g350(.A1(G16), .A2(G19), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n546), .B2(G16), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(G1341), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n727), .A2(G5), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G171), .B2(new_n727), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n780), .A2(G1961), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n777), .A2(G1341), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n775), .A2(new_n778), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n759), .A2(new_n769), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(G299), .A2(G16), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n727), .A2(G20), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT23), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(G1956), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n768), .A2(G2090), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n790), .A2(KEYINPUT96), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n727), .A2(G4), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n623), .B2(new_n727), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT91), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT90), .B(G1348), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT89), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n795), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n780), .A2(G1961), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT95), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n724), .B2(new_n725), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n799), .A2(new_n800), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n784), .A2(new_n792), .A3(new_n798), .A4(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(KEYINPUT96), .B1(new_n790), .B2(new_n791), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n593), .A2(G651), .ZN(new_n809));
  AND4_X1   g384(.A1(new_n809), .A2(new_n589), .A3(new_n596), .A4(new_n598), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(new_n727), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G6), .B2(new_n727), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT32), .B(G1981), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n812), .A2(new_n814), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n727), .A2(G22), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G166), .B2(new_n727), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(G1971), .Z(new_n819));
  NAND3_X1  g394(.A1(new_n815), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n586), .A2(new_n587), .ZN(new_n821));
  INV_X1    g396(.A(G74), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n498), .B1(new_n530), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(KEYINPUT87), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT87), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n585), .A2(new_n825), .A3(new_n586), .A4(new_n587), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n827), .A2(new_n727), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n727), .B2(G23), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT33), .B(G1976), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n829), .B(new_n830), .Z(new_n831));
  AOI21_X1  g406(.A(new_n820), .B1(new_n831), .B2(KEYINPUT88), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n829), .B(new_n830), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT88), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(KEYINPUT34), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT34), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n832), .A2(new_n838), .A3(new_n835), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n711), .A2(G25), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n461), .A2(G131), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n475), .A2(G119), .ZN(new_n842));
  OR2_X1    g417(.A1(G95), .A2(G2105), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n843), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n841), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n840), .B1(new_n846), .B2(new_n711), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT35), .B(G1991), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(G290), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n850), .A2(new_n727), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(new_n727), .B2(G24), .ZN(new_n852));
  INV_X1    g427(.A(G1986), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n849), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(new_n853), .B2(new_n852), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n837), .A2(new_n839), .A3(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n856), .A2(KEYINPUT36), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(KEYINPUT36), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n808), .B1(new_n857), .B2(new_n858), .ZN(G311));
  INV_X1    g434(.A(new_n858), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n856), .A2(KEYINPUT36), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n807), .B1(new_n860), .B2(new_n861), .ZN(G150));
  NAND3_X1  g437(.A1(new_n504), .A2(new_n508), .A3(G67), .ZN(new_n863));
  NAND2_X1  g438(.A1(G80), .A2(G543), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n498), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n504), .A2(new_n508), .A3(G93), .A4(new_n514), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n516), .A2(G55), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT98), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(KEYINPUT98), .B1(new_n865), .B2(new_n868), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(G860), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(KEYINPUT37), .Z(new_n876));
  NAND2_X1  g451(.A1(new_n623), .A2(G559), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n545), .A2(G651), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n879), .A2(new_n539), .A3(new_n541), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n871), .A2(new_n880), .A3(new_n872), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT97), .ZN(new_n882));
  NOR3_X1   g457(.A1(new_n880), .A2(new_n882), .A3(new_n869), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n863), .A2(new_n864), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(G651), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n866), .A2(new_n867), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT97), .B1(new_n546), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n881), .B1(new_n883), .B2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n878), .B(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n890), .A2(KEYINPUT39), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT99), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n893));
  AOI21_X1  g468(.A(G860), .B1(new_n890), .B2(KEYINPUT39), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n893), .B1(new_n892), .B2(new_n894), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n876), .B1(new_n895), .B2(new_n896), .ZN(G145));
  XNOR2_X1  g472(.A(new_n745), .B(KEYINPUT102), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n723), .A2(new_n754), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n496), .A2(KEYINPUT101), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n487), .A2(new_n495), .A3(new_n901), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n721), .A2(new_n722), .A3(new_n755), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n899), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n904), .B1(new_n899), .B2(new_n905), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n898), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n899), .A2(new_n905), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n903), .ZN(new_n911));
  AOI21_X1  g486(.A(KEYINPUT102), .B1(new_n739), .B2(new_n744), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(new_n912), .A3(new_n906), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n475), .A2(G130), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n463), .A2(G118), .ZN(new_n915));
  OAI21_X1  g490(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n917), .B1(G142), .B2(new_n461), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(new_n638), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(new_n846), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n909), .A2(new_n913), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT103), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n909), .A2(new_n913), .ZN(new_n923));
  INV_X1    g498(.A(new_n920), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n909), .A2(new_n913), .A3(new_n926), .A4(new_n920), .ZN(new_n927));
  XNOR2_X1  g502(.A(G160), .B(new_n647), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(G162), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n922), .A2(new_n925), .A3(new_n927), .A4(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n921), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n920), .B1(new_n909), .B2(new_n913), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G37), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n931), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(new_n511), .B2(new_n518), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n511), .A2(new_n518), .A3(new_n938), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n810), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(G166), .A2(KEYINPUT104), .ZN(new_n943));
  NAND3_X1  g518(.A1(G305), .A2(new_n939), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n824), .A2(new_n826), .ZN(new_n946));
  NAND2_X1  g521(.A1(G290), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n601), .A2(KEYINPUT80), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n605), .A2(new_n606), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n949), .A3(G651), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n950), .A2(new_n600), .A3(new_n824), .A4(new_n826), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n947), .A2(new_n951), .A3(KEYINPUT105), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n945), .A2(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n945), .A2(new_n952), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n947), .A2(new_n951), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n953), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT42), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n889), .B(new_n632), .Z(new_n960));
  NAND2_X1  g535(.A1(new_n615), .A2(new_n622), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(new_n567), .B2(new_n576), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT77), .B1(new_n554), .B2(new_n566), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n571), .A2(new_n575), .A3(new_n568), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n963), .A2(new_n964), .A3(new_n622), .A4(new_n615), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n960), .A2(new_n966), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n962), .A2(new_n965), .A3(KEYINPUT41), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT41), .B1(new_n962), .B2(new_n965), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n967), .B1(new_n970), .B2(new_n960), .ZN(new_n971));
  OR2_X1    g546(.A1(new_n971), .A2(KEYINPUT106), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(KEYINPUT106), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n959), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n973), .A2(new_n959), .ZN(new_n975));
  OAI21_X1  g550(.A(G868), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(G868), .B2(new_n873), .ZN(G295));
  OAI21_X1  g552(.A(new_n976), .B1(G868), .B2(new_n873), .ZN(G331));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n979));
  NAND3_X1  g554(.A1(G168), .A2(new_n533), .A3(new_n536), .ZN(new_n980));
  NAND2_X1  g555(.A1(G301), .A2(G286), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n889), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT107), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n882), .B1(new_n880), .B2(new_n869), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n546), .A2(new_n887), .A3(KEYINPUT97), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n988), .A2(new_n881), .A3(new_n982), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n889), .A2(new_n983), .A3(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n985), .A2(new_n966), .A3(new_n989), .A4(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n989), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n982), .B1(new_n988), .B2(new_n881), .ZN(new_n994));
  OAI22_X1  g569(.A1(new_n968), .A2(new_n969), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n992), .A2(new_n958), .A3(new_n995), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n996), .A2(new_n935), .ZN(new_n997));
  INV_X1    g572(.A(new_n958), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n991), .A2(new_n989), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n970), .B1(new_n985), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n984), .A2(new_n966), .A3(new_n989), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT108), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n984), .A2(new_n966), .A3(new_n1003), .A4(new_n989), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n998), .B1(new_n1000), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n997), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n992), .A2(new_n995), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n998), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1009), .A2(new_n1010), .A3(new_n935), .A4(new_n996), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n1007), .A2(KEYINPUT43), .B1(new_n1011), .B2(KEYINPUT110), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1011), .A2(KEYINPUT110), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n979), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n997), .A2(new_n1006), .A3(new_n1010), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT109), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n996), .A2(new_n935), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n958), .B1(new_n992), .B2(new_n995), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT43), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1016), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1017), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1014), .B1(new_n1022), .B2(new_n979), .ZN(G397));
  INV_X1    g598(.A(KEYINPUT45), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(new_n904), .B2(G1384), .ZN(new_n1025));
  AOI22_X1  g600(.A1(new_n461), .A2(G137), .B1(G101), .B2(new_n464), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n469), .A2(new_n470), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1026), .B(G40), .C1(new_n1027), .C2(new_n463), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(new_n853), .A3(new_n850), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1029), .A2(G1986), .A3(G290), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1032), .B(KEYINPUT111), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n723), .B(G1996), .ZN(new_n1034));
  INV_X1    g609(.A(G2067), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n754), .B(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1038));
  OR2_X1    g613(.A1(new_n846), .A2(new_n848), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n846), .A2(new_n848), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1033), .B1(new_n1029), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT125), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT123), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n1045));
  NOR2_X1   g620(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1046));
  INV_X1    g621(.A(new_n486), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n485), .B1(new_n636), .B2(new_n482), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n492), .A2(new_n494), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n636), .A2(G126), .A3(G2105), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1046), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G40), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n466), .A2(new_n471), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n1056));
  AOI21_X1  g631(.A(G1384), .B1(new_n487), .B2(new_n495), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1053), .B(new_n1055), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT115), .B1(new_n1058), .B2(G2084), .ZN(new_n1059));
  INV_X1    g634(.A(G1384), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n496), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(new_n1024), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1055), .B1(new_n1057), .B2(KEYINPUT45), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n730), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1028), .B1(new_n496), .B2(new_n1046), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1061), .A2(KEYINPUT50), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n1067));
  INV_X1    g642(.A(G2084), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1059), .A2(new_n1064), .A3(new_n1069), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1045), .B(G8), .C1(new_n1070), .C2(G286), .ZN(new_n1071));
  INV_X1    g646(.A(G8), .ZN(new_n1072));
  NOR2_X1   g647(.A1(G168), .A2(new_n1072), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1070), .A2(KEYINPUT122), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT122), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1071), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1073), .B1(new_n1070), .B2(G8), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1077), .A2(KEYINPUT51), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1044), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1070), .A2(KEYINPUT122), .A3(new_n1073), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1077), .A2(KEYINPUT51), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1084), .A2(KEYINPUT123), .A3(new_n1085), .A4(new_n1071), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1079), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1043), .B1(new_n1087), .B2(KEYINPUT62), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n1089));
  AOI211_X1 g664(.A(KEYINPUT125), .B(new_n1089), .C1(new_n1079), .C2(new_n1086), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1079), .A2(new_n1089), .A3(new_n1086), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1028), .B1(new_n1061), .B2(new_n1024), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n900), .A2(KEYINPUT45), .A3(new_n1060), .A4(new_n902), .ZN(new_n1093));
  AOI21_X1  g668(.A(G1971), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1058), .A2(G2090), .ZN(new_n1095));
  OAI21_X1  g670(.A(G8), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n582), .A2(G8), .A3(new_n583), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT55), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n582), .A2(new_n583), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1096), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1103), .B(G8), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n824), .A2(G1976), .A3(new_n826), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1072), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1106));
  INV_X1    g681(.A(G1976), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT52), .B1(G288), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1106), .ZN(new_n1111));
  INV_X1    g686(.A(G1981), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n594), .A2(new_n1112), .A3(new_n596), .A4(new_n598), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n520), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n589), .B(new_n595), .C1(new_n1114), .C2(new_n498), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(G1981), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT49), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1111), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1113), .A2(new_n1116), .A3(KEYINPUT49), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1110), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT112), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT112), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1105), .A2(new_n1124), .A3(new_n1106), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(KEYINPUT52), .A3(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1102), .A2(new_n1104), .A3(new_n1121), .A4(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(new_n1120), .A3(new_n1106), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1126), .A2(new_n1131), .A3(new_n1109), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1132), .A2(KEYINPUT124), .A3(new_n1104), .A4(new_n1102), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1092), .A2(new_n1093), .A3(new_n734), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT53), .ZN(new_n1135));
  INV_X1    g710(.A(G1961), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1134), .A2(new_n1135), .B1(new_n1136), .B2(new_n1058), .ZN(new_n1137));
  OR4_X1    g712(.A1(new_n1135), .A2(new_n1062), .A3(new_n1063), .A4(G2078), .ZN(new_n1138));
  AOI21_X1  g713(.A(G301), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1129), .A2(new_n1133), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1091), .A2(new_n1140), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1088), .A2(new_n1090), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1132), .A2(new_n1102), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT116), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1132), .A2(KEYINPUT116), .A3(new_n1102), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1104), .A2(KEYINPUT63), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1070), .A2(G8), .A3(G168), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1145), .A2(new_n1146), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1151), .B1(new_n1127), .B2(new_n1148), .ZN(new_n1152));
  INV_X1    g727(.A(G288), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1131), .A2(new_n1107), .A3(new_n1153), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1113), .B(KEYINPUT113), .Z(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n1106), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1121), .A2(new_n1126), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1157), .B(KEYINPUT114), .C1(new_n1104), .C2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT114), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1158), .A2(new_n1104), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1111), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1150), .A2(new_n1152), .B1(new_n1159), .B2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g739(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n1165));
  NOR2_X1   g740(.A1(new_n556), .A2(new_n560), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1165), .B1(new_n554), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n571), .A2(new_n575), .A3(KEYINPUT57), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(KEYINPUT56), .B(G2072), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1092), .A2(new_n1093), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1058), .A2(new_n789), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1169), .B1(new_n1173), .B2(KEYINPUT119), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1174), .B1(KEYINPUT119), .B2(new_n1173), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1061), .A2(new_n1028), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1058), .A2(new_n796), .B1(new_n1176), .B2(new_n1035), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(KEYINPUT118), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT118), .ZN(new_n1179));
  INV_X1    g754(.A(new_n796), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1180), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1061), .A2(G2067), .A3(new_n1028), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1179), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1178), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(new_n623), .ZN(new_n1186));
  AND3_X1   g761(.A1(new_n1171), .A2(new_n1169), .A3(new_n1172), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1175), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT60), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1189), .B1(new_n1178), .B2(new_n1183), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(KEYINPUT121), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1184), .A2(KEYINPUT60), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT121), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n961), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NOR3_X1   g769(.A1(new_n1190), .A2(KEYINPUT121), .A3(new_n623), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1191), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1185), .A2(new_n1189), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(G1996), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1092), .A2(new_n1093), .A3(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g775(.A(KEYINPUT58), .B(G1341), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1200), .B1(new_n1176), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1202), .A2(new_n546), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT59), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n1205));
  AOI22_X1  g780(.A1(new_n1203), .A2(new_n1204), .B1(new_n1187), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1206), .B1(new_n1204), .B2(new_n1203), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1169), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1208));
  OR2_X1    g783(.A1(new_n1208), .A2(KEYINPUT120), .ZN(new_n1209));
  AOI21_X1  g784(.A(KEYINPUT61), .B1(new_n1208), .B2(KEYINPUT120), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1187), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1207), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1188), .B1(new_n1198), .B2(new_n1212), .ZN(new_n1213));
  AND2_X1   g788(.A1(new_n1129), .A2(new_n1133), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1215));
  XNOR2_X1  g790(.A(G301), .B(KEYINPUT54), .ZN(new_n1216));
  AND4_X1   g791(.A1(KEYINPUT53), .A2(new_n1093), .A3(new_n734), .A4(new_n1055), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1216), .B1(new_n1025), .B2(new_n1217), .ZN(new_n1218));
  AOI22_X1  g793(.A1(new_n1215), .A2(new_n1216), .B1(new_n1218), .B2(new_n1137), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1087), .A2(new_n1214), .A3(new_n1219), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1164), .B1(new_n1213), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1042), .B1(new_n1142), .B2(new_n1221), .ZN(new_n1222));
  XOR2_X1   g797(.A(new_n1030), .B(KEYINPUT48), .Z(new_n1223));
  NAND2_X1  g798(.A1(new_n1041), .A2(new_n1029), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1223), .B1(new_n1224), .B2(KEYINPUT126), .ZN(new_n1225));
  OAI21_X1  g800(.A(new_n1225), .B1(KEYINPUT126), .B2(new_n1224), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1029), .A2(new_n1199), .ZN(new_n1227));
  OR2_X1    g802(.A1(new_n1227), .A2(KEYINPUT46), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1227), .A2(KEYINPUT46), .ZN(new_n1229));
  NAND3_X1  g804(.A1(new_n721), .A2(new_n722), .A3(new_n1036), .ZN(new_n1230));
  AOI22_X1  g805(.A1(new_n1228), .A2(new_n1229), .B1(new_n1029), .B2(new_n1230), .ZN(new_n1231));
  XOR2_X1   g806(.A(new_n1231), .B(KEYINPUT47), .Z(new_n1232));
  NOR3_X1   g807(.A1(new_n1034), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1233));
  NOR2_X1   g808(.A1(new_n754), .A2(G2067), .ZN(new_n1234));
  OAI21_X1  g809(.A(new_n1029), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g810(.A1(new_n1226), .A2(new_n1232), .A3(new_n1235), .ZN(new_n1236));
  INV_X1    g811(.A(new_n1236), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1222), .A2(new_n1237), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g813(.A1(new_n681), .A2(new_n457), .ZN(new_n1240));
  XNOR2_X1  g814(.A(new_n1240), .B(KEYINPUT127), .ZN(new_n1241));
  OAI21_X1  g815(.A(new_n1241), .B1(new_n708), .B2(new_n709), .ZN(new_n1242));
  AOI21_X1  g816(.A(new_n1242), .B1(new_n667), .B2(new_n668), .ZN(new_n1243));
  OAI211_X1 g817(.A(new_n1243), .B(new_n936), .C1(new_n1021), .C2(new_n1017), .ZN(G225));
  INV_X1    g818(.A(G225), .ZN(G308));
endmodule


