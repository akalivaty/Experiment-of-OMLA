//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961;
  INV_X1    g000(.A(KEYINPUT102), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(KEYINPUT22), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n208), .B(new_n203), .C1(KEYINPUT22), .C2(new_n206), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(KEYINPUT77), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT77), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n207), .A2(new_n213), .A3(new_n209), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT25), .ZN(new_n216));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(KEYINPUT68), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n216), .B1(new_n218), .B2(KEYINPUT23), .ZN(new_n219));
  INV_X1    g018(.A(G169gat), .ZN(new_n220));
  INV_X1    g019(.A(G176gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT67), .B1(new_n217), .B2(KEYINPUT23), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n229));
  INV_X1    g028(.A(G183gat), .ZN(new_n230));
  INV_X1    g029(.A(G190gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n231), .ZN(new_n233));
  NAND3_X1  g032(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT69), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n232), .A2(KEYINPUT69), .A3(new_n233), .A4(new_n234), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n219), .A2(new_n228), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n234), .B(KEYINPUT65), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(new_n230), .A3(new_n231), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n232), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n217), .A2(KEYINPUT23), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n225), .A2(new_n227), .A3(new_n247), .A4(new_n226), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n240), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n239), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n222), .A2(KEYINPUT26), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n222), .B(KEYINPUT68), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n226), .B(new_n251), .C1(new_n252), .C2(KEYINPUT26), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT27), .B(G183gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(new_n231), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT28), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT70), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n255), .A2(new_n257), .B1(G183gat), .B2(G190gat), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n253), .B(new_n258), .C1(new_n255), .C2(new_n257), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n250), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G226gat), .ZN(new_n261));
  INV_X1    g060(.A(G233gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(KEYINPUT29), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n265), .B1(new_n250), .B2(new_n259), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n215), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT78), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n250), .B(new_n259), .C1(new_n261), .C2(new_n262), .ZN(new_n269));
  INV_X1    g068(.A(new_n215), .ZN(new_n270));
  INV_X1    g069(.A(new_n260), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n269), .B(new_n270), .C1(new_n271), .C2(new_n265), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n267), .A2(new_n268), .A3(new_n272), .ZN(new_n273));
  OAI211_X1 g072(.A(KEYINPUT78), .B(new_n215), .C1(new_n264), .C2(new_n266), .ZN(new_n274));
  XNOR2_X1  g073(.A(G8gat), .B(G36gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(G64gat), .B(G92gat), .ZN(new_n276));
  XOR2_X1   g075(.A(new_n275), .B(new_n276), .Z(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n273), .A2(new_n274), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n278), .B1(new_n273), .B2(new_n274), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(KEYINPUT30), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT79), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n273), .A2(new_n274), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(new_n277), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT30), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n280), .A2(KEYINPUT79), .A3(KEYINPUT30), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n281), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G155gat), .ZN(new_n289));
  INV_X1    g088(.A(G162gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT2), .ZN(new_n292));
  NOR2_X1   g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G141gat), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT81), .B1(new_n295), .B2(G148gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT81), .ZN(new_n297));
  INV_X1    g096(.A(G148gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(new_n298), .A3(G141gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT80), .B(G141gat), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n296), .B(new_n299), .C1(new_n300), .C2(new_n298), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT82), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n296), .A2(new_n299), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT82), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n303), .B(new_n304), .C1(new_n298), .C2(new_n300), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n294), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(G141gat), .B(G148gat), .Z(new_n307));
  AND2_X1   g106(.A1(new_n307), .A2(new_n292), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n308), .A2(new_n291), .A3(new_n293), .ZN(new_n309));
  XOR2_X1   g108(.A(KEYINPUT83), .B(KEYINPUT3), .Z(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NOR3_X1   g110(.A1(new_n306), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G127gat), .B(G134gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT71), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n314), .B1(new_n315), .B2(KEYINPUT1), .ZN(new_n316));
  XNOR2_X1  g115(.A(G113gat), .B(G120gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(KEYINPUT1), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320));
  INV_X1    g119(.A(G113gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n321), .A2(G120gat), .ZN(new_n322));
  INV_X1    g121(.A(G120gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(G113gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n320), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  OR2_X1    g124(.A1(G127gat), .A2(G134gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(G127gat), .A2(G134gat), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n326), .A2(new_n327), .B1(KEYINPUT71), .B2(new_n320), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n319), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT3), .B1(new_n306), .B2(new_n309), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n313), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n306), .A2(new_n309), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n330), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT4), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G225gat), .A2(G233gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT72), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n330), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n319), .A2(KEYINPUT72), .A3(new_n329), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n334), .A2(KEYINPUT4), .A3(new_n342), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n333), .A2(new_n337), .A3(new_n338), .A4(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT5), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n331), .B1(new_n306), .B2(new_n309), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n335), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n338), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n345), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n309), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n302), .A2(new_n305), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n351), .B1(new_n352), .B2(new_n294), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n330), .B1(new_n353), .B2(KEYINPUT3), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n348), .B1(new_n354), .B2(new_n313), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT4), .B1(new_n334), .B2(new_n342), .ZN(new_n356));
  NOR4_X1   g155(.A1(new_n306), .A2(new_n331), .A3(new_n309), .A4(new_n336), .ZN(new_n357));
  NOR3_X1   g156(.A1(new_n356), .A2(new_n357), .A3(KEYINPUT5), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n350), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G1gat), .B(G29gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT0), .ZN(new_n362));
  XNOR2_X1  g161(.A(G57gat), .B(G85gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n360), .A2(KEYINPUT6), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT6), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n344), .A2(new_n349), .B1(new_n358), .B2(new_n355), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n367), .B1(new_n368), .B2(new_n364), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n350), .A2(new_n359), .A3(new_n364), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n366), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n288), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n260), .A2(KEYINPUT73), .A3(new_n342), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n319), .A2(KEYINPUT72), .A3(new_n329), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT72), .B1(new_n319), .B2(new_n329), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT73), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT73), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n340), .A2(new_n377), .A3(new_n341), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n376), .A2(new_n378), .A3(new_n250), .A4(new_n259), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n373), .A2(new_n379), .A3(G227gat), .A4(G233gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT32), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT33), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(G15gat), .B(G43gat), .Z(new_n384));
  XNOR2_X1  g183(.A(G71gat), .B(G99gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n381), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n386), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n380), .B(KEYINPUT32), .C1(new_n382), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n379), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT34), .ZN(new_n392));
  NAND2_X1  g191(.A1(G227gat), .A2(G233gat), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n392), .B1(new_n391), .B2(new_n393), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n390), .A2(KEYINPUT74), .A3(new_n396), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n387), .B(new_n389), .C1(new_n395), .C2(new_n394), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n396), .A2(KEYINPUT74), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(G228gat), .A2(G233gat), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n215), .B1(new_n312), .B2(KEYINPUT29), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT29), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n210), .A2(KEYINPUT84), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n211), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n210), .A2(KEYINPUT84), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n404), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n334), .B1(new_n408), .B2(new_n310), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n401), .B1(new_n403), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(new_n215), .B2(KEYINPUT29), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n401), .B1(new_n412), .B2(new_n353), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n413), .A2(new_n402), .A3(KEYINPUT85), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT85), .B1(new_n413), .B2(new_n402), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n410), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G78gat), .B(G106gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT31), .B(G50gat), .ZN(new_n418));
  XOR2_X1   g217(.A(new_n417), .B(new_n418), .Z(new_n419));
  NAND2_X1  g218(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT86), .B(G22gat), .ZN(new_n421));
  INV_X1    g220(.A(new_n419), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n410), .B(new_n422), .C1(new_n414), .C2(new_n415), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n421), .B1(new_n420), .B2(new_n423), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n400), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT35), .B1(new_n372), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n371), .A2(KEYINPUT90), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT90), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n366), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n424), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n433), .A2(new_n425), .A3(KEYINPUT35), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n390), .A2(new_n396), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n398), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n432), .A2(new_n434), .A3(new_n288), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n428), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n278), .A2(KEYINPUT37), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n279), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n267), .A2(new_n272), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT38), .B1(new_n441), .B2(KEYINPUT37), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT89), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n440), .A2(KEYINPUT89), .A3(new_n442), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT37), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n440), .B1(new_n448), .B2(new_n283), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n280), .B1(new_n449), .B2(KEYINPUT38), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n447), .A2(new_n450), .A3(new_n429), .A4(new_n431), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n433), .A2(new_n425), .ZN(new_n452));
  INV_X1    g251(.A(new_n281), .ZN(new_n453));
  INV_X1    g252(.A(new_n287), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT79), .B1(new_n280), .B2(KEYINPUT30), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT40), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT87), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n356), .A2(new_n357), .ZN(new_n459));
  AOI211_X1 g258(.A(KEYINPUT39), .B(new_n338), .C1(new_n459), .C2(new_n333), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n458), .B1(new_n460), .B2(new_n365), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n338), .B1(new_n459), .B2(new_n333), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT39), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n464), .A2(KEYINPUT87), .A3(new_n364), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n335), .A2(new_n338), .A3(new_n346), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n467), .A2(KEYINPUT88), .A3(KEYINPUT39), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT88), .B1(new_n467), .B2(KEYINPUT39), .ZN(new_n469));
  NOR3_X1   g268(.A1(new_n462), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n457), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n364), .B1(new_n350), .B2(new_n359), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n461), .B2(new_n465), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n472), .B1(new_n473), .B2(KEYINPUT40), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n456), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n451), .A2(new_n452), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n400), .A2(KEYINPUT36), .ZN(new_n477));
  XOR2_X1   g276(.A(KEYINPUT75), .B(KEYINPUT36), .Z(new_n478));
  OAI21_X1  g277(.A(KEYINPUT76), .B1(new_n436), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT76), .ZN(new_n480));
  INV_X1    g279(.A(new_n478), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n435), .A2(new_n480), .A3(new_n398), .A4(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n477), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n452), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n372), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n438), .B1(new_n476), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G43gat), .B(G50gat), .ZN(new_n490));
  INV_X1    g289(.A(G29gat), .ZN(new_n491));
  INV_X1    g290(.A(G36gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT14), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT14), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n494), .B1(G29gat), .B2(G36gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(G29gat), .A2(G36gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(KEYINPUT15), .B(new_n490), .C1(new_n496), .C2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT92), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n496), .B(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n498), .B1(new_n490), .B2(KEYINPUT15), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n502), .B1(KEYINPUT15), .B2(new_n490), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT17), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(G15gat), .B(G22gat), .Z(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT93), .ZN(new_n508));
  INV_X1    g307(.A(G1gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT16), .ZN(new_n510));
  XNOR2_X1  g309(.A(G15gat), .B(G22gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT93), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n508), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(G1gat), .B1(new_n508), .B2(new_n513), .ZN(new_n515));
  OAI21_X1  g314(.A(G8gat), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n508), .A2(new_n513), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n509), .ZN(new_n518));
  INV_X1    g317(.A(G8gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT16), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n508), .B(new_n513), .C1(new_n520), .C2(G1gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n499), .B(KEYINPUT17), .C1(new_n501), .C2(new_n503), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n506), .A2(new_n516), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(G229gat), .A2(G233gat), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n514), .A2(new_n515), .A3(G8gat), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n519), .B1(new_n518), .B2(new_n521), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n504), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n524), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n489), .B1(new_n529), .B2(KEYINPUT94), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT94), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n524), .A2(new_n528), .A3(new_n531), .A4(new_n525), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n524), .A2(new_n528), .A3(KEYINPUT18), .A4(new_n525), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n525), .B(KEYINPUT13), .Z(new_n535));
  NOR3_X1   g334(.A1(new_n526), .A2(new_n527), .A3(new_n504), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n501), .A2(new_n503), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n516), .A2(new_n522), .B1(new_n537), .B2(new_n499), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n535), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n533), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT91), .ZN(new_n543));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544));
  INV_X1    g343(.A(G197gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT11), .B(G169gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT12), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n542), .A2(new_n543), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n549), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n540), .B1(new_n530), .B2(new_n532), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n551), .B1(new_n552), .B2(KEYINPUT91), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n487), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g355(.A1(G71gat), .A2(G78gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(G71gat), .A2(G78gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G57gat), .B(G64gat), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G57gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(G64gat), .ZN(new_n564));
  INV_X1    g363(.A(G64gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(G57gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G71gat), .B(G78gat), .ZN(new_n568));
  INV_X1    g367(.A(new_n561), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n562), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT21), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(G127gat), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n516), .B(new_n522), .C1(new_n572), .C2(new_n571), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G183gat), .B(G211gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT96), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(new_n289), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n580), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n578), .A2(new_n584), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT8), .ZN(new_n590));
  NAND2_X1  g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT7), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(G85gat), .ZN(new_n594));
  INV_X1    g393(.A(G92gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n590), .A2(new_n593), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G99gat), .B(G106gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  AND3_X1   g400(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI22_X1  g403(.A1(KEYINPUT8), .A2(new_n589), .B1(new_n594), .B2(new_n595), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(new_n599), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n506), .A2(new_n523), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n598), .A2(new_n600), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n599), .B1(new_n604), .B2(new_n605), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AND2_X1   g410(.A1(G232gat), .A2(G233gat), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n504), .A2(new_n611), .B1(KEYINPUT41), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G190gat), .B(G218gat), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT97), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n612), .A2(KEYINPUT41), .ZN(new_n619));
  XNOR2_X1  g418(.A(G134gat), .B(G162gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n614), .A2(new_n616), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n618), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n621), .B1(new_n618), .B2(new_n622), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n588), .A2(new_n627), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n562), .B(new_n570), .C1(new_n609), .C2(new_n610), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n571), .A2(new_n606), .A3(new_n601), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G230gat), .A2(G233gat), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT100), .ZN(new_n634));
  XNOR2_X1  g433(.A(G120gat), .B(G148gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(G176gat), .B(G204gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT10), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n562), .A2(new_n570), .A3(KEYINPUT10), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n611), .A2(new_n642), .A3(KEYINPUT98), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT98), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n562), .A2(new_n570), .A3(KEYINPUT10), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n644), .B1(new_n607), .B2(new_n645), .ZN(new_n646));
  AOI22_X1  g445(.A1(new_n641), .A2(new_n631), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n632), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n640), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n631), .A2(new_n641), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n643), .A2(new_n646), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n652), .A2(KEYINPUT99), .A3(new_n632), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n632), .B(KEYINPUT101), .Z(new_n656));
  NOR2_X1   g455(.A1(new_n647), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n638), .B1(new_n634), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n628), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n202), .B1(new_n556), .B2(new_n661), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n435), .A2(new_n481), .A3(new_n398), .ZN(new_n663));
  AOI22_X1  g462(.A1(new_n663), .A2(new_n480), .B1(new_n400), .B2(KEYINPUT36), .ZN(new_n664));
  AOI22_X1  g463(.A1(new_n664), .A2(new_n479), .B1(new_n484), .B2(new_n372), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n451), .A2(new_n475), .A3(new_n452), .ZN(new_n666));
  AOI22_X1  g465(.A1(new_n665), .A2(new_n666), .B1(new_n428), .B2(new_n437), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(new_n554), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n668), .A2(KEYINPUT102), .A3(new_n660), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n662), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n368), .A2(new_n367), .A3(new_n364), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n472), .A2(KEYINPUT6), .ZN(new_n672));
  INV_X1    g471(.A(new_n370), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g475(.A(KEYINPUT16), .B(G8gat), .Z(new_n677));
  NAND3_X1  g476(.A1(new_n670), .A2(new_n456), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n288), .B1(new_n662), .B2(new_n669), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n519), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT42), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(G1325gat));
  INV_X1    g483(.A(G15gat), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n685), .A3(new_n436), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n483), .B1(new_n662), .B2(new_n669), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n686), .B1(new_n685), .B2(new_n687), .ZN(G1326gat));
  NAND2_X1  g487(.A1(new_n670), .A2(new_n484), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT43), .B(G22gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  NOR3_X1   g490(.A1(new_n588), .A2(new_n627), .A3(new_n659), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n668), .A2(new_n491), .A3(new_n674), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT45), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n695), .B1(new_n667), .B2(new_n627), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n487), .A2(KEYINPUT44), .A3(new_n626), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n659), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n555), .A2(new_n587), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT103), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n702), .A2(new_n674), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n694), .B1(new_n703), .B2(new_n491), .ZN(G1328gat));
  NAND4_X1  g503(.A1(new_n668), .A2(new_n492), .A3(new_n456), .A4(new_n692), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT46), .Z(new_n706));
  AND2_X1   g505(.A1(new_n702), .A2(new_n456), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(new_n707), .B2(new_n492), .ZN(G1329gat));
  INV_X1    g507(.A(new_n483), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n696), .A2(new_n697), .A3(new_n709), .A4(new_n701), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(G43gat), .ZN(new_n711));
  INV_X1    g510(.A(G43gat), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n668), .A2(new_n712), .A3(new_n436), .A4(new_n692), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT47), .B1(new_n713), .B2(KEYINPUT104), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1330gat));
  NAND4_X1  g515(.A1(new_n696), .A2(new_n697), .A3(new_n484), .A4(new_n701), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G50gat), .ZN(new_n718));
  INV_X1    g517(.A(G50gat), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n668), .A2(new_n719), .A3(new_n484), .A4(new_n692), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT48), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n721), .B(new_n723), .ZN(G1331gat));
  NOR3_X1   g523(.A1(new_n628), .A2(new_n555), .A3(new_n699), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n487), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n371), .B(KEYINPUT106), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g528(.A(new_n288), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n731), .A2(KEYINPUT107), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(KEYINPUT107), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1333gat));
  NAND2_X1  g535(.A1(new_n726), .A2(new_n436), .ZN(new_n737));
  INV_X1    g536(.A(G71gat), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n726), .A2(G71gat), .A3(new_n709), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n739), .B(new_n740), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n741), .B(new_n742), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n740), .B1(new_n747), .B2(new_n739), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n746), .A2(new_n748), .ZN(G1334gat));
  NAND2_X1  g548(.A1(new_n726), .A2(new_n484), .ZN(new_n750));
  XNOR2_X1  g549(.A(KEYINPUT110), .B(G78gat), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1335gat));
  NAND2_X1  g551(.A1(new_n554), .A2(new_n587), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT111), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n754), .A2(new_n659), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n698), .A2(new_n674), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G85gat), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n756), .A2(new_n757), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n667), .B2(new_n627), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n487), .A2(KEYINPUT113), .A3(new_n626), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n762), .A2(new_n763), .A3(new_n754), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n762), .A2(new_n763), .A3(KEYINPUT51), .A4(new_n754), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n674), .A2(new_n594), .A3(new_n659), .ZN(new_n769));
  OAI22_X1  g568(.A1(new_n759), .A2(new_n760), .B1(new_n768), .B2(new_n769), .ZN(G1336gat));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n696), .A2(new_n697), .A3(new_n456), .A4(new_n755), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G92gat), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n288), .A2(G92gat), .A3(new_n699), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n771), .B(new_n773), .C1(new_n768), .C2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(new_n766), .B2(new_n767), .ZN(new_n777));
  INV_X1    g576(.A(new_n773), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT52), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n779), .ZN(G1337gat));
  INV_X1    g579(.A(G99gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n436), .A2(new_n781), .A3(new_n659), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n698), .A2(new_n709), .A3(new_n755), .ZN(new_n783));
  OAI22_X1  g582(.A1(new_n768), .A2(new_n782), .B1(new_n783), .B2(new_n781), .ZN(G1338gat));
  XOR2_X1   g583(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n785));
  NAND4_X1  g584(.A1(new_n696), .A2(new_n697), .A3(new_n484), .A4(new_n755), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n786), .B2(G106gat), .ZN(new_n787));
  OR3_X1    g586(.A1(new_n452), .A2(G106gat), .A3(new_n699), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n768), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n788), .B1(new_n766), .B2(new_n767), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n786), .A2(new_n791), .A3(G106gat), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n791), .B1(new_n786), .B2(G106gat), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n790), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n789), .B1(new_n794), .B2(new_n795), .ZN(G1339gat));
  NOR3_X1   g595(.A1(new_n536), .A2(new_n538), .A3(new_n535), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n525), .B1(new_n524), .B2(new_n528), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n548), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n659), .B(new_n799), .C1(new_n542), .C2(new_n551), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n657), .A2(new_n801), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n802), .A2(KEYINPUT55), .A3(new_n638), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n801), .B1(new_n647), .B2(new_n656), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT99), .B1(new_n652), .B2(new_n632), .ZN(new_n806));
  AOI211_X1 g605(.A(new_n640), .B(new_n648), .C1(new_n650), .C2(new_n651), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n804), .B(new_n805), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n804), .B1(new_n654), .B2(new_n805), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n803), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n802), .A2(new_n638), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT116), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n812), .B1(new_n814), .B2(new_n808), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n655), .B(new_n811), .C1(new_n815), .C2(KEYINPUT55), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n800), .B1(new_n816), .B2(new_n554), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT117), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n819), .B(new_n800), .C1(new_n816), .C2(new_n554), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(new_n627), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n799), .B1(new_n542), .B2(new_n551), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n816), .A2(new_n627), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n588), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n660), .A2(new_n554), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT118), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n626), .B1(new_n817), .B2(KEYINPUT117), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n823), .B1(new_n830), .B2(new_n820), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n829), .B(new_n826), .C1(new_n831), .C2(new_n588), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n456), .A2(new_n371), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n833), .A2(new_n436), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n828), .A2(new_n452), .A3(new_n832), .A4(new_n834), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n835), .A2(new_n321), .A3(new_n554), .ZN(new_n836));
  INV_X1    g635(.A(new_n427), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n828), .A2(new_n837), .A3(new_n727), .A4(new_n832), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(new_n288), .A3(new_n555), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n836), .B1(new_n840), .B2(new_n321), .ZN(G1340gat));
  NAND2_X1  g640(.A1(new_n659), .A2(new_n323), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT119), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n839), .A2(new_n288), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(G120gat), .B1(new_n835), .B2(new_n699), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT120), .ZN(G1341gat));
  OAI21_X1  g646(.A(G127gat), .B1(new_n835), .B2(new_n587), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n839), .A2(new_n288), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n587), .A2(G127gat), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(G1342gat));
  NOR3_X1   g650(.A1(new_n456), .A2(G134gat), .A3(new_n627), .ZN(new_n852));
  XOR2_X1   g651(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n853));
  NAND3_X1  g652(.A1(new_n839), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n853), .ZN(new_n855));
  INV_X1    g654(.A(new_n852), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n838), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(G134gat), .B1(new_n835), .B2(new_n627), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n854), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT122), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n859), .B(new_n860), .ZN(G1343gat));
  AND2_X1   g660(.A1(new_n828), .A2(new_n832), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT124), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n709), .A2(new_n452), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n862), .A2(new_n863), .A3(new_n727), .A4(new_n864), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n456), .A2(G141gat), .A3(new_n554), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n828), .A2(new_n727), .A3(new_n832), .A4(new_n864), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT124), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT125), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n865), .A2(new_n871), .A3(new_n866), .A4(new_n868), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n828), .A2(new_n873), .A3(new_n484), .A4(new_n832), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n483), .A2(new_n833), .ZN(new_n875));
  XOR2_X1   g674(.A(KEYINPUT123), .B(KEYINPUT55), .Z(new_n876));
  OAI211_X1 g675(.A(new_n655), .B(new_n811), .C1(new_n815), .C2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n800), .B1(new_n877), .B2(new_n554), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n627), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n588), .B1(new_n879), .B2(new_n824), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n484), .B1(new_n827), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n875), .B1(new_n881), .B2(KEYINPUT57), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n874), .A2(new_n555), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT58), .B1(new_n883), .B2(new_n300), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n870), .A2(new_n872), .A3(new_n884), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n883), .A2(new_n300), .ZN(new_n886));
  NOR4_X1   g685(.A1(new_n867), .A2(G141gat), .A3(new_n456), .A4(new_n554), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT58), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n885), .A2(new_n888), .ZN(G1344gat));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n882), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n890), .B(G148gat), .C1(new_n891), .C2(new_n699), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n828), .A2(KEYINPUT57), .A3(new_n484), .A4(new_n832), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n881), .A2(new_n873), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n875), .A2(new_n699), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n298), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n892), .B1(new_n897), .B2(new_n890), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n865), .A2(new_n288), .A3(new_n868), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n659), .A2(new_n298), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(G1345gat));
  OAI21_X1  g700(.A(G155gat), .B1(new_n891), .B2(new_n587), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n588), .A2(new_n289), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n899), .B2(new_n903), .ZN(G1346gat));
  OAI21_X1  g703(.A(G162gat), .B1(new_n891), .B2(new_n627), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n626), .A2(new_n290), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n905), .B1(new_n899), .B2(new_n906), .ZN(G1347gat));
  NOR2_X1   g706(.A1(new_n727), .A2(new_n288), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n436), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT126), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n862), .A2(new_n452), .A3(new_n910), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(new_n220), .A3(new_n554), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n862), .A2(new_n371), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n427), .A2(new_n288), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n555), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n912), .B1(new_n917), .B2(new_n220), .ZN(G1348gat));
  OAI21_X1  g717(.A(G176gat), .B1(new_n911), .B2(new_n699), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n659), .A2(new_n221), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n919), .B1(new_n915), .B2(new_n920), .ZN(G1349gat));
  NAND2_X1  g720(.A1(new_n588), .A2(new_n254), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n913), .A2(new_n914), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(G183gat), .B1(new_n911), .B2(new_n587), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT60), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT60), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n924), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(G1350gat));
  OAI21_X1  g729(.A(G190gat), .B1(new_n911), .B2(new_n627), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT61), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n933), .B(G190gat), .C1(new_n911), .C2(new_n627), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n916), .A2(new_n231), .A3(new_n626), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1351gat));
  NAND2_X1  g736(.A1(new_n908), .A2(new_n483), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n938), .B1(new_n893), .B2(new_n894), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n940), .A2(new_n545), .A3(new_n554), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n709), .A2(new_n452), .A3(new_n288), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n913), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n555), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n941), .B1(new_n945), .B2(new_n545), .ZN(G1352gat));
  XOR2_X1   g745(.A(KEYINPUT127), .B(G204gat), .Z(new_n947));
  NAND2_X1  g746(.A1(new_n659), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(KEYINPUT62), .B1(new_n943), .B2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT62), .ZN(new_n950));
  INV_X1    g749(.A(new_n948), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n913), .A2(new_n950), .A3(new_n942), .A4(new_n951), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n940), .A2(new_n699), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n949), .B(new_n952), .C1(new_n953), .C2(new_n947), .ZN(G1353gat));
  NAND3_X1  g753(.A1(new_n944), .A2(new_n204), .A3(new_n588), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n588), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  OAI21_X1  g758(.A(G218gat), .B1(new_n940), .B2(new_n627), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n626), .A2(new_n205), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n960), .B1(new_n943), .B2(new_n961), .ZN(G1355gat));
endmodule


