

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582;

  XNOR2_X1 U323 ( .A(G1GAT), .B(KEYINPUT71), .ZN(n415) );
  AND2_X1 U324 ( .A1(n421), .A2(n459), .ZN(n422) );
  XNOR2_X1 U325 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U326 ( .A(n389), .B(n388), .ZN(n391) );
  XNOR2_X1 U327 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U328 ( .A(n373), .B(n360), .ZN(n558) );
  XOR2_X1 U329 ( .A(KEYINPUT64), .B(KEYINPUT78), .Z(n291) );
  XOR2_X1 U330 ( .A(n355), .B(n354), .Z(n292) );
  AND2_X1 U331 ( .A1(n567), .A2(n551), .ZN(n402) );
  NOR2_X1 U332 ( .A1(n425), .A2(n430), .ZN(n431) );
  XNOR2_X1 U333 ( .A(n387), .B(n386), .ZN(n388) );
  NOR2_X1 U334 ( .A1(n558), .A2(n423), .ZN(n424) );
  XOR2_X1 U335 ( .A(G57GAT), .B(KEYINPUT13), .Z(n395) );
  INV_X1 U336 ( .A(n396), .ZN(n397) );
  XOR2_X1 U337 ( .A(KEYINPUT73), .B(n395), .Z(n409) );
  XNOR2_X1 U338 ( .A(n409), .B(n397), .ZN(n398) );
  XNOR2_X1 U339 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U340 ( .A(n399), .B(n398), .ZN(n425) );
  XNOR2_X1 U341 ( .A(n379), .B(n378), .ZN(n504) );
  XNOR2_X1 U342 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n457) );
  XNOR2_X1 U343 ( .A(G211GAT), .B(G218GAT), .ZN(n293) );
  XNOR2_X1 U344 ( .A(n293), .B(KEYINPUT21), .ZN(n294) );
  XOR2_X1 U345 ( .A(n294), .B(KEYINPUT86), .Z(n296) );
  XNOR2_X1 U346 ( .A(G197GAT), .B(G204GAT), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n341) );
  XOR2_X1 U348 ( .A(KEYINPUT85), .B(KEYINPUT88), .Z(n298) );
  XNOR2_X1 U349 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n341), .B(n299), .ZN(n309) );
  XNOR2_X1 U352 ( .A(G106GAT), .B(G78GAT), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n300), .B(G148GAT), .ZN(n396) );
  XOR2_X1 U354 ( .A(G50GAT), .B(G162GAT), .Z(n356) );
  XOR2_X1 U355 ( .A(n396), .B(n356), .Z(n307) );
  XOR2_X1 U356 ( .A(G141GAT), .B(G22GAT), .Z(n363) );
  XOR2_X1 U357 ( .A(G155GAT), .B(KEYINPUT87), .Z(n302) );
  XNOR2_X1 U358 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n301) );
  XNOR2_X1 U359 ( .A(n302), .B(n301), .ZN(n321) );
  XOR2_X1 U360 ( .A(n321), .B(KEYINPUT23), .Z(n304) );
  NAND2_X1 U361 ( .A1(G228GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U362 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U363 ( .A(n363), .B(n305), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U365 ( .A(n309), .B(n308), .ZN(n465) );
  XOR2_X1 U366 ( .A(G57GAT), .B(KEYINPUT6), .Z(n311) );
  XNOR2_X1 U367 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n310) );
  XNOR2_X1 U368 ( .A(n311), .B(n310), .ZN(n329) );
  XOR2_X1 U369 ( .A(KEYINPUT78), .B(G127GAT), .Z(n313) );
  XNOR2_X1 U370 ( .A(G29GAT), .B(G134GAT), .ZN(n312) );
  XNOR2_X1 U371 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U372 ( .A(KEYINPUT89), .B(G148GAT), .Z(n315) );
  XNOR2_X1 U373 ( .A(G141GAT), .B(G120GAT), .ZN(n314) );
  XNOR2_X1 U374 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U375 ( .A(n317), .B(n316), .Z(n323) );
  XOR2_X1 U376 ( .A(G85GAT), .B(G162GAT), .Z(n319) );
  NAND2_X1 U377 ( .A1(G225GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U378 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U381 ( .A(n324), .B(KEYINPUT4), .Z(n327) );
  XNOR2_X1 U382 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n325), .B(KEYINPUT82), .ZN(n448) );
  XNOR2_X1 U384 ( .A(n448), .B(KEYINPUT5), .ZN(n326) );
  XNOR2_X1 U385 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n471) );
  INV_X1 U387 ( .A(n471), .ZN(n518) );
  XOR2_X1 U388 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n331) );
  XNOR2_X1 U389 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n330) );
  XNOR2_X1 U390 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U391 ( .A(n332), .B(G183GAT), .Z(n334) );
  XNOR2_X1 U392 ( .A(G169GAT), .B(G176GAT), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n449) );
  XOR2_X1 U394 ( .A(G92GAT), .B(G64GAT), .Z(n380) );
  XOR2_X1 U395 ( .A(KEYINPUT93), .B(n380), .Z(n336) );
  NAND2_X1 U396 ( .A1(G226GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U397 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U398 ( .A(G8GAT), .B(KEYINPUT79), .Z(n412) );
  XOR2_X1 U399 ( .A(n337), .B(n412), .Z(n343) );
  XOR2_X1 U400 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n339) );
  XNOR2_X1 U401 ( .A(G36GAT), .B(KEYINPUT90), .ZN(n338) );
  XNOR2_X1 U402 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U403 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U405 ( .A(n449), .B(n344), .Z(n520) );
  XOR2_X1 U406 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n346) );
  XNOR2_X1 U407 ( .A(G36GAT), .B(G29GAT), .ZN(n345) );
  XNOR2_X1 U408 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U409 ( .A(KEYINPUT70), .B(n347), .Z(n373) );
  XOR2_X1 U410 ( .A(G85GAT), .B(KEYINPUT75), .Z(n381) );
  XOR2_X1 U411 ( .A(G92GAT), .B(G99GAT), .Z(n349) );
  NAND2_X1 U412 ( .A1(G232GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U413 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U414 ( .A(n381), .B(n350), .ZN(n359) );
  XOR2_X1 U415 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n352) );
  XNOR2_X1 U416 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n351) );
  XNOR2_X1 U417 ( .A(n352), .B(n351), .ZN(n355) );
  XNOR2_X1 U418 ( .A(G190GAT), .B(G106GAT), .ZN(n353) );
  XNOR2_X1 U419 ( .A(n291), .B(n353), .ZN(n354) );
  XOR2_X1 U420 ( .A(G43GAT), .B(G134GAT), .Z(n443) );
  XNOR2_X1 U421 ( .A(n443), .B(n356), .ZN(n357) );
  XNOR2_X1 U422 ( .A(n292), .B(n357), .ZN(n358) );
  XNOR2_X1 U423 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U424 ( .A(KEYINPUT68), .B(KEYINPUT66), .Z(n362) );
  XNOR2_X1 U425 ( .A(KEYINPUT67), .B(KEYINPUT30), .ZN(n361) );
  XNOR2_X1 U426 ( .A(n362), .B(n361), .ZN(n367) );
  XOR2_X1 U427 ( .A(G43GAT), .B(G50GAT), .Z(n365) );
  XOR2_X1 U428 ( .A(n363), .B(n415), .Z(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U430 ( .A(n367), .B(n366), .Z(n369) );
  NAND2_X1 U431 ( .A1(G229GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n369), .B(n368), .ZN(n379) );
  XOR2_X1 U433 ( .A(KEYINPUT72), .B(KEYINPUT29), .Z(n371) );
  XNOR2_X1 U434 ( .A(G8GAT), .B(KEYINPUT69), .ZN(n370) );
  XNOR2_X1 U435 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U436 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U437 ( .A(G197GAT), .B(G113GAT), .Z(n375) );
  XNOR2_X1 U438 ( .A(G169GAT), .B(G15GAT), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n376) );
  INV_X1 U440 ( .A(n504), .ZN(n567) );
  INV_X1 U441 ( .A(KEYINPUT41), .ZN(n400) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n383) );
  XOR2_X1 U443 ( .A(G176GAT), .B(G204GAT), .Z(n382) );
  XNOR2_X1 U444 ( .A(n383), .B(n382), .ZN(n389) );
  XOR2_X1 U445 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n385) );
  XNOR2_X1 U446 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n385), .B(n384), .ZN(n387) );
  AND2_X1 U448 ( .A1(G230GAT), .A2(G233GAT), .ZN(n386) );
  INV_X1 U449 ( .A(KEYINPUT33), .ZN(n390) );
  XNOR2_X1 U450 ( .A(n391), .B(n390), .ZN(n394) );
  XNOR2_X1 U451 ( .A(G99GAT), .B(G71GAT), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n392), .B(G120GAT), .ZN(n446) );
  XNOR2_X1 U453 ( .A(n446), .B(KEYINPUT74), .ZN(n393) );
  XNOR2_X1 U454 ( .A(n394), .B(n393), .ZN(n399) );
  XNOR2_X1 U455 ( .A(n400), .B(n425), .ZN(n551) );
  INV_X1 U456 ( .A(KEYINPUT46), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n402), .B(n401), .ZN(n421) );
  XOR2_X1 U458 ( .A(G78GAT), .B(G155GAT), .Z(n404) );
  XNOR2_X1 U459 ( .A(G22GAT), .B(G211GAT), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U461 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n406) );
  XNOR2_X1 U462 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n420) );
  XOR2_X1 U465 ( .A(n409), .B(KEYINPUT80), .Z(n411) );
  NAND2_X1 U466 ( .A1(G231GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U467 ( .A(n411), .B(n410), .ZN(n418) );
  XOR2_X1 U468 ( .A(G15GAT), .B(G127GAT), .Z(n440) );
  XOR2_X1 U469 ( .A(n412), .B(n440), .Z(n414) );
  XNOR2_X1 U470 ( .A(G183GAT), .B(G71GAT), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n414), .B(n413), .ZN(n416) );
  XOR2_X1 U472 ( .A(n420), .B(n419), .Z(n459) );
  XOR2_X1 U473 ( .A(n422), .B(KEYINPUT110), .Z(n423) );
  XNOR2_X1 U474 ( .A(n424), .B(KEYINPUT47), .ZN(n435) );
  XOR2_X1 U475 ( .A(KEYINPUT45), .B(KEYINPUT111), .Z(n426) );
  XNOR2_X1 U476 ( .A(KEYINPUT65), .B(n426), .ZN(n429) );
  INV_X1 U477 ( .A(n459), .ZN(n574) );
  XNOR2_X1 U478 ( .A(KEYINPUT36), .B(KEYINPUT98), .ZN(n427) );
  XNOR2_X1 U479 ( .A(n427), .B(n558), .ZN(n577) );
  NAND2_X1 U480 ( .A1(n574), .A2(n577), .ZN(n428) );
  XOR2_X1 U481 ( .A(n429), .B(n428), .Z(n430) );
  XOR2_X1 U482 ( .A(KEYINPUT112), .B(n431), .Z(n432) );
  NOR2_X1 U483 ( .A1(n567), .A2(n432), .ZN(n433) );
  XNOR2_X1 U484 ( .A(KEYINPUT113), .B(n433), .ZN(n434) );
  NAND2_X1 U485 ( .A1(n435), .A2(n434), .ZN(n436) );
  XNOR2_X1 U486 ( .A(n436), .B(KEYINPUT48), .ZN(n546) );
  AND2_X1 U487 ( .A1(n520), .A2(n546), .ZN(n437) );
  XOR2_X1 U488 ( .A(n437), .B(KEYINPUT54), .Z(n438) );
  NOR2_X1 U489 ( .A1(n518), .A2(n438), .ZN(n566) );
  NAND2_X1 U490 ( .A1(n465), .A2(n566), .ZN(n439) );
  XNOR2_X1 U491 ( .A(n439), .B(KEYINPUT55), .ZN(n452) );
  XNOR2_X1 U492 ( .A(n440), .B(KEYINPUT20), .ZN(n441) );
  XNOR2_X1 U493 ( .A(n441), .B(KEYINPUT83), .ZN(n442) );
  XOR2_X1 U494 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U495 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U496 ( .A(n445), .B(n444), .ZN(n447) );
  XOR2_X1 U497 ( .A(n447), .B(n446), .Z(n451) );
  XNOR2_X1 U498 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U499 ( .A(n451), .B(n450), .ZN(n530) );
  NAND2_X1 U500 ( .A1(n452), .A2(n530), .ZN(n453) );
  XNOR2_X2 U501 ( .A(n453), .B(KEYINPUT121), .ZN(n562) );
  NAND2_X1 U502 ( .A1(n562), .A2(n551), .ZN(n456) );
  XOR2_X1 U503 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n454) );
  XNOR2_X1 U504 ( .A(n454), .B(G176GAT), .ZN(n455) );
  XNOR2_X1 U505 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  NAND2_X1 U506 ( .A1(n558), .A2(n562), .ZN(n458) );
  XNOR2_X1 U507 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XNOR2_X1 U508 ( .A(KEYINPUT96), .B(KEYINPUT34), .ZN(n480) );
  XOR2_X1 U509 ( .A(G1GAT), .B(KEYINPUT97), .Z(n478) );
  OR2_X1 U510 ( .A1(n504), .A2(n425), .ZN(n490) );
  NOR2_X1 U511 ( .A1(n459), .A2(n558), .ZN(n460) );
  XOR2_X1 U512 ( .A(KEYINPUT81), .B(n460), .Z(n461) );
  XNOR2_X1 U513 ( .A(n461), .B(KEYINPUT16), .ZN(n475) );
  XOR2_X1 U514 ( .A(n465), .B(KEYINPUT28), .Z(n525) );
  XNOR2_X1 U515 ( .A(KEYINPUT27), .B(n520), .ZN(n464) );
  NAND2_X1 U516 ( .A1(n518), .A2(n464), .ZN(n548) );
  NOR2_X1 U517 ( .A1(n525), .A2(n548), .ZN(n529) );
  XOR2_X1 U518 ( .A(n530), .B(KEYINPUT84), .Z(n462) );
  NAND2_X1 U519 ( .A1(n529), .A2(n462), .ZN(n474) );
  NOR2_X1 U520 ( .A1(n465), .A2(n530), .ZN(n463) );
  XNOR2_X1 U521 ( .A(n463), .B(KEYINPUT26), .ZN(n565) );
  NAND2_X1 U522 ( .A1(n464), .A2(n565), .ZN(n470) );
  NAND2_X1 U523 ( .A1(n520), .A2(n530), .ZN(n466) );
  NAND2_X1 U524 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U525 ( .A(n467), .B(KEYINPUT94), .ZN(n468) );
  XOR2_X1 U526 ( .A(KEYINPUT25), .B(n468), .Z(n469) );
  NAND2_X1 U527 ( .A1(n470), .A2(n469), .ZN(n472) );
  NAND2_X1 U528 ( .A1(n472), .A2(n471), .ZN(n473) );
  NAND2_X1 U529 ( .A1(n474), .A2(n473), .ZN(n486) );
  NAND2_X1 U530 ( .A1(n475), .A2(n486), .ZN(n505) );
  NOR2_X1 U531 ( .A1(n490), .A2(n505), .ZN(n476) );
  XOR2_X1 U532 ( .A(KEYINPUT95), .B(n476), .Z(n484) );
  NAND2_X1 U533 ( .A1(n484), .A2(n518), .ZN(n477) );
  XNOR2_X1 U534 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U535 ( .A(n480), .B(n479), .ZN(G1324GAT) );
  NAND2_X1 U536 ( .A1(n484), .A2(n520), .ZN(n481) );
  XNOR2_X1 U537 ( .A(n481), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U538 ( .A(G15GAT), .B(KEYINPUT35), .Z(n483) );
  NAND2_X1 U539 ( .A1(n484), .A2(n530), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n483), .B(n482), .ZN(G1326GAT) );
  NAND2_X1 U541 ( .A1(n484), .A2(n525), .ZN(n485) );
  XNOR2_X1 U542 ( .A(n485), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U543 ( .A(G29GAT), .B(KEYINPUT39), .Z(n493) );
  NAND2_X1 U544 ( .A1(n577), .A2(n486), .ZN(n487) );
  NOR2_X1 U545 ( .A1(n574), .A2(n487), .ZN(n488) );
  XOR2_X1 U546 ( .A(n488), .B(KEYINPUT37), .Z(n489) );
  XNOR2_X1 U547 ( .A(KEYINPUT99), .B(n489), .ZN(n517) );
  NOR2_X1 U548 ( .A1(n490), .A2(n517), .ZN(n491) );
  XNOR2_X1 U549 ( .A(n491), .B(KEYINPUT38), .ZN(n498) );
  NAND2_X1 U550 ( .A1(n518), .A2(n498), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NAND2_X1 U552 ( .A1(n498), .A2(n520), .ZN(n494) );
  XNOR2_X1 U553 ( .A(n494), .B(KEYINPUT100), .ZN(n495) );
  XNOR2_X1 U554 ( .A(G36GAT), .B(n495), .ZN(G1329GAT) );
  NAND2_X1 U555 ( .A1(n498), .A2(n530), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n496), .B(KEYINPUT40), .ZN(n497) );
  XNOR2_X1 U557 ( .A(G43GAT), .B(n497), .ZN(G1330GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n500) );
  NAND2_X1 U559 ( .A1(n525), .A2(n498), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U561 ( .A(G50GAT), .B(n501), .ZN(G1331GAT) );
  XNOR2_X1 U562 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n502), .B(KEYINPUT104), .ZN(n503) );
  XOR2_X1 U564 ( .A(KEYINPUT103), .B(n503), .Z(n507) );
  NAND2_X1 U565 ( .A1(n504), .A2(n551), .ZN(n516) );
  NOR2_X1 U566 ( .A1(n505), .A2(n516), .ZN(n512) );
  NAND2_X1 U567 ( .A1(n512), .A2(n518), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n507), .B(n506), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n512), .A2(n520), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n508), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U571 ( .A1(n512), .A2(n530), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n509), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n511) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(n515) );
  NAND2_X1 U576 ( .A1(n512), .A2(n525), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n513), .B(KEYINPUT105), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n515), .B(n514), .ZN(G1335GAT) );
  NOR2_X1 U579 ( .A1(n517), .A2(n516), .ZN(n526) );
  NAND2_X1 U580 ( .A1(n518), .A2(n526), .ZN(n519) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(n519), .ZN(G1336GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n522) );
  NAND2_X1 U583 ( .A1(n526), .A2(n520), .ZN(n521) );
  XNOR2_X1 U584 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(n523), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n526), .A2(n530), .ZN(n524) );
  XNOR2_X1 U587 ( .A(n524), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U588 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U589 ( .A(n527), .B(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  INV_X1 U591 ( .A(n546), .ZN(n532) );
  NAND2_X1 U592 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U593 ( .A1(n532), .A2(n531), .ZN(n541) );
  NAND2_X1 U594 ( .A1(n567), .A2(n541), .ZN(n533) );
  XNOR2_X1 U595 ( .A(G113GAT), .B(n533), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n535) );
  NAND2_X1 U597 ( .A1(n541), .A2(n551), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(n536), .ZN(G1341GAT) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(KEYINPUT116), .ZN(n540) );
  XOR2_X1 U601 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n538) );
  NAND2_X1 U602 ( .A1(n541), .A2(n574), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U606 ( .A1(n541), .A2(n558), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(n545) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT118), .Z(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  XOR2_X1 U610 ( .A(G141GAT), .B(KEYINPUT119), .Z(n550) );
  NAND2_X1 U611 ( .A1(n546), .A2(n565), .ZN(n547) );
  NOR2_X1 U612 ( .A1(n548), .A2(n547), .ZN(n557) );
  NAND2_X1 U613 ( .A1(n557), .A2(n567), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(G1344GAT) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n555) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n553) );
  NAND2_X1 U617 ( .A1(n557), .A2(n551), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n574), .A2(n557), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n556), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U623 ( .A(n559), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n561) );
  NAND2_X1 U625 ( .A1(n567), .A2(n562), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(G1348GAT) );
  XOR2_X1 U627 ( .A(G183GAT), .B(KEYINPUT123), .Z(n564) );
  NAND2_X1 U628 ( .A1(n562), .A2(n574), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(G1350GAT) );
  AND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n578) );
  NAND2_X1 U631 ( .A1(n578), .A2(n567), .ZN(n570) );
  XOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT60), .Z(n568) );
  XNOR2_X1 U633 ( .A(KEYINPUT59), .B(n568), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U636 ( .A1(n578), .A2(n425), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(n573), .ZN(G1353GAT) );
  XOR2_X1 U639 ( .A(G211GAT), .B(KEYINPUT125), .Z(n576) );
  NAND2_X1 U640 ( .A1(n578), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1354GAT) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n582) );
  XOR2_X1 U643 ( .A(KEYINPUT127), .B(KEYINPUT126), .Z(n580) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(G1355GAT) );
endmodule

