//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1186, new_n1187, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1237, new_n1238;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT64), .Z(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT65), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n209), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT66), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n223), .A2(new_n207), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  OAI22_X1  g0026(.A1(new_n220), .A2(KEYINPUT1), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NOR3_X1   g0027(.A1(new_n213), .A2(new_n222), .A3(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT67), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n232), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NAND3_X1  g0044(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n223), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n206), .A2(G20), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n249), .A2(G50), .A3(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n207), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n248), .ZN(new_n260));
  OAI221_X1 g0060(.A(new_n251), .B1(G50), .B2(new_n245), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  XOR2_X1   g0061(.A(new_n261), .B(KEYINPUT9), .Z(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G223), .ZN(new_n268));
  INV_X1    g0068(.A(G77), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G222), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n266), .ZN(new_n272));
  OAI221_X1 g0072(.A(new_n268), .B1(new_n269), .B2(new_n270), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT68), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(KEYINPUT68), .A2(G33), .A3(G41), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n223), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(KEYINPUT69), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT69), .ZN(new_n285));
  AOI211_X1 g0085(.A(new_n285), .B(new_n223), .C1(new_n281), .C2(new_n282), .ZN(new_n286));
  OAI211_X1 g0086(.A(G274), .B(new_n278), .C1(new_n284), .C2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G226), .ZN(new_n288));
  INV_X1    g0088(.A(new_n278), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n289), .B1(new_n284), .B2(new_n286), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n275), .B(new_n287), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT70), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n291), .B(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n262), .B1(new_n293), .B2(G190), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT74), .ZN(new_n295));
  AOI21_X1  g0095(.A(KEYINPUT10), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n293), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G200), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n294), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n298), .B(new_n294), .C1(new_n295), .C2(KEYINPUT10), .ZN(new_n301));
  AND2_X1   g0101(.A1(KEYINPUT71), .A2(G179), .ZN(new_n302));
  NOR2_X1   g0102(.A1(KEYINPUT71), .A2(G179), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n297), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n293), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n261), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n300), .A2(new_n301), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G13), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(G1), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G68), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G20), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  XOR2_X1   g0115(.A(new_n315), .B(KEYINPUT12), .Z(new_n316));
  INV_X1    g0116(.A(G33), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n207), .A2(new_n317), .ZN(new_n318));
  OAI221_X1 g0118(.A(new_n314), .B1(new_n254), .B2(new_n269), .C1(new_n202), .C2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(KEYINPUT11), .A3(new_n248), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n249), .A2(G68), .A3(new_n250), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n316), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT11), .B1(new_n319), .B2(new_n248), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT79), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  OAI211_X1 g0126(.A(G226), .B(new_n266), .C1(new_n263), .C2(new_n264), .ZN(new_n327));
  OAI211_X1 g0127(.A(G232), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G33), .A2(G97), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n274), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT75), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT75), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n330), .A2(new_n333), .A3(new_n274), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G274), .ZN(new_n336));
  INV_X1    g0136(.A(new_n223), .ZN(new_n337));
  INV_X1    g0137(.A(new_n282), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT68), .B1(G33), .B2(G41), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n285), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n283), .A2(KEYINPUT69), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n336), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n343), .A2(KEYINPUT76), .A3(new_n278), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT76), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n287), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n335), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G238), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT77), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n290), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n341), .A2(new_n342), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n351), .A2(KEYINPUT77), .A3(new_n289), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n348), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT13), .B1(new_n347), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT77), .B1(new_n351), .B2(new_n289), .ZN(new_n355));
  AOI211_X1 g0155(.A(new_n349), .B(new_n278), .C1(new_n341), .C2(new_n342), .ZN(new_n356));
  OAI21_X1  g0156(.A(G238), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT13), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n332), .A2(new_n334), .B1(new_n287), .B2(new_n345), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .A4(new_n344), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n354), .A2(new_n360), .A3(G179), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT78), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(KEYINPUT14), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n354), .A2(new_n360), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(G169), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n363), .A2(KEYINPUT14), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n362), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n306), .B1(new_n354), .B2(new_n360), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n367), .B1(new_n370), .B2(new_n364), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n326), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n324), .ZN(new_n373));
  INV_X1    g0173(.A(G200), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n365), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G190), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n354), .A2(new_n360), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n373), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT16), .ZN(new_n380));
  INV_X1    g0180(.A(G58), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n381), .A2(new_n313), .ZN(new_n382));
  OAI21_X1  g0182(.A(G20), .B1(new_n382), .B2(new_n201), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT80), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n257), .A2(new_n384), .A3(G159), .ZN(new_n385));
  INV_X1    g0185(.A(G159), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT80), .B1(new_n318), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n383), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT81), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n380), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n270), .B2(G20), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n313), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n390), .B1(new_n394), .B2(new_n388), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n392), .A2(new_n393), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G68), .ZN(new_n397));
  INV_X1    g0197(.A(new_n388), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n397), .A2(new_n389), .A3(new_n380), .A4(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n248), .ZN(new_n401));
  INV_X1    g0201(.A(new_n249), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n253), .A2(new_n250), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n402), .A2(new_n403), .B1(new_n245), .B2(new_n253), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n270), .A2(G223), .A3(new_n266), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G33), .A2(G87), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n270), .A2(G1698), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n407), .B(new_n408), .C1(new_n409), .C2(new_n288), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n274), .ZN(new_n411));
  OAI211_X1 g0211(.A(G232), .B(new_n289), .C1(new_n284), .C2(new_n286), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n287), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n306), .ZN(new_n414));
  INV_X1    g0214(.A(new_n304), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n406), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT18), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n413), .A2(new_n374), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(G190), .B2(new_n413), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n404), .B1(new_n400), .B2(new_n248), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT82), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n420), .A2(new_n421), .A3(KEYINPUT82), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(KEYINPUT17), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT17), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n420), .A2(new_n421), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT83), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n424), .A2(KEYINPUT83), .A3(KEYINPUT17), .A4(new_n425), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n418), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n270), .A2(G232), .A3(new_n266), .ZN(new_n433));
  INV_X1    g0233(.A(G107), .ZN(new_n434));
  OAI221_X1 g0234(.A(new_n433), .B1(new_n434), .B2(new_n270), .C1(new_n409), .C2(new_n348), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n274), .ZN(new_n436));
  INV_X1    g0236(.A(G244), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n436), .B(new_n287), .C1(new_n437), .C2(new_n290), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n438), .A2(G190), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n439), .B1(new_n374), .B2(new_n438), .ZN(new_n440));
  OAI22_X1  g0240(.A1(new_n252), .A2(new_n318), .B1(new_n207), .B2(new_n269), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT15), .B(G87), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n441), .A2(KEYINPUT72), .B1(new_n255), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(KEYINPUT72), .B2(new_n441), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n248), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n245), .A2(G77), .ZN(new_n447));
  XNOR2_X1  g0247(.A(new_n447), .B(KEYINPUT73), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n269), .B1(new_n206), .B2(G20), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n448), .B1(new_n249), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n440), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n451), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n438), .A2(new_n304), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n438), .A2(G169), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n309), .A2(new_n379), .A3(new_n432), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT5), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT87), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n460), .B2(G41), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n276), .A2(KEYINPUT87), .A3(KEYINPUT5), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n277), .A2(G1), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n464), .B1(new_n341), .B2(new_n342), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G270), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n351), .A2(G274), .A3(new_n464), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n270), .A2(G257), .A3(new_n266), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n265), .A2(G303), .ZN(new_n469));
  INV_X1    g0269(.A(G264), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n468), .B(new_n469), .C1(new_n409), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n274), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n466), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(G20), .B1(new_n317), .B2(G97), .ZN(new_n474));
  NAND3_X1  g0274(.A1(KEYINPUT86), .A2(G33), .A3(G283), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT86), .B1(G33), .B2(G283), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G116), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n247), .A2(new_n223), .B1(G20), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(KEYINPUT20), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT95), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT95), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n478), .A2(new_n483), .A3(KEYINPUT20), .A4(new_n480), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n478), .A2(new_n480), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT20), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n482), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n206), .A2(new_n479), .A3(G13), .A4(G20), .ZN(new_n489));
  XNOR2_X1  g0289(.A(new_n489), .B(KEYINPUT94), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n206), .A2(G33), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n245), .A2(new_n491), .A3(new_n223), .A4(new_n247), .ZN(new_n492));
  OR3_X1    g0292(.A1(new_n492), .A2(KEYINPUT93), .A3(new_n479), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT93), .B1(new_n492), .B2(new_n479), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n473), .A2(new_n496), .A3(G169), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT96), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT21), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT21), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n497), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G179), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n473), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n496), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n500), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  OR2_X1    g0306(.A1(new_n473), .A2(G190), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n473), .A2(new_n374), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n496), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT23), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n511), .A2(new_n207), .A3(G107), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT23), .B1(new_n434), .B2(G20), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G116), .ZN(new_n514));
  OAI22_X1  g0314(.A1(new_n512), .A2(new_n513), .B1(G20), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n270), .A2(new_n207), .A3(G87), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT22), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT22), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n270), .A2(new_n518), .A3(new_n207), .A4(G87), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n515), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  OR2_X1    g0320(.A1(new_n520), .A2(KEYINPUT24), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n260), .B1(new_n520), .B2(KEYINPUT24), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n311), .A2(G20), .A3(new_n434), .ZN(new_n524));
  OR2_X1    g0324(.A1(new_n524), .A2(KEYINPUT25), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(KEYINPUT25), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n525), .B(new_n526), .C1(new_n434), .C2(new_n492), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  AOI22_X1  g0329(.A1(G264), .A2(new_n465), .B1(new_n343), .B2(new_n464), .ZN(new_n530));
  OAI211_X1 g0330(.A(G250), .B(new_n266), .C1(new_n263), .C2(new_n264), .ZN(new_n531));
  OAI211_X1 g0331(.A(G257), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n532));
  INV_X1    g0332(.A(G294), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n531), .B(new_n532), .C1(new_n317), .C2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT97), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n534), .A2(new_n535), .A3(new_n274), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n535), .B1(new_n534), .B2(new_n274), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n306), .B1(new_n530), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n465), .A2(G264), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n534), .A2(new_n274), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n467), .A3(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n542), .A2(new_n503), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n529), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n530), .A2(new_n538), .A3(new_n376), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT98), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n530), .A2(new_n538), .A3(KEYINPUT98), .A4(new_n376), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n542), .A2(new_n374), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n527), .B1(new_n521), .B2(new_n522), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n545), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n265), .A2(new_n437), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n554), .A2(KEYINPUT85), .A3(KEYINPUT4), .A4(new_n266), .ZN(new_n555));
  NAND2_X1  g0355(.A1(KEYINPUT85), .A2(KEYINPUT4), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n270), .A2(G244), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n266), .B1(KEYINPUT85), .B2(KEYINPUT4), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OR2_X1    g0359(.A1(new_n476), .A2(new_n477), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n267), .A2(G250), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n555), .A2(new_n559), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n562), .A2(new_n274), .B1(new_n343), .B2(new_n464), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n465), .A2(G257), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(G190), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT88), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT88), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n563), .A2(new_n567), .A3(G190), .A4(new_n564), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g0369(.A(KEYINPUT84), .B(KEYINPUT6), .Z(new_n570));
  INV_X1    g0370(.A(G97), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n570), .B1(new_n571), .B2(G107), .ZN(new_n572));
  XNOR2_X1  g0372(.A(G97), .B(G107), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n572), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  OAI22_X1  g0374(.A1(new_n574), .A2(new_n207), .B1(new_n269), .B2(new_n318), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n434), .B1(new_n392), .B2(new_n393), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n248), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n245), .A2(G97), .ZN(new_n578));
  INV_X1    g0378(.A(new_n492), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n578), .B1(new_n579), .B2(G97), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n563), .A2(new_n564), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n581), .B1(G200), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n563), .A2(new_n304), .A3(new_n564), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT89), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT89), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n563), .A2(new_n586), .A3(new_n304), .A4(new_n564), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n582), .A2(new_n306), .B1(new_n577), .B2(new_n580), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n569), .A2(new_n583), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n270), .A2(new_n207), .A3(G68), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT19), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n207), .B1(new_n329), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(G87), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n571), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n593), .B1(G107), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n592), .B1(new_n329), .B2(G20), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n591), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n598), .A2(new_n248), .B1(new_n246), .B2(new_n442), .ZN(new_n599));
  OAI21_X1  g0399(.A(KEYINPUT92), .B1(new_n492), .B2(new_n594), .ZN(new_n600));
  OR3_X1    g0400(.A1(new_n492), .A2(KEYINPUT92), .A3(new_n594), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  MUX2_X1   g0402(.A(G250), .B(G274), .S(new_n463), .Z(new_n603));
  NAND2_X1  g0403(.A1(new_n351), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT90), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT90), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n351), .A2(new_n606), .A3(new_n603), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  OAI221_X1 g0408(.A(new_n514), .B1(new_n272), .B2(new_n348), .C1(new_n266), .C2(new_n557), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n274), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n602), .B1(new_n611), .B2(G200), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n605), .A2(new_n607), .B1(new_n274), .B2(new_n609), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(G190), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n611), .A2(new_n306), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n579), .A2(new_n443), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n599), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT91), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n613), .A2(new_n304), .ZN(new_n620));
  OR2_X1    g0420(.A1(new_n618), .A2(KEYINPUT91), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n616), .A2(new_n619), .A3(new_n620), .A4(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n510), .A2(new_n553), .A3(new_n590), .A4(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n458), .A2(new_n624), .ZN(G372));
  NAND2_X1  g0425(.A1(new_n365), .A2(G169), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(new_n363), .A3(KEYINPUT14), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n627), .A2(new_n371), .A3(new_n361), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n325), .ZN(new_n629));
  INV_X1    g0429(.A(new_n378), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n456), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n629), .A2(new_n631), .B1(new_n431), .B2(new_n430), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT18), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n416), .A2(new_n414), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(KEYINPUT100), .A3(new_n406), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT100), .B1(new_n634), .B2(new_n406), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n633), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT100), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n417), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(new_n635), .A3(KEYINPUT18), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n301), .B(new_n300), .C1(new_n632), .C2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n644), .A2(new_n308), .ZN(new_n645));
  INV_X1    g0445(.A(new_n615), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n569), .A2(new_n583), .B1(new_n551), .B2(new_n552), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n500), .A2(new_n544), .A3(new_n502), .A4(new_n505), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n588), .A2(new_n589), .ZN(new_n650));
  AOI211_X1 g0450(.A(KEYINPUT26), .B(new_n646), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n623), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT26), .B1(new_n652), .B2(new_n650), .ZN(new_n653));
  INV_X1    g0453(.A(new_n620), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT99), .ZN(new_n655));
  AOI211_X1 g0455(.A(new_n618), .B(new_n654), .C1(new_n655), .C2(new_n616), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n611), .A2(KEYINPUT99), .A3(new_n306), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n651), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n645), .B1(new_n458), .B2(new_n660), .ZN(G369));
  OR3_X1    g0461(.A1(new_n312), .A2(KEYINPUT27), .A3(G20), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT27), .B1(new_n312), .B2(G20), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT101), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(G343), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(G343), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n496), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n506), .B2(new_n509), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n506), .B2(new_n672), .ZN(new_n674));
  INV_X1    g0474(.A(G330), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n529), .A2(new_n671), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n553), .A2(new_n677), .B1(new_n545), .B2(new_n671), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n553), .A2(new_n506), .A3(new_n670), .A4(new_n677), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n544), .B2(new_n671), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n679), .A2(new_n681), .ZN(G399));
  INV_X1    g0482(.A(new_n210), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(G41), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n595), .A2(G107), .A3(G116), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G1), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n226), .B2(new_n685), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT31), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n473), .A2(new_n304), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n691), .A2(new_n611), .A3(new_n542), .A4(new_n582), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n563), .A2(new_n564), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n465), .A2(G264), .B1(new_n274), .B2(new_n534), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n693), .A2(new_n504), .A3(new_n694), .A4(new_n613), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT30), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n692), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n563), .A2(new_n694), .A3(new_n564), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(new_n611), .ZN(new_n699));
  AOI21_X1  g0499(.A(KEYINPUT30), .B1(new_n699), .B2(new_n504), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n671), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  OAI22_X1  g0501(.A1(new_n624), .A2(new_n671), .B1(new_n690), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n690), .B2(new_n701), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n675), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n646), .A2(new_n650), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT26), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n622), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n648), .A2(KEYINPUT102), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n499), .A2(KEYINPUT21), .B1(new_n496), .B2(new_n504), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT102), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n710), .A2(new_n711), .A3(new_n502), .A4(new_n544), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n709), .A2(new_n647), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n646), .B1(new_n713), .B2(new_n650), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n708), .B1(new_n714), .B2(KEYINPUT26), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n658), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(KEYINPUT29), .A3(new_n670), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT29), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n660), .B2(new_n671), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n704), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n689), .B1(new_n720), .B2(G1), .ZN(G364));
  NOR2_X1   g0521(.A1(new_n310), .A2(G20), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G45), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n685), .A2(G1), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT103), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n674), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n223), .B1(G20), .B2(new_n306), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n374), .A2(G179), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n731), .A2(G20), .A3(G190), .ZN(new_n732));
  INV_X1    g0532(.A(G303), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G179), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G190), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G20), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI221_X1 g0537(.A(new_n265), .B1(new_n732), .B2(new_n733), .C1(new_n737), .C2(new_n533), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n376), .A2(new_n374), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n415), .A2(G20), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR4_X1   g0541(.A1(new_n304), .A2(new_n207), .A3(new_n376), .A4(G200), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n741), .A2(G326), .B1(G322), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n207), .A2(G190), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n415), .A2(G200), .A3(new_n744), .ZN(new_n745));
  XOR2_X1   g0545(.A(KEYINPUT33), .B(G317), .Z(new_n746));
  OAI21_X1  g0546(.A(new_n743), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n415), .A2(new_n374), .A3(new_n744), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI211_X1 g0549(.A(new_n738), .B(new_n747), .C1(G311), .C2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n744), .A2(new_n734), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n751), .A2(KEYINPUT108), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(KEYINPUT108), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n744), .A2(new_n731), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n755), .A2(G329), .B1(G283), .B2(new_n757), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT109), .Z(new_n759));
  NAND2_X1  g0559(.A1(new_n750), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT107), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n732), .A2(new_n594), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n761), .B1(new_n762), .B2(new_n265), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(new_n269), .B2(new_n748), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n736), .A2(G97), .ZN(new_n765));
  OAI221_X1 g0565(.A(new_n765), .B1(new_n434), .B2(new_n756), .C1(new_n740), .C2(new_n202), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n762), .A2(new_n761), .A3(new_n265), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n745), .A2(new_n313), .ZN(new_n768));
  NOR4_X1   g0568(.A1(new_n764), .A2(new_n766), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n751), .A2(new_n386), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT106), .ZN(new_n771));
  XNOR2_X1  g0571(.A(KEYINPUT105), .B(KEYINPUT32), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n771), .B(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n742), .B(KEYINPUT104), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n769), .B(new_n773), .C1(new_n381), .C2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n730), .B1(new_n760), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n727), .A2(new_n729), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n683), .A2(new_n265), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n778), .A2(G355), .B1(new_n479), .B2(new_n683), .ZN(new_n779));
  INV_X1    g0579(.A(new_n226), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G45), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(new_n240), .B2(G45), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n210), .A2(new_n265), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n779), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n776), .B1(new_n777), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n724), .B1(new_n728), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n674), .A2(new_n675), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n676), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n786), .B1(new_n788), .B2(new_n724), .ZN(G396));
  INV_X1    g0589(.A(new_n724), .ZN(new_n790));
  INV_X1    g0590(.A(new_n456), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n671), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n453), .A2(new_n670), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n452), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n792), .B1(new_n794), .B2(new_n791), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(new_n660), .B2(new_n671), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n670), .B(new_n795), .C1(new_n651), .C2(new_n659), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n790), .B1(new_n799), .B2(new_n704), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n704), .B2(new_n799), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n756), .A2(new_n313), .ZN(new_n802));
  INV_X1    g0602(.A(new_n732), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n265), .B(new_n802), .C1(G50), .C2(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n381), .B2(new_n737), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G137), .A2(new_n741), .B1(new_n749), .B2(G159), .ZN(new_n806));
  INV_X1    g0606(.A(G150), .ZN(new_n807));
  INV_X1    g0607(.A(G143), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n806), .B1(new_n807), .B2(new_n745), .C1(new_n774), .C2(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT34), .Z(new_n810));
  AOI211_X1 g0610(.A(new_n805), .B(new_n810), .C1(G132), .C2(new_n755), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n749), .A2(G116), .B1(G294), .B2(new_n742), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n733), .B2(new_n740), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n270), .B1(new_n803), .B2(G107), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n814), .B(new_n765), .C1(new_n594), .C2(new_n756), .ZN(new_n815));
  INV_X1    g0615(.A(G311), .ZN(new_n816));
  INV_X1    g0616(.A(G283), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n754), .A2(new_n816), .B1(new_n817), .B2(new_n745), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n813), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n729), .B1(new_n811), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n729), .A2(new_n725), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n724), .B1(new_n269), .B2(new_n821), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n820), .B(new_n822), .C1(new_n726), .C2(new_n795), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n801), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G384));
  INV_X1    g0625(.A(KEYINPUT35), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n479), .B(new_n225), .C1(new_n574), .C2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n826), .B2(new_n574), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT36), .Z(new_n829));
  OAI211_X1 g0629(.A(new_n780), .B(G77), .C1(new_n381), .C2(new_n313), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n202), .A2(G68), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n206), .B(G13), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n372), .A2(new_n670), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  XOR2_X1   g0635(.A(KEYINPUT111), .B(KEYINPUT38), .Z(new_n836));
  NAND2_X1  g0636(.A1(new_n406), .A2(new_n665), .ZN(new_n837));
  AND3_X1   g0637(.A1(new_n420), .A2(new_n421), .A3(KEYINPUT82), .ZN(new_n838));
  AOI21_X1  g0638(.A(KEYINPUT82), .B1(new_n420), .B2(new_n421), .ZN(new_n839));
  NOR3_X1   g0639(.A1(new_n838), .A2(new_n839), .A3(new_n427), .ZN(new_n840));
  INV_X1    g0640(.A(new_n429), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n431), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n837), .B1(new_n642), .B2(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n422), .B(new_n837), .C1(new_n636), .C2(new_n637), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n838), .A2(new_n839), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT37), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n417), .A2(new_n846), .A3(new_n837), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n844), .A2(KEYINPUT37), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n836), .B1(new_n843), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT39), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n394), .A2(new_n388), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT16), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n405), .B1(new_n852), .B2(new_n260), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n634), .B2(new_n665), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n845), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n847), .A2(new_n845), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n853), .A2(new_n665), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n858), .B(KEYINPUT38), .C1(new_n432), .C2(new_n859), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n849), .A2(new_n850), .A3(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n417), .B(new_n633), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n859), .B1(new_n842), .B2(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n855), .A2(KEYINPUT37), .B1(new_n847), .B2(new_n845), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n850), .B1(new_n866), .B2(new_n860), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n835), .B1(new_n861), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n326), .A2(new_n670), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT110), .B1(new_n629), .B2(new_n630), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT110), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n871), .B(new_n378), .C1(new_n628), .C2(new_n325), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n869), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n871), .B1(new_n372), .B2(new_n378), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n629), .A2(KEYINPUT110), .A3(new_n630), .ZN(new_n875));
  INV_X1    g0675(.A(new_n869), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n792), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n798), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n866), .A2(new_n860), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n878), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n643), .A2(new_n664), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n868), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n458), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n717), .A2(new_n885), .A3(new_n719), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n645), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n884), .B(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT113), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n695), .A2(new_n696), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n699), .A2(KEYINPUT30), .A3(new_n504), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n890), .A2(new_n891), .A3(new_n692), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n889), .B(KEYINPUT31), .C1(new_n892), .C2(new_n671), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT113), .B1(new_n701), .B2(new_n690), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n895), .A2(new_n702), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n874), .A2(new_n876), .A3(new_n875), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n876), .B1(new_n874), .B2(new_n875), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n795), .B(new_n896), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT40), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n849), .B2(new_n860), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n878), .A2(new_n795), .A3(new_n881), .A4(new_n896), .ZN(new_n903));
  XNOR2_X1  g0703(.A(KEYINPUT112), .B(KEYINPUT40), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n900), .A2(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n895), .A2(new_n702), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n458), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n905), .B(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n888), .B1(new_n908), .B2(new_n675), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n206), .B2(new_n722), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n908), .A2(new_n888), .A3(new_n675), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n833), .B1(new_n910), .B2(new_n911), .ZN(G367));
  NOR2_X1   g0712(.A1(new_n236), .A2(new_n783), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n777), .B1(new_n210), .B2(new_n442), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n202), .A2(new_n748), .B1(new_n745), .B2(new_n386), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(G150), .B2(new_n742), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n736), .A2(G68), .ZN(new_n917));
  INV_X1    g0717(.A(G137), .ZN(new_n918));
  OAI221_X1 g0718(.A(new_n917), .B1(new_n381), .B2(new_n732), .C1(new_n918), .C2(new_n751), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n265), .B1(new_n757), .B2(G77), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n920), .A2(KEYINPUT116), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n741), .A2(G143), .B1(new_n920), .B2(KEYINPUT116), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n916), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n757), .A2(G97), .ZN(new_n925));
  INV_X1    g0725(.A(G317), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n925), .B(new_n265), .C1(new_n926), .C2(new_n751), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(G107), .B2(new_n736), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT115), .B1(new_n803), .B2(G116), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT46), .ZN(new_n930));
  INV_X1    g0730(.A(new_n745), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(G294), .ZN(new_n932));
  AOI22_X1  g0732(.A1(G283), .A2(new_n749), .B1(new_n741), .B2(G311), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n928), .A2(new_n930), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n774), .A2(new_n733), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n924), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT47), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n729), .B1(new_n936), .B2(new_n937), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n790), .B1(new_n913), .B2(new_n914), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT117), .ZN(new_n941));
  INV_X1    g0741(.A(new_n658), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n942), .A2(new_n646), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n671), .A2(new_n602), .ZN(new_n944));
  MUX2_X1   g0744(.A(new_n942), .B(new_n943), .S(new_n944), .Z(new_n945));
  INV_X1    g0745(.A(new_n727), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n941), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n723), .A2(G1), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n581), .A2(new_n671), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n590), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n650), .A2(new_n670), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(new_n681), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT45), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n953), .A2(new_n681), .ZN(new_n956));
  XOR2_X1   g0756(.A(KEYINPUT114), .B(KEYINPUT44), .Z(new_n957));
  XNOR2_X1  g0757(.A(new_n956), .B(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n679), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n506), .A2(new_n670), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n678), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n680), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(new_n676), .Z(new_n965));
  NAND3_X1  g0765(.A1(new_n961), .A2(new_n720), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n720), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n684), .B(KEYINPUT41), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n948), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NOR3_X1   g0769(.A1(new_n680), .A2(new_n950), .A3(KEYINPUT42), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n650), .B1(new_n950), .B2(new_n544), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n970), .B1(new_n971), .B2(new_n670), .ZN(new_n972));
  OAI21_X1  g0772(.A(KEYINPUT42), .B1(new_n680), .B2(new_n950), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n945), .A2(KEYINPUT43), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n960), .A2(new_n953), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n947), .B1(new_n969), .B2(new_n978), .ZN(G387));
  OAI211_X1 g0779(.A(new_n686), .B(new_n277), .C1(new_n313), .C2(new_n269), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n253), .A2(new_n202), .ZN(new_n981));
  XNOR2_X1  g0781(.A(KEYINPUT118), .B(KEYINPUT50), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n783), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n232), .B2(new_n277), .ZN(new_n986));
  INV_X1    g0786(.A(new_n778), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n986), .B1(G107), .B2(new_n210), .C1(new_n686), .C2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n724), .B1(new_n988), .B2(new_n777), .ZN(new_n989));
  INV_X1    g0789(.A(new_n751), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n803), .A2(G77), .B1(new_n990), .B2(G150), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n991), .A2(new_n270), .A3(new_n925), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n749), .A2(G68), .B1(G50), .B2(new_n742), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n993), .B1(new_n386), .B2(new_n740), .C1(new_n252), .C2(new_n745), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n992), .B(new_n994), .C1(new_n443), .C2(new_n736), .ZN(new_n995));
  AOI22_X1  g0795(.A1(G303), .A2(new_n749), .B1(new_n741), .B2(G322), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n816), .B2(new_n745), .C1(new_n774), .C2(new_n926), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n998), .A2(KEYINPUT48), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(KEYINPUT48), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n803), .A2(G294), .B1(new_n736), .B2(G283), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1003), .A2(KEYINPUT49), .ZN(new_n1004));
  INV_X1    g0804(.A(G326), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n265), .B1(new_n751), .B2(new_n1005), .C1(new_n479), .C2(new_n756), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(new_n1003), .B2(KEYINPUT49), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n995), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n989), .B1(new_n1008), .B2(new_n730), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(new_n678), .B2(new_n727), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n965), .B2(new_n948), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n720), .A2(new_n965), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1012), .A2(KEYINPUT119), .A3(new_n684), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n720), .B2(new_n965), .ZN(new_n1014));
  AOI21_X1  g0814(.A(KEYINPUT119), .B1(new_n1012), .B2(new_n684), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1011), .B1(new_n1014), .B2(new_n1015), .ZN(G393));
  NAND2_X1  g0816(.A1(new_n961), .A2(new_n948), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n953), .A2(new_n727), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT120), .Z(new_n1019));
  NOR2_X1   g0819(.A1(new_n243), .A2(new_n783), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n777), .B1(new_n571), .B2(new_n210), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n533), .A2(new_n748), .B1(new_n745), .B2(new_n733), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n803), .A2(G283), .B1(new_n990), .B2(G322), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1023), .B(new_n265), .C1(new_n434), .C2(new_n756), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1022), .B(new_n1024), .C1(G116), .C2(new_n736), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n742), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n1026), .A2(new_n816), .B1(new_n926), .B2(new_n740), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT52), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n1026), .A2(new_n386), .B1(new_n807), .B2(new_n740), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT51), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n202), .A2(new_n745), .B1(new_n748), .B2(new_n252), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n737), .A2(new_n269), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n270), .B1(new_n756), .B2(new_n594), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n732), .A2(new_n313), .B1(new_n751), .B2(new_n808), .ZN(new_n1034));
  NOR4_X1   g0834(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1025), .A2(new_n1028), .B1(new_n1030), .B2(new_n1035), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n790), .B1(new_n1020), .B2(new_n1021), .C1(new_n1036), .C2(new_n730), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n966), .A2(new_n684), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n961), .B1(new_n720), .B2(new_n965), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1017), .B1(new_n1019), .B2(new_n1037), .C1(new_n1038), .C2(new_n1039), .ZN(G390));
  NAND2_X1  g0840(.A1(new_n795), .A2(G330), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n906), .A2(new_n1041), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n878), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n849), .A2(new_n860), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n834), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n671), .B1(new_n715), .B2(new_n658), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n794), .A2(new_n791), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n879), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1045), .B1(new_n1049), .B2(new_n878), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n881), .A2(KEYINPUT39), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n849), .A2(new_n850), .A3(new_n860), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n878), .A2(new_n880), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1053), .B1(new_n1054), .B2(new_n834), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1043), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n834), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n861), .A2(new_n867), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n704), .A2(new_n878), .A3(new_n795), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n792), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n878), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1059), .B(new_n1060), .C1(new_n1063), .C2(new_n1045), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1056), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n885), .A2(G330), .A3(new_n896), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n886), .A2(new_n645), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n878), .B1(new_n704), .B2(new_n795), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n880), .B1(new_n1068), .B2(new_n1043), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1060), .B(new_n1061), .C1(new_n878), .C2(new_n1042), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1065), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1071), .A2(new_n1056), .A3(new_n1064), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1073), .A2(new_n684), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1056), .A2(new_n1064), .A3(new_n948), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n1026), .A2(new_n479), .B1(new_n571), .B2(new_n748), .ZN(new_n1077));
  NOR4_X1   g0877(.A1(new_n1032), .A2(new_n762), .A3(new_n802), .A4(new_n270), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1078), .B1(new_n434), .B2(new_n745), .C1(new_n533), .C2(new_n754), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1077), .B(new_n1079), .C1(G283), .C2(new_n741), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(KEYINPUT121), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n803), .A2(G150), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT53), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G132), .B2(new_n742), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n918), .B2(new_n745), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n270), .B1(new_n756), .B2(new_n202), .C1(new_n737), .C2(new_n386), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n755), .B2(G125), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT54), .B(G143), .Z(new_n1088));
  AOI22_X1  g0888(.A1(G128), .A2(new_n741), .B1(new_n749), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1081), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1080), .A2(KEYINPUT121), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n729), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n724), .B1(new_n252), .B2(new_n821), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1093), .B(new_n1094), .C1(new_n1053), .C2(new_n726), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1075), .A2(new_n1076), .A3(new_n1095), .ZN(G378));
  INV_X1    g0896(.A(new_n1067), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n261), .A2(new_n665), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n309), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n309), .A2(new_n1098), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1101), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n881), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n904), .B1(new_n899), .B2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n902), .A2(new_n878), .A3(new_n795), .A4(new_n896), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1106), .A2(G330), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1104), .B1(new_n1108), .B2(KEYINPUT123), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT123), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1106), .A2(new_n1110), .A3(G330), .A4(new_n1107), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n868), .A2(new_n882), .A3(new_n883), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1109), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n905), .A2(new_n884), .A3(new_n1110), .A4(G330), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1110), .B1(new_n905), .B2(G330), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1116), .B(new_n1117), .C1(new_n1118), .C2(new_n1104), .ZN(new_n1119));
  AOI221_X4 g0919(.A(KEYINPUT57), .B1(new_n1074), .B2(new_n1097), .C1(new_n1115), .C2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT57), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1074), .A2(new_n1097), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n684), .B1(new_n1120), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1122), .A2(new_n948), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n821), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n790), .B1(G50), .B2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT122), .Z(new_n1129));
  NAND2_X1  g0929(.A1(new_n741), .A2(G125), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n749), .A2(G137), .B1(G128), .B2(new_n742), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n803), .A2(new_n1088), .B1(new_n736), .B2(G150), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n931), .A2(G132), .ZN(new_n1133));
  AND4_X1   g0933(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n1135), .A2(KEYINPUT59), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(KEYINPUT59), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n317), .B(new_n276), .C1(new_n756), .C2(new_n386), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G124), .B2(new_n990), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1136), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(G97), .A2(new_n931), .B1(new_n749), .B2(new_n443), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n817), .B2(new_n754), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n270), .A2(G41), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(G77), .B2(new_n803), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1145), .B(new_n917), .C1(new_n381), .C2(new_n756), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n1026), .A2(new_n434), .B1(new_n479), .B2(new_n740), .ZN(new_n1147));
  NOR3_X1   g0947(.A1(new_n1142), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(KEYINPUT58), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1148), .A2(KEYINPUT58), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1144), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1151));
  AND4_X1   g0951(.A1(new_n1140), .A2(new_n1149), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1104), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1129), .B1(new_n730), .B2(new_n1152), .C1(new_n1153), .C2(new_n726), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1126), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1125), .A2(new_n1156), .ZN(G375));
  NAND3_X1  g0957(.A1(new_n1069), .A2(new_n1070), .A3(new_n1067), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1072), .A2(new_n968), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1062), .A2(new_n725), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n790), .B1(G68), .B2(new_n1127), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n434), .A2(new_n748), .B1(new_n740), .B2(new_n533), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G116), .B2(new_n931), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n755), .A2(G303), .B1(new_n742), .B2(G283), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n265), .B1(new_n756), .B2(new_n269), .C1(new_n571), .C2(new_n732), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n443), .B2(new_n736), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1164), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n755), .A2(G128), .B1(G159), .B2(new_n803), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT125), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n741), .A2(G132), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT124), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n270), .B1(new_n756), .B2(new_n381), .C1(new_n737), .C2(new_n202), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n931), .B2(new_n1088), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n807), .B2(new_n748), .C1(new_n918), .C2(new_n774), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1168), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1162), .B1(new_n1177), .B2(new_n729), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1160), .A2(new_n948), .B1(new_n1161), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1159), .A2(new_n1179), .ZN(G381));
  OR2_X1    g0980(.A1(G387), .A2(G390), .ZN(new_n1181));
  OR2_X1    g0981(.A1(G393), .A2(G396), .ZN(new_n1182));
  NOR4_X1   g0982(.A1(new_n1181), .A2(G384), .A3(G381), .A4(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(G375), .A2(G378), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(G407));
  INV_X1    g0985(.A(new_n1184), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n667), .A2(new_n668), .A3(G213), .ZN(new_n1187));
  OAI211_X1 g0987(.A(G407), .B(G213), .C1(new_n1186), .C2(new_n1187), .ZN(G409));
  NAND2_X1  g0988(.A1(G387), .A2(G390), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1181), .A2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(G393), .B(G396), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1190), .B(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT62), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(KEYINPUT126), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1125), .A2(G378), .A3(new_n1156), .ZN(new_n1195));
  INV_X1    g0995(.A(G378), .ZN(new_n1196));
  AND3_X1   g0996(.A1(new_n1122), .A2(new_n968), .A3(new_n1123), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1196), .B1(new_n1155), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1195), .A2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1158), .B(KEYINPUT60), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1200), .A2(new_n684), .A3(new_n1072), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n1179), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n824), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(G384), .A3(new_n1179), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1193), .A2(KEYINPUT126), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AND4_X1   g1008(.A1(new_n1187), .A2(new_n1199), .A3(new_n1206), .A4(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1187), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1208), .B1(new_n1211), .B2(new_n1206), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1194), .B1(new_n1209), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT61), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1210), .A2(G2897), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1205), .B(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1214), .B1(new_n1217), .B2(new_n1211), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1192), .B1(new_n1213), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1199), .A2(new_n1187), .A3(new_n1206), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT63), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1192), .B(new_n1214), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(KEYINPUT63), .B1(new_n1217), .B2(new_n1211), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1223), .B1(new_n1221), .B2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(KEYINPUT127), .B1(new_n1220), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1223), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1224), .A2(new_n1221), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT127), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1221), .A2(new_n1207), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1211), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1218), .B1(new_n1233), .B2(new_n1194), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1229), .B(new_n1230), .C1(new_n1234), .C2(new_n1192), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1226), .A2(new_n1235), .ZN(G405));
  XNOR2_X1  g1036(.A(new_n1192), .B(new_n1206), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(G375), .B(G378), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1237), .B(new_n1238), .ZN(G402));
endmodule


