//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n559, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n620, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1210, new_n1211, new_n1212, new_n1213;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT67), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT68), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G221), .A3(G219), .A4(G220), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  OR2_X1    g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT69), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  NAND2_X1  g032(.A1(G113), .A2(G2104), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n458), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n467), .B1(new_n461), .B2(KEYINPUT3), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n459), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n468), .A2(new_n469), .A3(new_n462), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(G137), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(G101), .A3(G2104), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n473), .B(KEYINPUT71), .ZN(new_n474));
  AND3_X1   g049(.A1(new_n466), .A2(new_n472), .A3(new_n474), .ZN(G160));
  NAND4_X1  g050(.A1(new_n468), .A2(new_n469), .A3(new_n471), .A4(new_n462), .ZN(new_n476));
  INV_X1    g051(.A(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n471), .A2(G112), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  OAI22_X1  g054(.A1(new_n476), .A2(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n470), .A2(G2105), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT72), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n480), .B1(new_n482), .B2(G124), .ZN(G162));
  INV_X1    g058(.A(new_n463), .ZN(new_n484));
  INV_X1    g059(.A(G138), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT73), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT73), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  AND3_X1   g065(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n468), .A2(new_n469), .A3(new_n486), .A4(new_n462), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n484), .A2(new_n491), .B1(new_n492), .B2(KEYINPUT4), .ZN(new_n493));
  AND2_X1   g068(.A1(G126), .A2(G2105), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n468), .A2(new_n469), .A3(new_n462), .A4(new_n494), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G114), .C2(new_n471), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n493), .A2(new_n498), .ZN(G164));
  AND2_X1   g074(.A1(KEYINPUT74), .A2(KEYINPUT5), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT74), .A2(KEYINPUT5), .ZN(new_n501));
  OAI21_X1  g076(.A(G543), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT75), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT75), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n506), .B(G543), .C1(new_n500), .C2(new_n501), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n503), .A2(new_n505), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  XOR2_X1   g085(.A(KEYINPUT76), .B(G88), .Z(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n508), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NAND4_X1  g090(.A1(new_n503), .A2(G62), .A3(new_n505), .A4(new_n507), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n512), .B(new_n514), .C1(new_n518), .C2(KEYINPUT77), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n518), .A2(KEYINPUT77), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(G166));
  OR2_X1    g096(.A1(KEYINPUT79), .A2(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT79), .A2(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n524), .B(new_n526), .ZN(new_n527));
  XOR2_X1   g102(.A(KEYINPUT78), .B(G51), .Z(new_n528));
  NAND2_X1  g103(.A1(new_n513), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n503), .A2(new_n505), .A3(new_n507), .ZN(new_n530));
  NAND2_X1  g105(.A1(G63), .A2(G651), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n527), .B(new_n529), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n509), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n532), .A2(new_n534), .ZN(G168));
  INV_X1    g110(.A(new_n505), .ZN(new_n536));
  OR2_X1    g111(.A1(KEYINPUT74), .A2(KEYINPUT5), .ZN(new_n537));
  NAND2_X1  g112(.A1(KEYINPUT74), .A2(KEYINPUT5), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n504), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n536), .B1(new_n539), .B2(new_n506), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT81), .B(G90), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n540), .A2(new_n503), .A3(new_n508), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n513), .A2(G52), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n503), .A2(G64), .A3(new_n505), .A4(new_n507), .ZN(new_n544));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n515), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n542), .B(new_n543), .C1(new_n546), .C2(KEYINPUT80), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n546), .A2(KEYINPUT80), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(G171));
  NAND2_X1  g124(.A1(new_n513), .A2(G43), .ZN(new_n550));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n509), .B2(new_n551), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n503), .A2(G56), .A3(new_n505), .A4(new_n507), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n515), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT82), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n530), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n508), .A2(G53), .A3(G543), .ZN(new_n567));
  AND2_X1   g142(.A1(KEYINPUT83), .A2(KEYINPUT9), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n567), .B(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G91), .ZN(new_n570));
  OAI211_X1 g145(.A(new_n566), .B(new_n569), .C1(new_n570), .C2(new_n509), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  OR2_X1    g148(.A1(new_n519), .A2(new_n520), .ZN(G303));
  NAND2_X1  g149(.A1(new_n513), .A2(G49), .ZN(new_n575));
  INV_X1    g150(.A(G87), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n509), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(G74), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n515), .B1(new_n530), .B2(new_n578), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n577), .A2(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(new_n513), .A2(G48), .ZN(new_n581));
  INV_X1    g156(.A(G86), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n509), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n503), .A2(G61), .A3(new_n505), .A4(new_n507), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n515), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n510), .A2(G85), .B1(G47), .B2(new_n513), .ZN(new_n589));
  NAND2_X1  g164(.A1(G72), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G60), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n530), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G651), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n530), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(G54), .B2(new_n513), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  OAI21_X1  g175(.A(KEYINPUT84), .B1(new_n509), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  NOR3_X1   g177(.A1(new_n509), .A2(KEYINPUT84), .A3(new_n600), .ZN(new_n603));
  NOR3_X1   g178(.A1(new_n602), .A2(KEYINPUT10), .A3(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  OR3_X1    g180(.A1(new_n509), .A2(KEYINPUT84), .A3(new_n600), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(new_n601), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n599), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(KEYINPUT85), .ZN(new_n609));
  OAI21_X1  g184(.A(KEYINPUT10), .B1(new_n602), .B2(new_n603), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n606), .A2(new_n605), .A3(new_n601), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT85), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n612), .A2(new_n613), .A3(new_n599), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n595), .B1(new_n615), .B2(G868), .ZN(G284));
  OAI21_X1  g191(.A(new_n595), .B1(new_n615), .B2(G868), .ZN(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n569), .B1(new_n570), .B2(new_n509), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(G651), .B2(new_n565), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n618), .B1(new_n620), .B2(G868), .ZN(G297));
  XOR2_X1   g196(.A(G297), .B(KEYINPUT86), .Z(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n615), .B1(new_n623), .B2(G860), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT87), .ZN(G148));
  INV_X1    g200(.A(new_n614), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n613), .B1(new_n612), .B2(new_n599), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g206(.A(G135), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n471), .A2(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  OAI22_X1  g209(.A1(new_n476), .A2(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n482), .B2(G123), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n637), .A2(G2096), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(G2096), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT88), .B(KEYINPUT12), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n471), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2100), .Z(new_n644));
  NAND3_X1  g219(.A1(new_n638), .A2(new_n639), .A3(new_n644), .ZN(G156));
  INV_X1    g220(.A(G14), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(KEYINPUT14), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  AND2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT89), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n646), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n661), .B2(new_n658), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT90), .ZN(G401));
  XOR2_X1   g239(.A(KEYINPUT91), .B(KEYINPUT18), .Z(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2096), .B(G2100), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT92), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2072), .B(G2078), .Z(new_n675));
  INV_X1    g250(.A(new_n665), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n675), .B1(new_n668), .B2(new_n676), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n674), .A2(new_n677), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(G227));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT93), .ZN(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  NAND3_X1  g264(.A1(new_n686), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n686), .B1(new_n688), .B2(new_n689), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n688), .A2(new_n689), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n691), .B(new_n694), .C1(new_n685), .C2(new_n693), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G1981), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n695), .A2(G1981), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n683), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n695), .A2(G1981), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n700), .A2(G1986), .A3(new_n696), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT94), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n699), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n704), .B1(new_n699), .B2(new_n701), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n682), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n707), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n709), .A2(new_n681), .A3(new_n705), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n708), .A2(new_n710), .ZN(G229));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G26), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  INV_X1    g289(.A(G140), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n476), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n717));
  INV_X1    g292(.A(G116), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(G2105), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n482), .B2(G128), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n714), .B1(new_n722), .B2(new_n712), .ZN(new_n723));
  INV_X1    g298(.A(G2067), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT30), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n726), .A2(G28), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n712), .B1(new_n726), .B2(G28), .ZN(new_n728));
  AND2_X1   g303(.A1(KEYINPUT31), .A2(G11), .ZN(new_n729));
  NOR2_X1   g304(.A1(KEYINPUT31), .A2(G11), .ZN(new_n730));
  OAI22_X1  g305(.A1(new_n727), .A2(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n636), .B2(G29), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT101), .B(KEYINPUT24), .ZN(new_n733));
  INV_X1    g308(.A(G34), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n735), .A2(new_n712), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT102), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G29), .B2(G160), .ZN(new_n740));
  INV_X1    g315(.A(G2084), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n712), .A2(G27), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G164), .B2(new_n712), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT104), .B(G2078), .Z(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n725), .A2(new_n732), .A3(new_n742), .A4(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G16), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G20), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT23), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n620), .B2(new_n748), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1956), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n748), .A2(G21), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G168), .B2(new_n748), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1966), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n712), .A2(G32), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT26), .Z(new_n758));
  NAND3_X1  g333(.A1(new_n471), .A2(G105), .A3(G2104), .ZN(new_n759));
  INV_X1    g334(.A(G141), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n758), .B(new_n759), .C1(new_n760), .C2(new_n476), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n482), .B2(G129), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n756), .B1(new_n762), .B2(new_n712), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT27), .B(G1996), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NOR4_X1   g340(.A1(new_n747), .A2(new_n752), .A3(new_n755), .A4(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G29), .A2(G35), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G162), .B2(G29), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT29), .ZN(new_n769));
  INV_X1    g344(.A(G2090), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G16), .A2(G19), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n556), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT98), .B(G1341), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(G115), .A2(G2104), .ZN(new_n776));
  INV_X1    g351(.A(G127), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n463), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G2105), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT100), .Z(new_n780));
  INV_X1    g355(.A(KEYINPUT99), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT25), .Z(new_n783));
  INV_X1    g358(.A(G139), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n476), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n780), .B1(new_n781), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n785), .A2(new_n781), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(new_n712), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n712), .B2(G33), .ZN(new_n790));
  INV_X1    g365(.A(G2072), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n790), .A2(new_n791), .B1(new_n773), .B2(new_n774), .ZN(new_n792));
  AND4_X1   g367(.A1(new_n766), .A2(new_n771), .A3(new_n775), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n748), .A2(G5), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G171), .B2(new_n748), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n795), .A2(G1961), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n795), .A2(G1961), .ZN(new_n797));
  OR3_X1    g372(.A1(new_n790), .A2(KEYINPUT103), .A3(new_n791), .ZN(new_n798));
  OAI21_X1  g373(.A(KEYINPUT103), .B1(new_n790), .B2(new_n791), .ZN(new_n799));
  AOI211_X1 g374(.A(new_n796), .B(new_n797), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n748), .A2(G4), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n615), .B2(new_n748), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT97), .B(G1348), .Z(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n802), .A2(new_n804), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n793), .A2(new_n800), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n748), .A2(G23), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G288), .B2(G16), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT33), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G1976), .ZN(new_n814));
  INV_X1    g389(.A(G1976), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n811), .A2(new_n815), .A3(new_n812), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  OR2_X1    g392(.A1(G16), .A2(G22), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G303), .B2(new_n748), .ZN(new_n819));
  INV_X1    g394(.A(G1971), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n748), .A2(G6), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n587), .B2(new_n748), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT32), .B(G1981), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT95), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n824), .B(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n821), .A2(new_n822), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(KEYINPUT34), .B1(new_n817), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT96), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n814), .A2(new_n816), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n832), .A2(new_n822), .A3(new_n821), .A4(new_n827), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n833), .A2(KEYINPUT96), .A3(KEYINPUT34), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n833), .A2(KEYINPUT34), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n712), .A2(G25), .ZN(new_n837));
  INV_X1    g412(.A(G131), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n476), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n840));
  INV_X1    g415(.A(G107), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n840), .B1(new_n841), .B2(G2105), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n482), .B2(G119), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n837), .B1(new_n845), .B2(new_n712), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT35), .B(G1991), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  MUX2_X1   g423(.A(G24), .B(G290), .S(G16), .Z(new_n849));
  OR2_X1    g424(.A1(new_n849), .A2(G1986), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(G1986), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n848), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n836), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n835), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT36), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT36), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n835), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n807), .B1(new_n855), .B2(new_n857), .ZN(G311));
  INV_X1    g433(.A(new_n807), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n835), .A2(new_n853), .A3(new_n856), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n856), .B1(new_n835), .B2(new_n853), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(G150));
  NAND2_X1  g437(.A1(G80), .A2(G543), .ZN(new_n863));
  INV_X1    g438(.A(G67), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n530), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(G651), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n513), .A2(G55), .ZN(new_n867));
  INV_X1    g442(.A(G93), .ZN(new_n868));
  OAI211_X1 g443(.A(KEYINPUT105), .B(new_n867), .C1(new_n509), .C2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n540), .A2(G93), .A3(new_n503), .A4(new_n508), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT105), .B1(new_n871), .B2(new_n867), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n866), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(KEYINPUT106), .B(G860), .Z(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT37), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n615), .A2(G559), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT38), .ZN(new_n879));
  INV_X1    g454(.A(new_n556), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n873), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n556), .B(new_n866), .C1(new_n872), .C2(new_n870), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n879), .B(new_n883), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n884), .A2(KEYINPUT39), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n875), .B1(new_n884), .B2(KEYINPUT39), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n877), .B1(new_n885), .B2(new_n886), .ZN(G145));
  INV_X1    g462(.A(KEYINPUT72), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n481), .B(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(G128), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n720), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n491), .A2(new_n484), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n495), .A2(new_n497), .A3(KEYINPUT107), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT107), .B1(new_n495), .B2(new_n497), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n891), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n897), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n493), .B1(new_n900), .B2(new_n895), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n722), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n902), .A3(new_n762), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n762), .B1(new_n899), .B2(new_n902), .ZN(new_n905));
  OAI211_X1 g480(.A(KEYINPUT108), .B(new_n788), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n899), .A2(new_n902), .ZN(new_n907));
  INV_X1    g482(.A(new_n762), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n788), .A2(KEYINPUT108), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(new_n786), .B2(new_n787), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n909), .A2(new_n910), .A3(new_n912), .A4(new_n903), .ZN(new_n913));
  INV_X1    g488(.A(new_n642), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n845), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G119), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n843), .B1(new_n889), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n642), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n470), .A2(G142), .A3(new_n471), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT109), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n471), .A2(G118), .ZN(new_n921));
  OAI21_X1  g496(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n922));
  INV_X1    g497(.A(G130), .ZN(new_n923));
  OAI221_X1 g498(.A(new_n920), .B1(new_n921), .B2(new_n922), .C1(new_n889), .C2(new_n923), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n915), .A2(new_n918), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n924), .B1(new_n915), .B2(new_n918), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n906), .A2(new_n913), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n927), .B1(new_n906), .B2(new_n913), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g505(.A(G162), .B(new_n636), .Z(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(G160), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n906), .A2(new_n913), .ZN(new_n934));
  INV_X1    g509(.A(new_n927), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n906), .A2(new_n913), .A3(new_n927), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n932), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT110), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI211_X1 g515(.A(KEYINPUT110), .B(new_n939), .C1(new_n928), .C2(new_n929), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n933), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g519(.A1(new_n881), .A2(new_n882), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n615), .A2(new_n623), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n945), .B1(new_n615), .B2(new_n623), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n612), .A2(new_n620), .A3(new_n599), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n620), .B1(new_n612), .B2(new_n599), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n947), .A2(new_n948), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n628), .A2(new_n883), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT41), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(new_n950), .B2(new_n951), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n608), .A2(G299), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n957), .A2(KEYINPUT41), .A3(new_n949), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n954), .A2(new_n946), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT42), .B1(new_n953), .B2(new_n959), .ZN(new_n960));
  XOR2_X1   g535(.A(G290), .B(G288), .Z(new_n961));
  NOR2_X1   g536(.A1(G303), .A2(new_n587), .ZN(new_n962));
  NOR2_X1   g537(.A1(G166), .A2(G305), .ZN(new_n963));
  OR3_X1    g538(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT41), .B1(new_n957), .B2(new_n949), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n957), .A2(KEYINPUT41), .A3(new_n949), .ZN(new_n969));
  OAI22_X1  g544(.A1(new_n947), .A2(new_n948), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n954), .B(new_n946), .C1(new_n951), .C2(new_n950), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n960), .A2(new_n967), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n967), .B1(new_n960), .B2(new_n973), .ZN(new_n975));
  OAI21_X1  g550(.A(G868), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n874), .A2(G868), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(G295));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n977), .ZN(G331));
  OAI21_X1  g554(.A(G286), .B1(new_n547), .B2(new_n548), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n546), .A2(KEYINPUT80), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n546), .A2(KEYINPUT80), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n542), .A2(new_n543), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n981), .A2(G168), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n945), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n881), .A2(new_n980), .A3(new_n984), .A4(new_n882), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n883), .A2(KEYINPUT111), .A3(new_n980), .A4(new_n984), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n969), .A2(new_n968), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n986), .A2(new_n993), .A3(new_n988), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n945), .A2(new_n985), .A3(KEYINPUT112), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n991), .A2(new_n992), .B1(new_n996), .B2(new_n952), .ZN(new_n997));
  AOI21_X1  g572(.A(G37), .B1(new_n997), .B2(new_n966), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n952), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n956), .A2(new_n989), .A3(new_n958), .A4(new_n990), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n967), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT43), .B1(new_n998), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(new_n966), .A3(new_n1000), .ZN(new_n1004));
  INV_X1    g579(.A(G37), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT43), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n989), .A2(new_n990), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n952), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n956), .A2(new_n994), .A3(new_n958), .A4(new_n995), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n966), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n1006), .A2(new_n1007), .A3(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT44), .B1(new_n1003), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1007), .B1(new_n998), .B2(new_n1002), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1006), .A2(KEYINPUT43), .A3(new_n1011), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1013), .A2(new_n1017), .ZN(G397));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(new_n901), .B2(G1384), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n466), .A2(new_n472), .A3(G40), .A4(new_n474), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n762), .B(G1996), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n722), .B(G2067), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n845), .B(new_n847), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(G290), .B(G1986), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1022), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1021), .ZN(new_n1031));
  INV_X1    g606(.A(G1384), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(new_n898), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(G8), .ZN(new_n1034));
  OAI21_X1  g609(.A(G1981), .B1(new_n586), .B2(KEYINPUT114), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n586), .B2(new_n583), .ZN(new_n1036));
  INV_X1    g611(.A(new_n583), .ZN(new_n1037));
  INV_X1    g612(.A(new_n586), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(KEYINPUT114), .A4(G1981), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1036), .A2(new_n1039), .A3(KEYINPUT115), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1034), .B1(new_n1040), .B2(KEYINPUT49), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT49), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1036), .A2(new_n1039), .A3(KEYINPUT115), .A4(new_n1043), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1042), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1033), .B(G8), .C1(G288), .C2(new_n815), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(G288), .B2(new_n815), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1051));
  OAI22_X1  g626(.A1(new_n1045), .A2(new_n1046), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G8), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n898), .A2(KEYINPUT45), .A3(new_n1032), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1032), .B1(new_n493), .B2(new_n498), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1019), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n1031), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n820), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1021), .B1(new_n1055), .B2(KEYINPUT50), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n898), .A2(new_n1060), .A3(new_n1032), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1059), .A2(new_n770), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1053), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(G8), .B1(new_n519), .B2(new_n520), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n1067));
  OAI211_X1 g642(.A(KEYINPUT55), .B(G8), .C1(new_n519), .C2(new_n520), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1067), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1063), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1031), .B1(new_n1055), .B2(KEYINPUT50), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1060), .B1(new_n898), .B2(new_n1032), .ZN(new_n1073));
  OR3_X1    g648(.A1(new_n1072), .A2(new_n1073), .A3(G2090), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1053), .B1(new_n1074), .B2(new_n1058), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1071), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1052), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1057), .B2(G2078), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1082));
  INV_X1    g657(.A(G1961), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1080), .A2(G2078), .ZN(new_n1085));
  OAI211_X1 g660(.A(KEYINPUT45), .B(new_n1032), .C1(new_n493), .C2(new_n498), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1020), .A2(new_n1031), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1081), .A2(new_n1084), .A3(new_n1087), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1088), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT123), .B1(new_n1088), .B2(G171), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1966), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1031), .A2(new_n1086), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT45), .B1(new_n898), .B2(new_n1032), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1059), .A2(new_n1061), .A3(new_n741), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(G8), .ZN(new_n1099));
  OR3_X1    g674(.A1(G168), .A2(KEYINPUT121), .A3(new_n1053), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT121), .B1(G168), .B2(new_n1053), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1099), .A2(KEYINPUT122), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT122), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1053), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1103), .A2(new_n1107), .A3(KEYINPUT51), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1098), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n1107), .B2(KEYINPUT51), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT62), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  OR2_X1    g686(.A1(new_n1107), .A2(KEYINPUT51), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1103), .A2(new_n1107), .A3(KEYINPUT51), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .A4(new_n1109), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1079), .A2(new_n1092), .A3(new_n1111), .A4(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(G288), .A2(G1976), .ZN(new_n1117));
  XOR2_X1   g692(.A(new_n1117), .B(KEYINPUT117), .Z(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1119));
  OR2_X1    g694(.A1(G305), .A2(G1981), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1034), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1105), .A2(new_n1123), .A3(G168), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1123), .B1(new_n1105), .B2(G168), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT63), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1071), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1051), .A2(new_n1049), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1046), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1121), .A2(new_n1122), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1134));
  OAI22_X1  g709(.A1(new_n1124), .A2(new_n1125), .B1(new_n1076), .B2(new_n1063), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT63), .B1(new_n1052), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1116), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1112), .A2(new_n1113), .A3(new_n1109), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1071), .A2(new_n1077), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1020), .A2(new_n1031), .A3(new_n1054), .A4(new_n1085), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1081), .A2(new_n1084), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(G171), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1142), .B(KEYINPUT54), .C1(G171), .C2(new_n1088), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1133), .A2(new_n1138), .A3(new_n1139), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1082), .A2(new_n803), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1033), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n724), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT57), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n620), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(G1956), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1151), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1152));
  NAND2_X1  g727(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT56), .B(G2072), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1054), .A2(new_n1056), .A3(new_n1031), .A4(new_n1154), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1150), .A2(new_n1152), .A3(new_n1153), .A4(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n615), .A2(new_n1148), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT120), .B1(new_n626), .B2(new_n627), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n609), .A2(new_n1163), .A3(new_n614), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1145), .A2(new_n1147), .A3(KEYINPUT60), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1162), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT60), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1148), .A2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1165), .A2(new_n609), .A3(new_n1163), .A4(new_n614), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1167), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  XOR2_X1   g746(.A(KEYINPUT58), .B(G1341), .Z(new_n1172));
  NAND2_X1  g747(.A1(new_n1033), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(G1996), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1054), .A2(new_n1056), .A3(new_n1174), .A4(new_n1031), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n880), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT59), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1177), .A2(KEYINPUT119), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1176), .B(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1160), .A2(new_n1156), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(KEYINPUT61), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1160), .A2(new_n1182), .A3(new_n1156), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1179), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1161), .B1(new_n1171), .B2(new_n1184), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n1141), .A2(G171), .ZN(new_n1186));
  AOI21_X1  g761(.A(KEYINPUT54), .B1(new_n1091), .B2(new_n1186), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1144), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1030), .B1(new_n1137), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1022), .A2(new_n1174), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(KEYINPUT46), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1024), .A2(new_n762), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(new_n1022), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT125), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1194), .B(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1196), .B(KEYINPUT47), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1022), .A2(new_n683), .A3(new_n593), .A4(new_n589), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1198), .ZN(new_n1199));
  AOI22_X1  g774(.A1(new_n1028), .A2(new_n1022), .B1(KEYINPUT48), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1200), .B1(KEYINPUT48), .B2(new_n1199), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n845), .A2(new_n847), .ZN(new_n1202));
  XOR2_X1   g777(.A(new_n1202), .B(KEYINPUT124), .Z(new_n1203));
  OAI22_X1  g778(.A1(new_n1203), .A2(new_n1025), .B1(G2067), .B2(new_n891), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1022), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1201), .A2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1197), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1189), .A2(new_n1207), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g783(.A(G319), .B1(new_n678), .B2(new_n679), .ZN(new_n1210));
  XOR2_X1   g784(.A(new_n1210), .B(KEYINPUT126), .Z(new_n1211));
  NAND2_X1  g785(.A1(new_n663), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g786(.A(new_n1212), .B1(new_n708), .B2(new_n710), .ZN(new_n1213));
  OAI211_X1 g787(.A(new_n943), .B(new_n1213), .C1(new_n1015), .C2(new_n1016), .ZN(G225));
  INV_X1    g788(.A(G225), .ZN(G308));
endmodule


