//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT32), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT64), .A2(G143), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(G146), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n195), .A2(new_n197), .A3(new_n199), .ZN(new_n200));
  AND2_X1   g014(.A1(KEYINPUT64), .A2(G143), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT64), .A2(G143), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n196), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n196), .A2(G143), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n203), .A2(new_n205), .B1(G128), .B2(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n200), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G134), .B(G137), .ZN(new_n210));
  INV_X1    g024(.A(G131), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OR2_X1    g026(.A1(KEYINPUT67), .A2(KEYINPUT11), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT67), .A2(KEYINPUT11), .ZN(new_n214));
  INV_X1    g028(.A(G137), .ZN(new_n215));
  AOI22_X1  g029(.A1(new_n213), .A2(new_n214), .B1(G134), .B2(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT67), .A2(KEYINPUT11), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(G134), .ZN(new_n218));
  INV_X1    g032(.A(G134), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G137), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n217), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT68), .B(G131), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n212), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n209), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(G131), .B1(new_n216), .B2(new_n221), .ZN(new_n226));
  INV_X1    g040(.A(new_n214), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n218), .B1(new_n227), .B2(new_n217), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n228), .B(new_n223), .C1(new_n217), .C2(new_n210), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT0), .B(G128), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n231), .B1(new_n203), .B2(new_n205), .ZN(new_n232));
  AND2_X1   g046(.A1(KEYINPUT0), .A2(G128), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n195), .A2(new_n197), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n195), .A2(KEYINPUT65), .A3(new_n197), .A4(new_n233), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n232), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n230), .B1(new_n238), .B2(KEYINPUT66), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n240));
  AOI211_X1 g054(.A(new_n240), .B(new_n232), .C1(new_n236), .C2(new_n237), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n225), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT30), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT70), .B1(new_n200), .B2(new_n207), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n195), .A2(new_n197), .A3(new_n199), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT64), .B(G143), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n204), .B1(new_n248), .B2(new_n196), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n198), .B1(new_n197), .B2(KEYINPUT1), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n246), .B(new_n247), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n245), .A2(new_n224), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n236), .A2(new_n237), .ZN(new_n253));
  INV_X1    g067(.A(new_n232), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n230), .A3(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n252), .A2(new_n255), .A3(KEYINPUT30), .ZN(new_n256));
  INV_X1    g070(.A(G116), .ZN(new_n257));
  INV_X1    g071(.A(G119), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(G116), .A2(G119), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT2), .B(G113), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  XOR2_X1   g077(.A(KEYINPUT2), .B(G113), .Z(new_n264));
  NAND2_X1  g078(.A1(new_n259), .A2(new_n260), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT69), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n263), .A2(new_n266), .A3(KEYINPUT69), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n256), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n244), .A2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n269), .A2(new_n270), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(new_n252), .A3(new_n255), .ZN(new_n275));
  INV_X1    g089(.A(G237), .ZN(new_n276));
  INV_X1    g090(.A(G953), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n277), .A3(G210), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n278), .A2(KEYINPUT27), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(KEYINPUT27), .ZN(new_n280));
  OR3_X1    g094(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT26), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n278), .B(KEYINPUT27), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT26), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n281), .A2(G101), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(G101), .B1(new_n281), .B2(new_n283), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n275), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT71), .B1(new_n273), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n290));
  AOI211_X1 g104(.A(new_n290), .B(new_n287), .C1(new_n244), .C2(new_n272), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT31), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT31), .B1(new_n273), .B2(new_n288), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n275), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n296), .B1(new_n242), .B2(new_n271), .ZN(new_n297));
  XOR2_X1   g111(.A(KEYINPUT73), .B(KEYINPUT28), .Z(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI22_X1  g113(.A1(new_n297), .A2(new_n299), .B1(KEYINPUT28), .B2(new_n296), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n286), .B(KEYINPUT72), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT74), .B1(new_n295), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT31), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n256), .A2(new_n271), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n305), .B1(new_n243), .B2(new_n242), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n290), .B1(new_n306), .B2(new_n287), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n273), .A2(KEYINPUT71), .A3(new_n288), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n304), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI211_X1 g123(.A(KEYINPUT74), .B(new_n302), .C1(new_n309), .C2(new_n293), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n190), .B1(new_n303), .B2(new_n311), .ZN(new_n312));
  OR2_X1    g126(.A1(new_n301), .A2(KEYINPUT29), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n300), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n274), .B1(new_n252), .B2(new_n255), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n296), .A2(new_n315), .ZN(new_n316));
  MUX2_X1   g130(.A(new_n296), .B(new_n316), .S(KEYINPUT28), .Z(new_n317));
  AND2_X1   g131(.A1(new_n317), .A2(new_n286), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n273), .A2(new_n275), .ZN(new_n319));
  INV_X1    g133(.A(new_n286), .ZN(new_n320));
  AOI21_X1  g134(.A(KEYINPUT29), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n314), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G902), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G472), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n302), .B1(new_n309), .B2(new_n293), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT74), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n188), .B1(new_n328), .B2(new_n310), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n312), .B(new_n325), .C1(new_n329), .C2(KEYINPUT32), .ZN(new_n330));
  OAI21_X1  g144(.A(G214), .B1(G237), .B2(G902), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT81), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(G234), .A2(G237), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(G952), .A3(new_n277), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(KEYINPUT97), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n334), .A2(G902), .A3(G953), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT21), .B(G898), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G107), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G104), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT3), .B1(new_n343), .B2(KEYINPUT79), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n345), .A2(new_n346), .A3(new_n342), .A4(G104), .ZN(new_n347));
  INV_X1    g161(.A(G104), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G107), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n344), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G101), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n351), .A2(KEYINPUT4), .ZN(new_n352));
  INV_X1    g166(.A(G101), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n344), .A2(new_n353), .A3(new_n347), .A4(new_n349), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n351), .A2(KEYINPUT4), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n271), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n261), .A2(new_n262), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n265), .A2(KEYINPUT5), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT5), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(new_n258), .A3(G116), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G113), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n357), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n353), .B1(new_n343), .B2(new_n349), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT80), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n363), .A2(new_n354), .A3(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G110), .B(G122), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n356), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT85), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT85), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n356), .A2(new_n371), .A3(new_n367), .A4(new_n368), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n343), .A2(new_n349), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n365), .B1(new_n374), .B2(new_n353), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n364), .A2(KEYINPUT80), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n354), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n363), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n368), .B(KEYINPUT8), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n361), .B1(new_n358), .B2(KEYINPUT87), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT87), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n265), .A2(new_n381), .A3(KEYINPUT5), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n357), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n378), .B(new_n379), .C1(new_n377), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT88), .ZN(new_n385));
  OR2_X1    g199(.A1(new_n383), .A2(new_n377), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT88), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n386), .A2(new_n387), .A3(new_n378), .A4(new_n379), .ZN(new_n388));
  INV_X1    g202(.A(G125), .ZN(new_n389));
  MUX2_X1   g203(.A(new_n238), .B(new_n209), .S(new_n389), .Z(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT86), .B(G224), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(G953), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT7), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n385), .A2(new_n388), .B1(new_n390), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT89), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n397), .B1(new_n390), .B2(new_n395), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n209), .A2(G125), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n238), .A2(new_n389), .ZN(new_n400));
  OAI211_X1 g214(.A(KEYINPUT89), .B(new_n394), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n373), .A2(new_n396), .A3(new_n402), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n403), .A2(new_n323), .ZN(new_n404));
  OAI21_X1  g218(.A(G210), .B1(G237), .B2(G902), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(KEYINPUT84), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n356), .A2(KEYINPUT82), .A3(new_n367), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n368), .B(KEYINPUT83), .Z(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(KEYINPUT82), .B1(new_n356), .B2(new_n367), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n356), .A2(new_n367), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT82), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n416), .A2(new_n407), .A3(new_n409), .A4(new_n410), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n370), .A2(KEYINPUT6), .A3(new_n372), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n413), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n390), .B(new_n393), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n404), .A2(new_n405), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n405), .B1(new_n404), .B2(new_n421), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n333), .B(new_n341), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n198), .A2(G119), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT23), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n258), .A2(G128), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G110), .ZN(new_n431));
  XNOR2_X1  g245(.A(G125), .B(G140), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT16), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT16), .ZN(new_n434));
  INV_X1    g248(.A(G140), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n435), .A3(G125), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n433), .A2(G146), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(G146), .B1(new_n433), .B2(new_n436), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n431), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n425), .A2(new_n428), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(KEYINPUT75), .ZN(new_n441));
  XOR2_X1   g255(.A(KEYINPUT24), .B(G110), .Z(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT76), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n441), .A2(KEYINPUT76), .A3(new_n442), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n439), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OAI22_X1  g262(.A1(new_n441), .A2(new_n442), .B1(G110), .B2(new_n430), .ZN(new_n449));
  INV_X1    g263(.A(new_n437), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n432), .A2(new_n196), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n277), .A2(G221), .A3(G234), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(KEYINPUT22), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(G137), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n448), .A2(new_n452), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n455), .ZN(new_n457));
  INV_X1    g271(.A(new_n452), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n457), .B1(new_n458), .B2(new_n447), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT77), .ZN(new_n461));
  INV_X1    g275(.A(G217), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n462), .B1(G234), .B2(new_n323), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(G902), .ZN(new_n464));
  XOR2_X1   g278(.A(new_n464), .B(KEYINPUT78), .Z(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(KEYINPUT25), .B1(new_n460), .B2(G902), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT25), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n456), .A2(new_n459), .A3(new_n469), .A4(new_n323), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n463), .A3(new_n470), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT9), .B(G234), .ZN(new_n473));
  OAI21_X1  g287(.A(G221), .B1(new_n473), .B2(G902), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G469), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(new_n323), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n195), .A2(new_n197), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n198), .B1(new_n203), .B2(KEYINPUT1), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n246), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n366), .A3(new_n354), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT10), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n377), .A2(new_n482), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(new_n245), .A3(new_n251), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n352), .A2(new_n238), .A3(new_n355), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n230), .ZN(new_n488));
  INV_X1    g302(.A(new_n230), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n483), .A2(new_n485), .A3(new_n486), .A4(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(G110), .B(G140), .ZN(new_n491));
  INV_X1    g305(.A(G227), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(G953), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n491), .B(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n208), .A2(new_n377), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n481), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT12), .B1(new_n498), .B2(new_n230), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT12), .ZN(new_n500));
  AOI211_X1 g314(.A(new_n500), .B(new_n489), .C1(new_n481), .C2(new_n497), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n490), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n488), .A2(new_n496), .B1(new_n502), .B2(new_n494), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n477), .B1(new_n503), .B2(G469), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n499), .A2(new_n501), .ZN(new_n505));
  INV_X1    g319(.A(new_n490), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n505), .A2(new_n506), .A3(new_n494), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n495), .B1(new_n488), .B2(new_n490), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n476), .B(new_n323), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n475), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n472), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(KEYINPUT94), .B1(new_n248), .B2(new_n198), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT94), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n193), .A2(new_n513), .A3(G128), .A4(new_n194), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT13), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT13), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n198), .A2(G143), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G134), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n515), .A2(new_n219), .A3(new_n519), .ZN(new_n522));
  INV_X1    g336(.A(G122), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G116), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n257), .A2(G122), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT93), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n524), .A2(new_n525), .A3(KEYINPUT93), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(G107), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n528), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n342), .B1(new_n530), .B2(new_n526), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n522), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n521), .A2(new_n533), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n473), .A2(new_n462), .A3(G953), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT95), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n536), .B1(new_n525), .B2(KEYINPUT14), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT14), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n538), .A2(new_n257), .A3(KEYINPUT95), .A4(G122), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n525), .A2(KEYINPUT14), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n537), .A2(new_n524), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT96), .B1(new_n541), .B2(G107), .ZN(new_n542));
  INV_X1    g356(.A(new_n531), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n541), .A2(KEYINPUT96), .A3(G107), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n219), .B1(new_n515), .B2(new_n519), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n544), .B(new_n545), .C1(new_n522), .C2(new_n546), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n534), .A2(new_n535), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n535), .B1(new_n534), .B2(new_n547), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n323), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(G478), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n551), .A2(KEYINPUT15), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n534), .A2(new_n547), .ZN(new_n554));
  INV_X1    g368(.A(new_n535), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n534), .A2(new_n547), .A3(new_n535), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n552), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n323), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n553), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n437), .A2(new_n438), .ZN(new_n563));
  INV_X1    g377(.A(G214), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n564), .A2(G237), .A3(G953), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G143), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n248), .B2(new_n565), .ZN(new_n567));
  INV_X1    g381(.A(new_n223), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(KEYINPUT17), .A3(new_n568), .ZN(new_n569));
  OR2_X1    g383(.A1(new_n248), .A2(new_n565), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n570), .A2(new_n223), .A3(new_n566), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n567), .A2(new_n568), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n563), .B(new_n569), .C1(new_n573), .C2(KEYINPUT17), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n435), .A2(G125), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n389), .A2(G140), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(G146), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n451), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT90), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n578), .A2(new_n451), .A3(KEYINPUT90), .ZN(new_n582));
  NAND2_X1  g396(.A1(KEYINPUT18), .A2(G131), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n581), .A2(new_n582), .B1(new_n584), .B2(new_n567), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n586), .B1(new_n567), .B2(new_n584), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n570), .A2(KEYINPUT91), .A3(new_n583), .A4(new_n566), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(G113), .B(G122), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(new_n348), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT92), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n574), .A2(new_n590), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n592), .B1(new_n574), .B2(new_n590), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n323), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G475), .ZN(new_n598));
  NOR2_X1   g412(.A1(G475), .A2(G902), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT19), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n577), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n432), .A2(KEYINPUT19), .ZN(new_n603));
  AOI21_X1  g417(.A(G146), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n437), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n573), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n590), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n592), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n574), .A2(new_n590), .A3(new_n594), .ZN(new_n610));
  AOI211_X1 g424(.A(KEYINPUT20), .B(new_n600), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT20), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n585), .A2(new_n589), .B1(new_n605), .B2(new_n573), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n610), .B1(new_n592), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n612), .B1(new_n614), .B2(new_n599), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n598), .B1(new_n611), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n562), .A2(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n424), .A2(new_n511), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n330), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT98), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n623));
  AOI21_X1  g437(.A(G478), .B1(new_n558), .B2(new_n323), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT33), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n625), .B1(new_n548), .B2(new_n549), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n556), .A2(KEYINPUT33), .A3(new_n557), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n551), .A2(G902), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n624), .B1(new_n629), .B2(KEYINPUT99), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n626), .A2(new_n627), .A3(new_n631), .A4(new_n628), .ZN(new_n632));
  AOI211_X1 g446(.A(KEYINPUT100), .B(new_n617), .C1(new_n630), .C2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n629), .A2(KEYINPUT99), .ZN(new_n635));
  INV_X1    g449(.A(new_n624), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n632), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n634), .B1(new_n637), .B2(new_n616), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n623), .B1(new_n639), .B2(new_n424), .ZN(new_n640));
  INV_X1    g454(.A(new_n424), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n641), .B(KEYINPUT101), .C1(new_n638), .C2(new_n633), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n323), .B1(new_n303), .B2(new_n311), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(G472), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n329), .A2(new_n511), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT34), .B(G104), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G6));
  INV_X1    g465(.A(new_n405), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n419), .A2(new_n420), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n403), .A2(new_n323), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n404), .A2(new_n421), .A3(new_n405), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n332), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n611), .ZN(new_n658));
  INV_X1    g472(.A(new_n615), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n598), .A2(KEYINPUT102), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n598), .A2(KEYINPUT102), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n662), .A2(new_n561), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n657), .A2(new_n664), .A3(new_n341), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n641), .A2(KEYINPUT103), .A3(new_n664), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n648), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT35), .B(G107), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  AOI21_X1  g486(.A(new_n329), .B1(new_n644), .B2(G472), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n448), .A2(new_n452), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n457), .A2(KEYINPUT36), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n466), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n471), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT104), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n471), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n424), .A2(new_n618), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n673), .A2(new_n510), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT37), .B(G110), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT105), .B(KEYINPUT106), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G12));
  OAI21_X1  g502(.A(new_n333), .B1(new_n422), .B2(new_n423), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n510), .A2(new_n679), .A3(new_n681), .ZN(new_n690));
  INV_X1    g504(.A(G900), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n337), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n336), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n662), .A2(new_n561), .A3(new_n663), .A4(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n689), .A2(new_n690), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n330), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G128), .ZN(G30));
  INV_X1    g512(.A(new_n510), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n693), .B(KEYINPUT39), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT40), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n187), .B1(new_n303), .B2(new_n311), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n189), .ZN(new_n704));
  INV_X1    g518(.A(G472), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n289), .A2(new_n291), .ZN(new_n706));
  INV_X1    g520(.A(new_n301), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n706), .B1(new_n707), .B2(new_n316), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n705), .B1(new_n708), .B2(new_n323), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n328), .A2(new_n310), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n709), .B1(new_n710), .B2(new_n190), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n704), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n655), .A2(new_n656), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT38), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n561), .A2(new_n616), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n715), .A2(new_n678), .A3(new_n332), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n702), .A2(new_n712), .A3(new_n714), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT107), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n248), .ZN(G45));
  NAND3_X1  g533(.A1(new_n637), .A2(new_n616), .A3(new_n694), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n689), .A2(new_n690), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n330), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT108), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n330), .A2(new_n724), .A3(new_n721), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G146), .ZN(G48));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n323), .B1(new_n507), .B2(new_n508), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(G469), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n509), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n728), .B1(new_n731), .B2(new_n475), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n730), .A2(KEYINPUT109), .A3(new_n474), .A4(new_n509), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(new_n472), .A3(new_n733), .ZN(new_n734));
  AOI22_X1  g548(.A1(new_n710), .A2(new_n190), .B1(G472), .B2(new_n324), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n734), .B1(new_n704), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n643), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT41), .B(G113), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT110), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n737), .B(new_n739), .ZN(G15));
  NAND2_X1  g554(.A1(new_n669), .A2(new_n736), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G116), .ZN(G18));
  NAND2_X1  g556(.A1(new_n732), .A2(new_n733), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n743), .B1(new_n704), .B2(new_n735), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n683), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G119), .ZN(G21));
  OAI21_X1  g560(.A(new_n295), .B1(new_n707), .B2(new_n317), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n187), .ZN(new_n748));
  AOI21_X1  g562(.A(G902), .B1(new_n328), .B2(new_n310), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n472), .B(new_n748), .C1(new_n749), .C2(new_n705), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n732), .A2(new_n341), .A3(new_n733), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n715), .A2(KEYINPUT111), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n550), .A2(new_n552), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n559), .B1(new_n558), .B2(new_n323), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n616), .B(new_n754), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(KEYINPUT112), .B1(new_n689), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n757), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n754), .B1(new_n561), .B2(new_n616), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n657), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n752), .B1(new_n759), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n751), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G122), .ZN(G24));
  OAI211_X1 g581(.A(new_n678), .B(new_n748), .C1(new_n749), .C2(new_n705), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n743), .A2(new_n689), .A3(new_n720), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G125), .ZN(G27));
  NAND3_X1  g586(.A1(new_n655), .A2(new_n333), .A3(new_n656), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n773), .A2(new_n720), .A3(new_n699), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n312), .A2(new_n325), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT32), .B1(new_n710), .B2(new_n187), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n472), .B(new_n774), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT42), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n330), .A2(KEYINPUT42), .A3(new_n472), .A4(new_n774), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G131), .ZN(G33));
  NOR3_X1   g596(.A1(new_n773), .A2(new_n695), .A3(new_n699), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n472), .B(new_n783), .C1(new_n775), .C2(new_n776), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G134), .ZN(G36));
  NAND2_X1  g599(.A1(new_n645), .A2(new_n703), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n637), .A2(new_n617), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT43), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n786), .A2(new_n678), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT113), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n789), .A2(new_n678), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n673), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n795), .A3(KEYINPUT44), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n422), .A2(new_n423), .A3(new_n332), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(new_n794), .B2(KEYINPUT44), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n496), .A2(new_n488), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n502), .A2(new_n494), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT45), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n476), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n503), .A2(KEYINPUT45), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n477), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n807), .A2(KEYINPUT46), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n509), .B1(new_n807), .B2(KEYINPUT46), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n474), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n700), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n797), .A2(new_n800), .A3(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G137), .ZN(G39));
  XOR2_X1   g627(.A(new_n810), .B(KEYINPUT47), .Z(new_n814));
  NOR4_X1   g628(.A1(new_n330), .A2(new_n472), .A3(new_n720), .A4(new_n773), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  INV_X1    g631(.A(new_n472), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n818), .A2(new_n787), .A3(new_n475), .A4(new_n332), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n731), .B(KEYINPUT49), .Z(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OR3_X1    g635(.A1(new_n821), .A2(new_n712), .A3(new_n714), .ZN(new_n822));
  INV_X1    g636(.A(new_n712), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n798), .A2(new_n732), .A3(new_n733), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n824), .A2(new_n818), .A3(new_n336), .ZN(new_n825));
  INV_X1    g639(.A(new_n637), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n823), .A2(new_n825), .A3(new_n617), .A4(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n827), .B(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n810), .B(KEYINPUT47), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n731), .A2(new_n474), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n773), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n336), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n789), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n750), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n824), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n833), .A2(new_n836), .B1(new_n769), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT50), .ZN(new_n839));
  AOI211_X1 g653(.A(new_n333), .B(new_n714), .C1(KEYINPUT116), .C2(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n835), .A2(new_n743), .A3(new_n750), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n842), .A2(new_n843), .A3(KEYINPUT50), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n840), .B(new_n841), .C1(KEYINPUT116), .C2(new_n839), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n829), .A2(new_n838), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT51), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n841), .A2(new_n657), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n818), .B1(new_n704), .B2(new_n735), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n837), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT48), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n277), .A2(G952), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT119), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n823), .B(new_n825), .C1(new_n638), .C2(new_n633), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n849), .A2(new_n852), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT118), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n846), .A2(new_n857), .A3(new_n847), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n857), .B1(new_n846), .B2(new_n847), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n848), .B(new_n856), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n769), .A2(new_n770), .B1(new_n330), .B2(new_n696), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n759), .A2(new_n764), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n699), .A2(new_n678), .A3(new_n693), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n712), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n725), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n724), .B1(new_n330), .B2(new_n721), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n862), .B(new_n865), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n726), .A2(KEYINPUT52), .A3(new_n862), .A4(new_n865), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n645), .A2(new_n774), .A3(new_n678), .A4(new_n748), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n662), .A2(new_n562), .A3(new_n663), .A4(new_n694), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n690), .A2(new_n773), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n875), .B1(new_n775), .B2(new_n776), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n784), .A2(new_n873), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n736), .B1(new_n643), .B2(new_n669), .ZN(new_n878));
  AOI22_X1  g692(.A1(new_n683), .A2(new_n744), .B1(new_n751), .B2(new_n765), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n781), .A2(new_n877), .A3(new_n878), .A4(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n826), .A2(new_n617), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n645), .A2(new_n646), .A3(new_n641), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n620), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT114), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT114), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n620), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n562), .A2(new_n616), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n645), .A2(new_n646), .A3(new_n641), .A4(new_n887), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n684), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n884), .A2(new_n886), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n880), .A2(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n872), .A2(new_n891), .A3(KEYINPUT53), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT53), .B1(new_n872), .B2(new_n891), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT54), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n872), .A2(new_n891), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT53), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n872), .A2(new_n891), .A3(KEYINPUT53), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n894), .A2(new_n900), .A3(KEYINPUT115), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT115), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n897), .A2(new_n902), .A3(new_n898), .A4(new_n899), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n861), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(G952), .A2(G953), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n822), .B1(new_n904), .B2(new_n905), .ZN(G75));
  XNOR2_X1  g720(.A(new_n419), .B(new_n420), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT55), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n323), .B1(new_n897), .B2(new_n899), .ZN(new_n909));
  AOI211_X1 g723(.A(KEYINPUT56), .B(new_n908), .C1(new_n909), .C2(G210), .ZN(new_n910));
  INV_X1    g724(.A(new_n908), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n897), .A2(new_n899), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n912), .A2(G210), .A3(G902), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT56), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n277), .A2(G952), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n910), .A2(new_n915), .A3(new_n916), .ZN(G51));
  XNOR2_X1  g731(.A(new_n477), .B(KEYINPUT57), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT54), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n898), .B1(new_n897), .B2(new_n899), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n507), .A2(new_n508), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n909), .A2(new_n806), .A3(new_n805), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n916), .B1(new_n923), .B2(new_n924), .ZN(G54));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n926));
  AND2_X1   g740(.A1(KEYINPUT58), .A2(G475), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n909), .A2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n614), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n916), .B1(new_n928), .B2(new_n929), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n909), .A2(KEYINPUT120), .A3(new_n614), .A4(new_n927), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(G60));
  NAND2_X1  g747(.A1(new_n626), .A2(new_n627), .ZN(new_n934));
  NAND2_X1  g748(.A1(G478), .A2(G902), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT59), .Z(new_n936));
  NOR2_X1   g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n919), .B2(new_n920), .ZN(new_n938));
  INV_X1    g752(.A(new_n916), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n936), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n901), .A2(new_n903), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n940), .B1(new_n934), .B2(new_n942), .ZN(G63));
  NAND2_X1  g757(.A1(G217), .A2(G902), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT60), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n676), .B(new_n946), .C1(new_n892), .C2(new_n893), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n945), .B1(new_n897), .B2(new_n899), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n947), .B(new_n939), .C1(new_n948), .C2(new_n461), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(G66));
  NAND2_X1  g765(.A1(new_n878), .A2(new_n879), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n890), .A2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT121), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n953), .A2(new_n954), .A3(new_n277), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n890), .A2(new_n952), .ZN(new_n956));
  OAI21_X1  g770(.A(KEYINPUT121), .B1(new_n956), .B2(G953), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT122), .ZN(new_n959));
  OAI21_X1  g773(.A(G953), .B1(new_n391), .B2(new_n338), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n959), .B1(new_n958), .B2(new_n960), .ZN(new_n962));
  INV_X1    g776(.A(G898), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n419), .B1(new_n963), .B2(G953), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  OR3_X1    g779(.A1(new_n961), .A2(new_n962), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n965), .B1(new_n961), .B2(new_n962), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(G69));
  OAI21_X1  g782(.A(G953), .B1(new_n492), .B2(new_n691), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT126), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n244), .A2(new_n256), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n602), .A2(new_n603), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT123), .Z(new_n973));
  XOR2_X1   g787(.A(new_n971), .B(new_n973), .Z(new_n974));
  AND2_X1   g788(.A1(new_n726), .A2(new_n862), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n975), .A2(KEYINPUT62), .A3(new_n717), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n726), .A2(new_n717), .A3(new_n862), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT62), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI22_X1  g793(.A1(new_n976), .A2(new_n979), .B1(new_n814), .B2(new_n815), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n881), .A2(new_n887), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT124), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n982), .A2(new_n701), .A3(new_n850), .A4(new_n798), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n812), .A2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT125), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(KEYINPUT125), .B1(new_n812), .B2(new_n983), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n980), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n974), .B1(new_n988), .B2(new_n277), .ZN(new_n989));
  AND4_X1   g803(.A1(new_n781), .A2(new_n975), .A3(new_n784), .A4(new_n816), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n799), .B1(new_n792), .B2(new_n796), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n850), .A2(new_n863), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n811), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(G953), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n277), .A2(G900), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n974), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n970), .B1(new_n989), .B2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n970), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n984), .B(new_n985), .ZN(new_n1000));
  AOI21_X1  g814(.A(G953), .B1(new_n1000), .B2(new_n980), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n999), .B(new_n996), .C1(new_n1001), .C2(new_n974), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n998), .A2(new_n1002), .ZN(G72));
  NAND3_X1  g817(.A1(new_n990), .A2(new_n956), .A3(new_n993), .ZN(new_n1004));
  NAND2_X1  g818(.A1(G472), .A2(G902), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT63), .Z(new_n1006));
  NAND2_X1  g820(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n1007), .A2(new_n320), .A3(new_n275), .A4(new_n273), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1006), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n319), .A2(new_n320), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1009), .B1(new_n706), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n912), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1008), .A2(new_n939), .A3(new_n1012), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n980), .B(new_n956), .C1(new_n986), .C2(new_n987), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT127), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1014), .A2(new_n1015), .A3(new_n1006), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n1016), .A2(new_n286), .A3(new_n319), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1014), .ZN(new_n1018));
  OAI21_X1  g832(.A(KEYINPUT127), .B1(new_n1018), .B2(new_n1009), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1013), .B1(new_n1017), .B2(new_n1019), .ZN(G57));
endmodule


