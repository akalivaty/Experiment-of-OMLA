//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI21_X1  g0005(.A(G50), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT65), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G77), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n211), .B1(new_n203), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n202), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n210), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT66), .Z(new_n222));
  INV_X1    g0022(.A(KEYINPUT1), .ZN(new_n223));
  AND2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n222), .A2(new_n223), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n204), .A2(new_n205), .ZN(new_n226));
  INV_X1    g0026(.A(G50), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AND2_X1   g0031(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n210), .A2(G13), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n233), .B(G250), .C1(G257), .C2(G264), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT0), .Z(new_n235));
  NOR4_X1   g0035(.A1(new_n224), .A2(new_n225), .A3(new_n232), .A4(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n217), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT67), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  AOI21_X1  g0052(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G77), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n254), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  MUX2_X1   g0061(.A(G222), .B(G223), .S(G1698), .Z(new_n262));
  OAI21_X1  g0062(.A(new_n261), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n253), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT68), .B(G45), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n265), .B(new_n266), .C1(G41), .C2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G226), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(KEYINPUT69), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT69), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G1), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(G41), .B2(G45), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n254), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n263), .B(new_n268), .C1(new_n269), .C2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G169), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(G179), .B2(new_n276), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n229), .B1(new_n210), .B2(new_n258), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT70), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OR3_X1    g0084(.A1(new_n283), .A2(new_n202), .A3(KEYINPUT8), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n230), .A2(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n288), .B1(G150), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n207), .A2(G20), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n281), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n273), .A2(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(new_n280), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G50), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n270), .A2(new_n272), .A3(G13), .A4(G20), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n296), .B1(G50), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n279), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT10), .ZN(new_n301));
  OR3_X1    g0101(.A1(new_n292), .A2(KEYINPUT9), .A3(new_n298), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT9), .B1(new_n292), .B2(new_n298), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n276), .A2(G200), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(new_n276), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n301), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n304), .A2(new_n301), .A3(new_n308), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n300), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n274), .A2(G244), .A3(new_n254), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n313), .A2(new_n268), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n257), .A2(new_n259), .ZN(new_n315));
  INV_X1    g0115(.A(G1698), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(G232), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G107), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(new_n315), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n260), .A2(new_n212), .A3(new_n316), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n253), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n314), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G190), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n297), .A2(new_n281), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT71), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n297), .A2(new_n281), .A3(KEYINPUT71), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n327), .A2(new_n293), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G77), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G20), .A2(G77), .ZN(new_n331));
  INV_X1    g0131(.A(new_n289), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT15), .B(G87), .ZN(new_n333));
  OAI221_X1 g0133(.A(new_n331), .B1(new_n282), .B2(new_n332), .C1(new_n287), .C2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n297), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n334), .A2(new_n280), .B1(new_n255), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n322), .A2(G200), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n324), .A2(new_n330), .A3(new_n336), .A4(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n322), .A2(new_n277), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n330), .A2(new_n336), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n339), .B(new_n340), .C1(G179), .C2(new_n322), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n312), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT80), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n286), .A2(new_n297), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n295), .B2(new_n286), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT16), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT7), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n315), .B2(G20), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n260), .A2(KEYINPUT7), .A3(new_n230), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n203), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n202), .A2(new_n203), .ZN(new_n353));
  OAI21_X1  g0153(.A(G20), .B1(new_n226), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n289), .A2(G159), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n348), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT77), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n358), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n281), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n354), .A2(new_n355), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT75), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n258), .B2(KEYINPUT3), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n256), .A2(KEYINPUT75), .A3(G33), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(new_n365), .A3(new_n259), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n349), .B1(new_n366), .B2(new_n230), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n349), .A3(new_n230), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G68), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n362), .B(KEYINPUT16), .C1(new_n367), .C2(new_n369), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n370), .B(KEYINPUT76), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n347), .B1(new_n361), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n274), .A2(G232), .A3(new_n254), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n268), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT79), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n373), .A2(KEYINPUT79), .A3(new_n268), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(new_n306), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n269), .A2(G1698), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(G223), .B2(G1698), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n366), .A2(new_n380), .B1(new_n258), .B2(new_n213), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n253), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n382), .B(KEYINPUT78), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n374), .B1(new_n253), .B2(new_n381), .ZN(new_n384));
  OAI22_X1  g0184(.A1(new_n378), .A2(new_n383), .B1(new_n384), .B2(G200), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n372), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT17), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n361), .A2(new_n371), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n346), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT18), .ZN(new_n391));
  INV_X1    g0191(.A(G179), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n376), .A2(new_n392), .A3(new_n377), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n393), .A2(new_n383), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n384), .A2(G169), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n390), .A2(new_n391), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n396), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT18), .B1(new_n372), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n372), .A2(KEYINPUT17), .A3(new_n385), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n388), .A2(new_n397), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n332), .A2(new_n227), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n287), .A2(new_n255), .B1(new_n230), .B2(G68), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n280), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT73), .ZN(new_n406));
  OR2_X1    g0206(.A1(new_n406), .A2(KEYINPUT11), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(KEYINPUT11), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n329), .A2(G68), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n335), .A2(new_n203), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT12), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n407), .A2(new_n408), .A3(new_n409), .A4(new_n411), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n412), .B(KEYINPUT74), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n268), .B1(new_n275), .B2(new_n212), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n217), .A2(G1698), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n315), .B(new_n415), .C1(G226), .C2(G1698), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G97), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n254), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OR2_X1    g0218(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT13), .ZN(new_n420));
  OR3_X1    g0220(.A1(new_n414), .A2(KEYINPUT13), .A3(new_n418), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(G190), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT72), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n420), .A2(new_n423), .A3(new_n421), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n419), .A2(KEYINPUT72), .A3(KEYINPUT13), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(G200), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n413), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n413), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n424), .A2(G169), .A3(new_n425), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT14), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT14), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n424), .A2(new_n432), .A3(G169), .A4(new_n425), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n420), .A2(G179), .A3(new_n421), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n428), .B1(new_n429), .B2(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n343), .A2(new_n344), .A3(new_n402), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n429), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n312), .A2(new_n427), .A3(new_n438), .A4(new_n342), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT80), .B1(new_n439), .B2(new_n401), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n364), .A2(new_n365), .A3(new_n259), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n442), .A2(KEYINPUT22), .A3(new_n230), .A4(G87), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT23), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(new_n318), .A3(G20), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT87), .ZN(new_n446));
  INV_X1    g0246(.A(G116), .ZN(new_n447));
  OAI22_X1  g0247(.A1(new_n445), .A2(new_n446), .B1(new_n287), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(new_n446), .B2(new_n445), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT23), .B1(new_n230), .B2(G107), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT86), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT22), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n230), .A2(G87), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n453), .B1(new_n260), .B2(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n443), .A2(new_n449), .A3(new_n452), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT24), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n452), .A2(new_n455), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT24), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n458), .A2(new_n459), .A3(new_n443), .A4(new_n449), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n281), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n270), .A2(new_n272), .A3(G33), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n297), .A2(new_n281), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G107), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n335), .A2(KEYINPUT25), .A3(new_n318), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT25), .B1(new_n335), .B2(new_n318), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n219), .A2(G1698), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(G250), .B2(G1698), .ZN(new_n470));
  INV_X1    g0270(.A(G294), .ZN(new_n471));
  OAI22_X1  g0271(.A1(new_n366), .A2(new_n470), .B1(new_n258), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n253), .ZN(new_n473));
  XOR2_X1   g0273(.A(KEYINPUT5), .B(G41), .Z(new_n474));
  NAND3_X1  g0274(.A1(new_n270), .A2(new_n272), .A3(G45), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n265), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n254), .B(G264), .C1(new_n474), .C2(new_n475), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n473), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G200), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(new_n306), .B2(new_n479), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n468), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT88), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT88), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n468), .A2(new_n485), .A3(new_n482), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n318), .B1(new_n350), .B2(new_n351), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT6), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n489), .A2(new_n218), .A3(G107), .ZN(new_n490));
  XNOR2_X1  g0290(.A(G97), .B(G107), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n490), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  OAI22_X1  g0292(.A1(new_n492), .A2(new_n230), .B1(new_n255), .B2(new_n332), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n280), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n463), .A2(G97), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n335), .A2(new_n218), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n257), .A2(new_n259), .A3(G250), .A4(G1698), .ZN(new_n500));
  AND2_X1   g0300(.A1(KEYINPUT4), .A2(G244), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n257), .A2(new_n259), .A3(new_n501), .A4(new_n316), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G283), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT4), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n364), .A2(new_n365), .A3(G244), .A4(new_n259), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n505), .B1(new_n506), .B2(G1698), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n254), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n254), .B(G257), .C1(new_n474), .C2(new_n475), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n477), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G190), .ZN(new_n512));
  INV_X1    g0312(.A(G200), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n499), .B(new_n512), .C1(new_n513), .C2(new_n511), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n392), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n277), .B1(new_n508), .B2(new_n510), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n498), .A3(new_n516), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n479), .A2(new_n277), .ZN(new_n519));
  OAI221_X1 g0319(.A(new_n519), .B1(G179), .B2(new_n479), .C1(new_n461), .C2(new_n467), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n487), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n254), .B(G270), .C1(new_n474), .C2(new_n475), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n477), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G264), .A2(G1698), .ZN(new_n524));
  INV_X1    g0324(.A(G303), .ZN(new_n525));
  OAI22_X1  g0325(.A1(new_n366), .A2(new_n524), .B1(new_n315), .B2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n442), .A2(KEYINPUT84), .A3(G257), .A4(new_n316), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT84), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n316), .A2(G257), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n366), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n526), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n523), .B1(new_n531), .B2(new_n254), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n327), .A2(G116), .A3(new_n328), .A4(new_n462), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n503), .B(new_n230), .C1(G33), .C2(new_n218), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n447), .A2(G20), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n534), .A2(new_n280), .A3(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT20), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n534), .A2(new_n280), .A3(KEYINPUT20), .A4(new_n535), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n538), .A2(new_n539), .B1(new_n447), .B2(new_n335), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n277), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n532), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT21), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT85), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT85), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n532), .A2(new_n541), .A3(new_n545), .A4(KEYINPUT21), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n533), .A2(new_n540), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n548), .A2(G179), .A3(new_n523), .ZN(new_n549));
  OR2_X1    g0349(.A1(new_n531), .A2(new_n254), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n549), .A2(new_n550), .B1(new_n542), .B2(new_n543), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n548), .B1(new_n532), .B2(G200), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n306), .B2(new_n532), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n547), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n203), .A2(G20), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n364), .A2(new_n365), .A3(new_n555), .A4(new_n259), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n230), .B1(new_n417), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n213), .A2(new_n218), .A3(new_n318), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n557), .B1(new_n287), .B2(new_n218), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n556), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n280), .ZN(new_n563));
  INV_X1    g0363(.A(new_n333), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n564), .A2(new_n297), .A3(new_n281), .A4(new_n462), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n564), .A2(new_n297), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n563), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT83), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n566), .B1(new_n562), .B2(new_n280), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(KEYINPUT83), .A3(new_n565), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  OR2_X1    g0373(.A1(new_n214), .A2(KEYINPUT81), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n475), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(G274), .B1(KEYINPUT81), .B2(G250), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n270), .A2(new_n576), .A3(new_n272), .A4(G45), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n254), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT82), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n442), .A2(new_n580), .A3(G244), .A4(G1698), .ZN(new_n581));
  OAI21_X1  g0381(.A(KEYINPUT82), .B1(new_n506), .B2(new_n316), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n212), .A2(G1698), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n364), .A2(new_n365), .A3(new_n583), .A4(new_n259), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G33), .A2(G116), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n581), .A2(new_n582), .A3(new_n586), .ZN(new_n587));
  AOI211_X1 g0387(.A(G179), .B(new_n579), .C1(new_n587), .C2(new_n253), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n573), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n253), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n578), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n277), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(G200), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n463), .A2(G87), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n571), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n579), .B1(new_n587), .B2(new_n253), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n595), .B1(new_n596), .B2(G190), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n589), .A2(new_n592), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n521), .A2(new_n554), .A3(new_n599), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n441), .A2(new_n600), .ZN(G372));
  NAND3_X1  g0401(.A1(new_n590), .A2(new_n392), .A3(new_n578), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n592), .A2(new_n602), .A3(new_n572), .A4(new_n570), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n515), .A2(new_n498), .A3(new_n516), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n593), .A2(new_n597), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n603), .A2(KEYINPUT26), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT92), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT92), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n598), .A2(new_n608), .A3(KEYINPUT26), .A4(new_n604), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n590), .A2(KEYINPUT89), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT89), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n587), .A2(new_n612), .A3(new_n253), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n579), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n589), .B1(new_n614), .B2(G169), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n597), .B1(new_n614), .B2(new_n513), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT90), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n617), .B1(new_n615), .B2(new_n616), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n604), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT26), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n610), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n602), .A2(new_n572), .A3(new_n570), .ZN(new_n623));
  INV_X1    g0423(.A(new_n613), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n612), .B1(new_n587), .B2(new_n253), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n578), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n623), .B1(new_n277), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(KEYINPUT93), .B1(new_n622), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n607), .A2(new_n609), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n590), .A2(G190), .A3(new_n578), .ZN(new_n630));
  INV_X1    g0430(.A(new_n595), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n626), .B2(G200), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT90), .B1(new_n627), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n517), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n629), .B1(new_n636), .B2(KEYINPUT26), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT93), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(new_n638), .A3(new_n615), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n485), .B1(new_n468), .B2(new_n482), .ZN(new_n640));
  NOR4_X1   g0440(.A1(new_n481), .A2(new_n461), .A3(KEYINPUT88), .A4(new_n467), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n518), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n547), .A2(new_n520), .A3(new_n551), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT91), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n634), .A2(new_n635), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n487), .A2(new_n518), .A3(new_n643), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n618), .A2(new_n619), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT91), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n628), .A2(new_n639), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n441), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n397), .A2(new_n399), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n388), .A2(new_n400), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(new_n428), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n438), .A2(new_n341), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n310), .A2(new_n311), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n300), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n654), .A2(new_n662), .ZN(G369));
  NAND2_X1  g0463(.A1(new_n547), .A2(new_n551), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n230), .A2(G13), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n273), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G343), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n670), .B1(new_n533), .B2(new_n540), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n554), .A2(new_n671), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n672), .A2(new_n673), .A3(KEYINPUT94), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(KEYINPUT94), .B2(new_n672), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  INV_X1    g0476(.A(new_n520), .ZN(new_n677));
  INV_X1    g0477(.A(new_n670), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n461), .B2(new_n467), .ZN(new_n679));
  XOR2_X1   g0479(.A(new_n679), .B(KEYINPUT95), .Z(new_n680));
  AOI21_X1  g0480(.A(new_n677), .B1(new_n680), .B2(new_n487), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n520), .A2(new_n678), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n676), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n680), .A2(new_n487), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n520), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n664), .A2(new_n670), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n682), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n686), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n233), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n559), .A2(G116), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G1), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n228), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n697), .B1(new_n698), .B2(new_n695), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT28), .ZN(new_n700));
  INV_X1    g0500(.A(G330), .ZN(new_n701));
  NOR4_X1   g0501(.A1(new_n521), .A2(new_n554), .A3(new_n599), .A4(new_n678), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT31), .ZN(new_n703));
  AND4_X1   g0503(.A1(G179), .A2(new_n523), .A3(new_n478), .A4(new_n473), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n704), .A2(new_n550), .A3(new_n596), .A4(new_n511), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT30), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(KEYINPUT30), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n479), .A2(new_n392), .ZN(new_n708));
  AOI211_X1 g0508(.A(new_n511), .B(new_n708), .C1(new_n550), .C2(new_n523), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n706), .A2(new_n707), .B1(new_n626), .B2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT96), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n678), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n705), .B(KEYINPUT30), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n709), .A2(new_n626), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n713), .A2(new_n711), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n703), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n710), .A2(new_n703), .A3(new_n670), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT97), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n702), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n716), .A2(KEYINPUT97), .A3(new_n718), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n701), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT98), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n637), .A2(new_n615), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n725), .A2(KEYINPUT93), .B1(new_n651), .B2(new_n648), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n678), .B1(new_n726), .B2(new_n639), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n724), .B1(new_n727), .B2(KEYINPUT29), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n653), .A2(new_n670), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT29), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n729), .A2(KEYINPUT98), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n599), .A2(KEYINPUT26), .A3(new_n517), .ZN(new_n733));
  AOI211_X1 g0533(.A(new_n627), .B(new_n733), .C1(new_n645), .C2(new_n647), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n620), .A2(KEYINPUT26), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n678), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(KEYINPUT29), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n723), .B1(new_n732), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n700), .B1(new_n738), .B2(G1), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT99), .ZN(G364));
  AOI21_X1  g0540(.A(new_n266), .B1(new_n665), .B2(G45), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n694), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n743), .B1(new_n675), .B2(G330), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n675), .A2(G330), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G13), .A2(G33), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n675), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n743), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n229), .B1(G20), .B2(new_n277), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n230), .A2(new_n392), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G190), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n315), .B1(new_n757), .B2(new_n255), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n755), .A2(G190), .A3(new_n513), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n758), .B1(G58), .B2(new_n760), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n306), .A2(G179), .A3(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n230), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n755), .A2(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n306), .ZN(new_n766));
  AOI22_X1  g0566(.A1(G97), .A2(new_n764), .B1(new_n766), .B2(G50), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n230), .A2(G179), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n756), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G159), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n768), .A2(new_n306), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n771), .A2(KEYINPUT32), .B1(G107), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n761), .A2(new_n767), .A3(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n768), .A2(G190), .A3(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n213), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n765), .A2(G190), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n778), .B1(new_n771), .B2(KEYINPUT32), .C1(new_n780), .C2(new_n203), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n775), .A2(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n760), .A2(G322), .B1(new_n770), .B2(G329), .ZN(new_n783));
  INV_X1    g0583(.A(new_n757), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n315), .B1(new_n784), .B2(G311), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n766), .A2(G326), .ZN(new_n787));
  XNOR2_X1  g0587(.A(KEYINPUT33), .B(G317), .ZN(new_n788));
  INV_X1    g0588(.A(new_n776), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n779), .A2(new_n788), .B1(new_n789), .B2(G303), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n764), .A2(G294), .B1(new_n773), .B2(G283), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n786), .A2(new_n787), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n754), .B1(new_n782), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n749), .A2(new_n753), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n693), .A2(new_n260), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n795), .A2(G355), .B1(new_n447), .B2(new_n693), .ZN(new_n796));
  INV_X1    g0596(.A(G45), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n248), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n442), .A2(new_n693), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n698), .B2(new_n267), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n796), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n752), .B(new_n793), .C1(new_n794), .C2(new_n801), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n744), .A2(new_n746), .B1(new_n751), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(G396));
  NAND2_X1  g0604(.A1(new_n678), .A2(new_n340), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n338), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n341), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n341), .A2(new_n678), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n748), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n766), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n813), .A2(new_n525), .B1(new_n772), .B2(new_n213), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G97), .A2(new_n764), .B1(new_n779), .B2(G283), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n315), .B1(new_n770), .B2(G311), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n760), .A2(G294), .B1(new_n784), .B2(G116), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n814), .B(new_n818), .C1(G107), .C2(new_n789), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT100), .Z(new_n820));
  AOI22_X1  g0620(.A1(G137), .A2(new_n766), .B1(new_n779), .B2(G150), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT101), .ZN(new_n822));
  INV_X1    g0622(.A(G143), .ZN(new_n823));
  INV_X1    g0623(.A(G159), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n822), .B1(new_n823), .B2(new_n759), .C1(new_n824), .C2(new_n757), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT34), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G132), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n442), .B1(new_n828), .B2(new_n769), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n763), .A2(new_n202), .B1(new_n776), .B2(new_n227), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n772), .A2(new_n203), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n825), .B2(new_n826), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n820), .B1(new_n827), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n753), .A2(new_n747), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n834), .A2(new_n753), .B1(new_n255), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n752), .B1(new_n812), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n729), .A2(new_n809), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n653), .A2(new_n670), .A3(new_n810), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(new_n723), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n838), .B1(new_n842), .B2(new_n743), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT102), .Z(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(G384));
  INV_X1    g0645(.A(new_n492), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n846), .A2(KEYINPUT35), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(KEYINPUT35), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n847), .A2(G116), .A3(new_n231), .A4(new_n848), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT36), .Z(new_n850));
  OAI211_X1 g0650(.A(new_n228), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n227), .A2(G68), .ZN(new_n852));
  AOI211_X1 g0652(.A(G13), .B(new_n273), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n662), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n737), .A2(new_n441), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT98), .B1(new_n729), .B2(new_n730), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n724), .B(KEYINPUT29), .C1(new_n653), .C2(new_n670), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT107), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT107), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n857), .B(new_n862), .C1(new_n858), .C2(new_n859), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n855), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n362), .B1(new_n367), .B2(new_n369), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n281), .B1(new_n865), .B2(new_n348), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n371), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n346), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n669), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n401), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n868), .A2(new_n396), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n386), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT104), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n390), .A2(new_n875), .A3(new_n396), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT104), .B1(new_n372), .B2(new_n398), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n390), .A2(new_n669), .ZN(new_n878));
  XOR2_X1   g0678(.A(KEYINPUT105), .B(KEYINPUT37), .Z(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n372), .B2(new_n385), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n876), .A2(new_n877), .A3(new_n878), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n874), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n871), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n871), .A2(new_n882), .A3(KEYINPUT38), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n386), .B1(new_n372), .B2(new_n398), .ZN(new_n887));
  INV_X1    g0687(.A(new_n669), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n372), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n879), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n881), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n401), .A2(new_n889), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT38), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT106), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n885), .B(new_n886), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT39), .ZN(new_n896));
  INV_X1    g0696(.A(new_n886), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n897), .A2(new_n893), .ZN(new_n898));
  NOR2_X1   g0698(.A1(KEYINPUT106), .A2(KEYINPUT39), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n438), .A2(new_n678), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n901), .A2(new_n902), .B1(new_n655), .B2(new_n888), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n438), .B(new_n427), .C1(new_n413), .C2(new_n670), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n429), .B(new_n678), .C1(new_n428), .C2(new_n435), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n808), .B(KEYINPUT103), .Z(new_n908));
  AOI21_X1  g0708(.A(new_n907), .B1(new_n840), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n885), .A2(new_n886), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n903), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n864), .B(new_n912), .Z(new_n913));
  INV_X1    g0713(.A(new_n702), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n713), .A2(new_n714), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n670), .B1(new_n915), .B2(KEYINPUT96), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n710), .A2(new_n711), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n916), .A2(KEYINPUT31), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n914), .A2(new_n716), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n809), .B1(new_n904), .B2(new_n905), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n919), .B(new_n920), .C1(new_n897), .C2(new_n893), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT40), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n919), .A2(new_n920), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT40), .B1(new_n885), .B2(new_n886), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n441), .A2(new_n919), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n701), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n927), .B2(new_n926), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n913), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n273), .B2(new_n665), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n913), .A2(new_n929), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n854), .B1(new_n931), .B2(new_n932), .ZN(G367));
  INV_X1    g0733(.A(new_n799), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n794), .B1(new_n233), .B2(new_n333), .C1(new_n934), .C2(new_n243), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n935), .A2(new_n743), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n780), .A2(new_n471), .B1(new_n772), .B2(new_n218), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(G311), .B2(new_n766), .ZN(new_n938));
  INV_X1    g0738(.A(G283), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n763), .A2(new_n318), .B1(new_n757), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT115), .ZN(new_n941));
  INV_X1    g0741(.A(G317), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n759), .A2(new_n525), .B1(new_n769), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT46), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n776), .A2(new_n944), .A3(new_n447), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n943), .A2(new_n945), .A3(new_n442), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n944), .B1(new_n776), .B2(new_n447), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT116), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n938), .A2(new_n941), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n763), .A2(new_n203), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(G150), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n951), .B1(new_n759), .B2(new_n952), .C1(new_n823), .C2(new_n813), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT117), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n260), .B1(new_n784), .B2(G50), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n773), .A2(G77), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n955), .B(new_n956), .C1(new_n780), .C2(new_n824), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT118), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n789), .A2(G58), .B1(new_n770), .B2(G137), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n958), .B2(new_n959), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n949), .B1(new_n954), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT47), .Z(new_n963));
  NOR2_X1   g0763(.A1(new_n670), .A2(new_n631), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n615), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n647), .B2(new_n964), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT108), .Z(new_n967));
  OAI221_X1 g0767(.A(new_n936), .B1(new_n754), .B2(new_n963), .C1(new_n967), .C2(new_n750), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT112), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n514), .A2(new_n517), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n499), .A2(new_n670), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n970), .A2(new_n971), .B1(new_n517), .B2(new_n670), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT109), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n691), .A2(new_n969), .A3(new_n973), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n681), .A2(new_n689), .B1(new_n520), .B2(new_n678), .ZN(new_n975));
  INV_X1    g0775(.A(new_n973), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT112), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT45), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n977), .A2(new_n974), .A3(KEYINPUT45), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT44), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n691), .B2(new_n973), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n975), .A2(new_n976), .A3(KEYINPUT44), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n980), .A2(KEYINPUT113), .A3(new_n981), .A4(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT114), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n978), .A2(new_n979), .B1(new_n984), .B2(new_n983), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n981), .ZN(new_n990));
  OAI21_X1  g0790(.A(KEYINPUT113), .B1(new_n685), .B2(KEYINPUT114), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n988), .A2(new_n685), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n683), .B(new_n689), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(new_n676), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n738), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n694), .B(KEYINPUT41), .Z(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n742), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(KEYINPUT111), .B1(new_n686), .B2(new_n976), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT111), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n685), .A2(new_n1003), .A3(new_n973), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1000), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n683), .A2(new_n690), .A3(new_n973), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT42), .Z(new_n1008));
  AOI21_X1  g0808(.A(new_n604), .B1(new_n973), .B2(new_n677), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n678), .B1(new_n1009), .B2(KEYINPUT110), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(KEYINPUT110), .B2(new_n1009), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1002), .B1(new_n1000), .B2(new_n1004), .ZN(new_n1015));
  OR3_X1    g0815(.A1(new_n1006), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1014), .B1(new_n1006), .B2(new_n1015), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n968), .B1(new_n999), .B2(new_n1018), .ZN(G387));
  AOI21_X1  g0819(.A(new_n695), .B1(new_n738), .B2(new_n994), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n738), .B2(new_n994), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n240), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n934), .B1(new_n1022), .B2(new_n267), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n696), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1023), .B1(new_n1024), .B2(new_n795), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n282), .A2(G50), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT50), .Z(new_n1027));
  OAI21_X1  g0827(.A(new_n797), .B1(new_n203), .B2(new_n255), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n1027), .A2(new_n1024), .A3(new_n1028), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n1025), .A2(new_n1029), .B1(G107), .B2(new_n233), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n752), .B1(new_n1030), .B2(new_n794), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n763), .A2(new_n333), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n255), .B2(new_n776), .C1(new_n824), .C2(new_n813), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n760), .A2(G50), .B1(new_n770), .B2(G150), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n366), .B1(new_n773), .B2(G97), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1035), .B(new_n1036), .C1(new_n203), .C2(new_n757), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n780), .A2(new_n286), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n1034), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n764), .A2(G283), .B1(new_n789), .B2(G294), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n759), .A2(new_n942), .B1(new_n757), .B2(new_n525), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT119), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G311), .A2(new_n779), .B1(new_n766), .B2(G322), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n1042), .B2(new_n1041), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT48), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1040), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT120), .Z(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n1048), .B2(new_n1047), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1051), .A2(KEYINPUT49), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n442), .B1(G326), .B2(new_n770), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n447), .B2(new_n772), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n1051), .B2(KEYINPUT49), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1039), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1031), .B1(new_n1056), .B2(new_n754), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n684), .B2(new_n749), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n994), .B2(new_n742), .ZN(new_n1059));
  AOI21_X1  g0859(.A(KEYINPUT121), .B1(new_n1021), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1021), .A2(KEYINPUT121), .A3(new_n1059), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(G393));
  NAND2_X1  g0863(.A1(new_n738), .A2(new_n994), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT122), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n989), .A2(new_n685), .A3(new_n1065), .A4(new_n981), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n686), .A2(KEYINPUT122), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n685), .A2(new_n1065), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n990), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1064), .A2(new_n1066), .A3(new_n1069), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1070), .B(new_n694), .C1(new_n1064), .C2(new_n992), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1066), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT123), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n741), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1069), .A2(KEYINPUT123), .A3(new_n1066), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n976), .A2(new_n749), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n794), .B1(new_n218), .B2(new_n233), .C1(new_n934), .C2(new_n251), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n743), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G317), .A2(new_n766), .B1(new_n760), .B2(G311), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT52), .Z(new_n1080));
  NOR2_X1   g0880(.A1(new_n757), .A2(new_n471), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n315), .B(new_n1081), .C1(G322), .C2(new_n770), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n779), .A2(G303), .B1(new_n773), .B2(G107), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n764), .A2(G116), .B1(new_n789), .B2(G283), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1080), .A2(new_n1082), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT124), .Z(new_n1086));
  OAI22_X1  g0886(.A1(new_n813), .A2(new_n952), .B1(new_n824), .B2(new_n759), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT51), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n757), .A2(new_n282), .B1(new_n769), .B2(new_n823), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1089), .A2(new_n366), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n763), .A2(new_n255), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n203), .A2(new_n776), .B1(new_n772), .B2(new_n213), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1091), .B(new_n1092), .C1(G50), .C2(new_n779), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1088), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1086), .A2(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT125), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1078), .B1(new_n1096), .B2(new_n753), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1074), .A2(new_n1075), .B1(new_n1076), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1071), .A2(new_n1098), .ZN(G390));
  AOI21_X1  g0899(.A(new_n752), .B1(new_n286), .B2(new_n835), .ZN(new_n1100));
  INV_X1    g0900(.A(G128), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n813), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n779), .A2(G137), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n227), .B2(new_n772), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1102), .B(new_n1104), .C1(G159), .C2(new_n764), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n776), .A2(new_n952), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT53), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(KEYINPUT54), .B(G143), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n759), .A2(new_n828), .B1(new_n757), .B2(new_n1108), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n260), .B(new_n1109), .C1(G125), .C2(new_n770), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1105), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1091), .B1(G283), .B2(new_n766), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n759), .A2(new_n447), .B1(new_n769), .B2(new_n471), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n260), .B1(new_n757), .B2(new_n218), .ZN(new_n1114));
  NOR4_X1   g0914(.A1(new_n1113), .A2(new_n1114), .A3(new_n777), .A4(new_n831), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1112), .B(new_n1115), .C1(new_n318), .C2(new_n780), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1100), .B1(new_n754), .B2(new_n1117), .C1(new_n901), .C2(new_n748), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n895), .A2(KEYINPUT39), .B1(new_n898), .B2(new_n899), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n909), .B2(new_n902), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT126), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n723), .A2(new_n1121), .A3(new_n810), .A4(new_n906), .ZN(new_n1122));
  AOI21_X1  g0922(.A(KEYINPUT31), .B1(new_n916), .B2(new_n917), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n720), .B1(new_n1123), .B2(new_n717), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1124), .A2(new_n722), .A3(new_n914), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1125), .A2(G330), .A3(new_n810), .A4(new_n906), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(KEYINPUT126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n736), .A2(new_n807), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n808), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n906), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n902), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n891), .A2(new_n892), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n886), .B1(new_n1133), .B2(KEYINPUT38), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1120), .A2(new_n1128), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1134), .A2(new_n1132), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n906), .B2(new_n1130), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n840), .A2(new_n908), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n906), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1132), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1138), .B1(new_n1141), .B2(new_n1119), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n919), .A2(G330), .A3(new_n920), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1136), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1118), .B1(new_n1144), .B2(new_n741), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n441), .A2(G330), .A3(new_n919), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n919), .A2(G330), .A3(new_n810), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1130), .B1(new_n907), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1128), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1125), .A2(G330), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n907), .B1(new_n1150), .B2(new_n809), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n1143), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n1139), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1149), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n864), .A2(new_n1146), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n695), .B1(new_n1155), .B2(new_n1144), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1120), .A2(new_n1128), .A3(new_n1135), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1143), .B1(new_n1120), .B2(new_n1135), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1146), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n855), .B(new_n1160), .C1(new_n861), .C2(new_n863), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1159), .A2(new_n1161), .A3(new_n1154), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1145), .B1(new_n1156), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(G378));
  INV_X1    g0964(.A(new_n312), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1165), .B(new_n669), .C1(new_n292), .C2(new_n298), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n312), .B1(new_n299), .B2(new_n888), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(KEYINPUT40), .A2(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1171), .B1(new_n1172), .B2(new_n701), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1171), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n926), .A2(G330), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n912), .A2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n903), .A2(new_n1173), .A3(new_n1175), .A4(new_n911), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1171), .A2(new_n747), .ZN(new_n1180));
  NOR3_X1   g0980(.A1(new_n753), .A2(G50), .A3(new_n747), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n766), .A2(G125), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n780), .B2(new_n828), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n760), .A2(G128), .B1(new_n784), .B2(G137), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n776), .B2(new_n1108), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1183), .B(new_n1185), .C1(G150), .C2(new_n764), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n773), .A2(G159), .ZN(new_n1190));
  AOI211_X1 g0990(.A(G33), .B(G41), .C1(new_n770), .C2(G124), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n759), .A2(new_n318), .B1(new_n769), .B2(new_n939), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n951), .B1(new_n255), .B2(new_n776), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(new_n564), .C2(new_n784), .ZN(new_n1195));
  INV_X1    g0995(.A(G41), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n813), .A2(new_n447), .B1(new_n772), .B2(new_n202), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G97), .B2(new_n779), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1195), .A2(new_n1196), .A3(new_n366), .A4(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT58), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1202));
  AOI21_X1  g1002(.A(G50), .B1(new_n258), .B2(new_n1196), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n442), .B2(G41), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1192), .A2(new_n1201), .A3(new_n1202), .A4(new_n1204), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n752), .B(new_n1181), .C1(new_n1205), .C2(new_n753), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1179), .A2(new_n742), .B1(new_n1180), .B2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n862), .B1(new_n732), .B2(new_n857), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n863), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n662), .B(new_n1146), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n1159), .B2(new_n1154), .ZN(new_n1211));
  AND4_X1   g1011(.A1(new_n911), .A2(new_n903), .A3(new_n1173), .A4(new_n1175), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n911), .A2(new_n903), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1213));
  OAI21_X1  g1013(.A(KEYINPUT57), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n694), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1149), .A2(new_n1153), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1161), .B1(new_n1144), .B2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(KEYINPUT57), .B1(new_n1217), .B2(new_n1179), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1207), .B1(new_n1215), .B2(new_n1218), .ZN(G375));
  NAND2_X1  g1019(.A1(new_n907), .A2(new_n747), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n447), .A2(new_n780), .B1(new_n813), .B2(new_n471), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G97), .B2(new_n789), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n759), .A2(new_n939), .B1(new_n757), .B2(new_n318), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n315), .B(new_n1223), .C1(G303), .C2(new_n770), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1222), .A2(new_n956), .A3(new_n1033), .A4(new_n1224), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n757), .A2(new_n952), .B1(new_n769), .B2(new_n1101), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G137), .B2(new_n760), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1108), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G50), .A2(new_n764), .B1(new_n779), .B2(new_n1228), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n766), .A2(G132), .B1(new_n789), .B2(G159), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n366), .B1(new_n773), .B2(G58), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1227), .A2(new_n1229), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n754), .B1(new_n1225), .B2(new_n1232), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n752), .B(new_n1233), .C1(new_n203), .C2(new_n835), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1154), .A2(new_n742), .B1(new_n1220), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1155), .A2(new_n998), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1154), .B1(new_n864), .B2(new_n1146), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(G381));
  NAND3_X1  g1038(.A1(new_n1061), .A2(new_n803), .A3(new_n1062), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1239), .A2(G381), .ZN(new_n1240));
  INV_X1    g1040(.A(G375), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(G384), .A2(G387), .A3(G390), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .A4(new_n1163), .ZN(G407));
  INV_X1    g1043(.A(G343), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(G213), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(G375), .A2(G378), .A3(new_n1245), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT127), .Z(new_n1247));
  NAND3_X1  g1047(.A1(new_n1247), .A2(G213), .A3(G407), .ZN(G409));
  NOR2_X1   g1048(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1211), .A2(new_n1249), .A3(new_n997), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1180), .A2(new_n1206), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n1249), .B2(new_n741), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1163), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(G375), .B2(new_n1163), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1245), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1237), .B1(KEYINPUT60), .B2(new_n1155), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1210), .A2(KEYINPUT60), .A3(new_n1216), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n694), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1235), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(G384), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n844), .B(new_n1235), .C1(new_n1256), .C2(new_n1258), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1244), .A2(G213), .A3(G2897), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1263), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1260), .A2(new_n1261), .A3(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1255), .A2(new_n1264), .A3(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1254), .A2(new_n1262), .A3(new_n1245), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT62), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT61), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT62), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1254), .A2(new_n1262), .A3(new_n1271), .A4(new_n1245), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1267), .A2(new_n1269), .A3(new_n1270), .A4(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G390), .B(new_n968), .C1(new_n999), .C2(new_n1018), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(G387), .A2(new_n1071), .A3(new_n1098), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1062), .ZN(new_n1277));
  OAI21_X1  g1077(.A(G396), .B1(new_n1277), .B2(new_n1060), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1239), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1276), .A2(new_n1279), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1274), .A2(new_n1278), .A3(new_n1239), .A4(new_n1275), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1273), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT63), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1282), .B1(new_n1284), .B2(new_n1268), .ZN(new_n1285));
  OR2_X1    g1085(.A1(new_n1268), .A2(new_n1284), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1285), .A2(new_n1286), .A3(new_n1270), .A4(new_n1267), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1283), .A2(new_n1287), .ZN(G405));
  INV_X1    g1088(.A(new_n1262), .ZN(new_n1289));
  AND2_X1   g1089(.A1(G375), .A2(new_n1163), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(G375), .A2(new_n1163), .ZN(new_n1291));
  OR3_X1    g1091(.A1(new_n1289), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1282), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1289), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1292), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1293), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(G402));
endmodule


