//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 1 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n551,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n576, new_n577, new_n578, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1144, new_n1145, new_n1146, new_n1147;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(KEYINPUT66), .A3(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n459), .A2(G2104), .ZN(new_n464));
  NAND4_X1  g039(.A1(new_n460), .A2(new_n462), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G137), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n464), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n461), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n467), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NAND4_X1  g052(.A1(new_n460), .A2(new_n462), .A3(G2105), .A4(new_n464), .ZN(new_n478));
  INV_X1    g053(.A(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n480), .B(new_n481), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n485), .B1(new_n466), .B2(G136), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n482), .A2(new_n486), .ZN(G162));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(G114), .B2(new_n463), .ZN(new_n490));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n478), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT4), .B1(new_n465), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g069(.A(KEYINPUT68), .B(KEYINPUT4), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n493), .A2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n495), .A2(new_n469), .A3(new_n464), .A4(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n492), .B1(new_n494), .B2(new_n497), .ZN(G164));
  AND2_X1   g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n502), .A2(G62), .ZN(new_n509));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  XNOR2_X1  g085(.A(new_n510), .B(KEYINPUT69), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n508), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n507), .A2(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n515), .B1(new_n516), .B2(KEYINPUT70), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G51), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT72), .B(G89), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n516), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(G63), .A2(G651), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n502), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT71), .ZN(new_n531));
  XOR2_X1   g106(.A(new_n531), .B(KEYINPUT7), .Z(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(G168));
  NAND2_X1  g108(.A1(new_n522), .A2(G52), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n501), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n501), .A2(new_n506), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n537), .A2(G651), .B1(new_n538), .B2(G90), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(G171));
  AOI22_X1  g116(.A1(new_n502), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n508), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n522), .A2(G43), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n538), .A2(G81), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  XOR2_X1   g125(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n551));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(new_n538), .A2(G91), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n502), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n556), .B2(new_n508), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT70), .B1(new_n504), .B2(new_n505), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n521), .A2(new_n560), .A3(G53), .A4(G543), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT74), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n517), .A2(KEYINPUT74), .A3(G53), .A4(new_n521), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT9), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT75), .A4(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g144(.A(KEYINPUT76), .B(KEYINPUT9), .Z(new_n570));
  NOR2_X1   g145(.A1(new_n561), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n559), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  AOI211_X1 g148(.A(KEYINPUT77), .B(new_n571), .C1(new_n567), .C2(new_n568), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n558), .B1(new_n573), .B2(new_n574), .ZN(G299));
  NOR2_X1   g150(.A1(G171), .A2(KEYINPUT78), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n534), .A2(KEYINPUT78), .A3(new_n539), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G301));
  INV_X1    g154(.A(G168), .ZN(G286));
  NAND2_X1  g155(.A1(new_n522), .A2(G49), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n581), .B(new_n582), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n502), .A2(G74), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n584), .A2(G651), .B1(G87), .B2(new_n538), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n586), .B(new_n587), .ZN(G288));
  NAND3_X1  g163(.A1(new_n502), .A2(KEYINPUT81), .A3(G61), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n501), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n589), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G651), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n502), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n506), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(new_n508), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n522), .A2(G47), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n538), .A2(G85), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(new_n538), .A2(G92), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT10), .Z(new_n605));
  NAND2_X1  g180(.A1(new_n522), .A2(G54), .ZN(new_n606));
  XNOR2_X1  g181(.A(KEYINPUT82), .B(G66), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n502), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  AND2_X1   g184(.A1(G79), .A2(G543), .ZN(new_n610));
  OAI21_X1  g185(.A(G651), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n605), .A2(new_n606), .A3(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(new_n578), .B2(G868), .ZN(G284));
  AOI21_X1  g189(.A(new_n613), .B1(new_n578), .B2(G868), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n569), .A2(new_n572), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(KEYINPUT77), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n571), .B1(new_n567), .B2(new_n568), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n559), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n557), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n616), .B1(new_n621), .B2(G868), .ZN(G297));
  OAI21_X1  g197(.A(new_n616), .B1(new_n621), .B2(G868), .ZN(G280));
  INV_X1    g198(.A(new_n612), .ZN(new_n624));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G860), .ZN(G148));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n546), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n612), .A2(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(new_n627), .ZN(G323));
  XNOR2_X1  g205(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n631));
  XNOR2_X1  g206(.A(G323), .B(new_n631), .ZN(G282));
  NAND2_X1  g207(.A1(new_n466), .A2(G135), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT84), .Z(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  INV_X1    g210(.A(G111), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n635), .A2(KEYINPUT85), .B1(new_n636), .B2(G2105), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(KEYINPUT85), .B2(new_n635), .ZN(new_n638));
  INV_X1    g213(.A(new_n478), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G123), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n634), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2096), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(G2096), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2100), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n642), .A2(new_n643), .A3(new_n647), .ZN(G156));
  XOR2_X1   g223(.A(KEYINPUT86), .B(KEYINPUT14), .Z(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2430), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n651), .B2(new_n652), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n654), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  AND3_X1   g237(.A1(new_n661), .A2(G14), .A3(new_n662), .ZN(G401));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n666), .A2(KEYINPUT17), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  AOI21_X1  g243(.A(KEYINPUT18), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n666), .B2(KEYINPUT18), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n669), .B(new_n671), .Z(new_n672));
  XOR2_X1   g247(.A(G2096), .B(G2100), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G227));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT19), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n679), .A2(new_n680), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  MUX2_X1   g261(.A(new_n686), .B(new_n685), .S(new_n678), .Z(new_n687));
  NOR2_X1   g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT87), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1991), .B(G1996), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n691), .A2(new_n692), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n691), .A2(new_n692), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n694), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n696), .A2(new_n699), .ZN(G229));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G25), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n466), .A2(G131), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT88), .ZN(new_n704));
  OAI21_X1  g279(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n705));
  INV_X1    g280(.A(G107), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(G2105), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n639), .B2(G119), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n702), .B1(new_n710), .B2(new_n701), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT35), .B(G1991), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(G16), .A2(G24), .ZN(new_n714));
  INV_X1    g289(.A(G290), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(G16), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT89), .B(G1986), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G22), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G166), .B2(new_n719), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G1971), .ZN(new_n722));
  MUX2_X1   g297(.A(G6), .B(G305), .S(G16), .Z(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT32), .B(G1981), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  NOR3_X1   g301(.A1(new_n722), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n719), .A2(G23), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n583), .A2(new_n585), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n719), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT33), .B(G1976), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n730), .A2(new_n732), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n727), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n713), .B(new_n718), .C1(new_n735), .C2(KEYINPUT34), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(KEYINPUT34), .B2(new_n735), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT36), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n719), .A2(G20), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT23), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n621), .B2(new_n719), .ZN(new_n741));
  INV_X1    g316(.A(G1956), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n719), .A2(G5), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G171), .B2(new_n719), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT97), .Z(new_n746));
  INV_X1    g321(.A(G1961), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G34), .ZN(new_n749));
  AOI21_X1  g324(.A(G29), .B1(new_n749), .B2(KEYINPUT24), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(KEYINPUT24), .B2(new_n749), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n476), .B2(new_n701), .ZN(new_n752));
  INV_X1    g327(.A(G2084), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT27), .B(G1996), .ZN(new_n755));
  OAI21_X1  g330(.A(KEYINPUT93), .B1(G29), .B2(G32), .ZN(new_n756));
  INV_X1    g331(.A(G141), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n465), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n639), .A2(G129), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT92), .ZN(new_n761));
  NAND3_X1  g336(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT26), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g339(.A1(KEYINPUT26), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n764), .A2(new_n765), .B1(new_n474), .B2(G105), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n759), .A2(new_n760), .A3(new_n761), .A4(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G129), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n766), .B1(new_n478), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(KEYINPUT92), .B1(new_n769), .B2(new_n758), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(G29), .ZN(new_n772));
  MUX2_X1   g347(.A(KEYINPUT93), .B(new_n756), .S(new_n772), .Z(new_n773));
  OAI211_X1 g348(.A(new_n748), .B(new_n754), .C1(new_n755), .C2(new_n773), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT98), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n547), .A2(G16), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G16), .B2(G19), .ZN(new_n777));
  INV_X1    g352(.A(G1341), .ZN(new_n778));
  NAND2_X1  g353(.A1(G115), .A2(G2104), .ZN(new_n779));
  INV_X1    g354(.A(G127), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n470), .B2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT25), .ZN(new_n782));
  NAND2_X1  g357(.A1(G103), .A2(G2104), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(G2105), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n463), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n781), .A2(G2105), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n466), .A2(G139), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  MUX2_X1   g363(.A(G33), .B(new_n788), .S(G29), .Z(new_n789));
  AOI22_X1  g364(.A1(new_n777), .A2(new_n778), .B1(G2072), .B2(new_n789), .ZN(new_n790));
  OAI221_X1 g365(.A(new_n790), .B1(new_n778), .B2(new_n777), .C1(new_n753), .C2(new_n752), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT30), .B(G28), .ZN(new_n792));
  OR2_X1    g367(.A1(KEYINPUT31), .A2(G11), .ZN(new_n793));
  NAND2_X1  g368(.A1(KEYINPUT31), .A2(G11), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n792), .A2(new_n701), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(G168), .A2(new_n719), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n719), .B2(G21), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT94), .B(G1966), .ZN(new_n798));
  OAI221_X1 g373(.A(new_n795), .B1(G2072), .B2(new_n789), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n791), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n797), .A2(new_n798), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT96), .Z(new_n802));
  NOR2_X1   g377(.A1(G4), .A2(G16), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT90), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n612), .B2(new_n719), .ZN(new_n805));
  INV_X1    g380(.A(G1348), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n641), .A2(new_n701), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT95), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n701), .A2(G26), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT28), .ZN(new_n812));
  INV_X1    g387(.A(G128), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n463), .A2(G116), .ZN(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n815));
  OAI22_X1  g390(.A1(new_n478), .A2(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n466), .A2(KEYINPUT91), .A3(G140), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT91), .ZN(new_n818));
  INV_X1    g393(.A(G140), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n465), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n816), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n812), .B1(new_n821), .B2(new_n701), .ZN(new_n822));
  INV_X1    g397(.A(G2067), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n800), .A2(new_n802), .A3(new_n810), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n701), .A2(G35), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G162), .B2(new_n701), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT29), .Z(new_n828));
  INV_X1    g403(.A(G2090), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n701), .A2(G27), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(G164), .B2(new_n701), .ZN(new_n832));
  INV_X1    g407(.A(G2078), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n830), .B(new_n834), .C1(new_n747), .C2(new_n746), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n773), .A2(new_n755), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n828), .B2(new_n829), .ZN(new_n837));
  NOR4_X1   g412(.A1(new_n775), .A2(new_n825), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n738), .A2(new_n743), .A3(new_n838), .ZN(G150));
  INV_X1    g414(.A(G150), .ZN(G311));
  NAND2_X1  g415(.A1(new_n624), .A2(G559), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT38), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n522), .A2(G55), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n538), .A2(G93), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n843), .B(new_n844), .C1(new_n508), .C2(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n846), .A2(new_n546), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n546), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n842), .B(new_n850), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n852), .A2(new_n853), .A3(G860), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n846), .A2(G860), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT37), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n854), .A2(new_n856), .ZN(G145));
  XNOR2_X1  g432(.A(new_n641), .B(new_n476), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n767), .A2(new_n770), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n817), .A2(new_n820), .ZN(new_n861));
  INV_X1    g436(.A(new_n816), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(G164), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n494), .A2(new_n497), .ZN(new_n865));
  INV_X1    g440(.A(new_n492), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n821), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n860), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n863), .A2(G164), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n821), .A2(new_n867), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n771), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(KEYINPUT100), .B1(new_n786), .B2(new_n787), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n873), .A2(KEYINPUT99), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n869), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n788), .A2(KEYINPUT99), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(KEYINPUT99), .B2(new_n873), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n877), .B1(new_n869), .B2(new_n872), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n710), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n877), .ZN(new_n880));
  INV_X1    g455(.A(new_n872), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n771), .B1(new_n870), .B2(new_n871), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n869), .A2(new_n872), .A3(new_n874), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n883), .A2(new_n709), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n466), .A2(G142), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n639), .A2(G130), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n463), .A2(G118), .ZN(new_n888));
  OAI21_X1  g463(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n886), .B(new_n887), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n890), .B(new_n645), .Z(new_n891));
  NAND3_X1  g466(.A1(new_n879), .A2(new_n885), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT102), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n891), .B1(new_n879), .B2(new_n885), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n859), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n879), .A2(new_n885), .ZN(new_n897));
  INV_X1    g472(.A(new_n891), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n899), .A2(new_n893), .A3(new_n892), .A4(new_n858), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(G162), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n901), .B(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(KEYINPUT101), .B(G37), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g481(.A1(new_n846), .A2(new_n627), .ZN(new_n907));
  XNOR2_X1  g482(.A(G303), .B(G305), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n729), .A2(new_n715), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n586), .A2(G290), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n908), .B1(new_n911), .B2(KEYINPUT104), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(KEYINPUT104), .B2(new_n911), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n909), .A2(new_n914), .A3(new_n910), .A4(new_n908), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n916), .B(new_n917), .Z(new_n918));
  NAND2_X1  g493(.A1(G299), .A2(new_n612), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n558), .B(new_n624), .C1(new_n573), .C2(new_n574), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(KEYINPUT41), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT41), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n919), .A2(new_n924), .A3(new_n920), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  XOR2_X1   g501(.A(new_n849), .B(KEYINPUT103), .Z(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(new_n629), .ZN(new_n928));
  MUX2_X1   g503(.A(new_n922), .B(new_n926), .S(new_n928), .Z(new_n929));
  XNOR2_X1  g504(.A(new_n918), .B(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n907), .B1(new_n930), .B2(new_n627), .ZN(G295));
  OAI21_X1  g506(.A(new_n907), .B1(new_n930), .B2(new_n627), .ZN(G331));
  NOR2_X1   g507(.A1(G168), .A2(G171), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n933), .B1(new_n578), .B2(G168), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(new_n850), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n926), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n934), .B(new_n849), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n922), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT106), .B1(new_n913), .B2(new_n915), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n938), .B(new_n936), .C1(new_n916), .C2(KEYINPUT106), .ZN(new_n942));
  INV_X1    g517(.A(G37), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  OR2_X1    g519(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n945));
  INV_X1    g520(.A(new_n916), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n925), .A2(KEYINPUT107), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n919), .A2(new_n948), .A3(new_n924), .A4(new_n920), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(new_n923), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n951), .A3(new_n935), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n938), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n951), .B1(new_n950), .B2(new_n935), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n946), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n904), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n936), .A2(new_n938), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n956), .B1(new_n957), .B2(new_n916), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n945), .B(KEYINPUT44), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n955), .A2(new_n960), .A3(new_n958), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI211_X1 g542(.A(KEYINPUT109), .B(KEYINPUT44), .C1(new_n963), .C2(new_n964), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n961), .B1(new_n967), .B2(new_n968), .ZN(G397));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n867), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(G160), .A2(G40), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G1996), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n977), .A2(new_n860), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n978), .B(KEYINPUT111), .Z(new_n979));
  INV_X1    g554(.A(new_n975), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n821), .B(G2067), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n975), .A2(G1996), .A3(new_n860), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT112), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n979), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n710), .A2(new_n712), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n710), .A2(new_n712), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n975), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  OR2_X1    g564(.A1(G290), .A2(G1986), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(G290), .A2(G1986), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n992), .B(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n989), .B1(new_n975), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G8), .ZN(new_n996));
  AND2_X1   g571(.A1(G160), .A2(G40), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n973), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT114), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT114), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n973), .A2(new_n997), .A3(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(G164), .A2(G1384), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT45), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n971), .A2(KEYINPUT50), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1007), .A3(new_n997), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  AOI22_X1  g584(.A1(new_n1004), .A2(new_n798), .B1(new_n753), .B2(new_n1009), .ZN(new_n1010));
  AOI211_X1 g585(.A(KEYINPUT51), .B(new_n996), .C1(new_n1010), .C2(G168), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n996), .B1(new_n1010), .B2(G168), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(G168), .B2(new_n1010), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1011), .B1(new_n1013), .B2(KEYINPUT51), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT120), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n619), .B2(new_n557), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT116), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n621), .A2(KEYINPUT57), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n973), .A2(new_n1003), .A3(new_n997), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT56), .B(G2072), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1021), .A2(new_n1022), .B1(new_n1008), .B2(new_n742), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1023), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1018), .A2(new_n1019), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT61), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1015), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n974), .A2(new_n971), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1008), .A2(new_n806), .B1(new_n823), .B2(new_n1030), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1031), .A2(new_n612), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1031), .A2(new_n612), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT60), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT60), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1031), .A2(new_n1035), .A3(new_n624), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1021), .A2(new_n976), .ZN(new_n1039));
  XOR2_X1   g614(.A(KEYINPUT58), .B(G1341), .Z(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n974), .B2(new_n971), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1038), .B1(new_n1042), .B2(new_n547), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1042), .A2(new_n1038), .A3(new_n547), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(KEYINPUT59), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT59), .ZN(new_n1047));
  AOI211_X1 g622(.A(KEYINPUT118), .B(new_n546), .C1(new_n1039), .C2(new_n1041), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1047), .B1(new_n1043), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1037), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(KEYINPUT119), .B(KEYINPUT61), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1027), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1024), .A2(KEYINPUT120), .A3(KEYINPUT61), .A4(new_n1026), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1029), .A2(new_n1050), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1025), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1033), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1026), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1057), .B(KEYINPUT117), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n973), .A2(new_n1003), .A3(new_n997), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(new_n1061), .B2(G2078), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1062), .B(KEYINPUT121), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1060), .A2(G2078), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .A4(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1008), .A2(new_n747), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1063), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT54), .B1(new_n1067), .B2(new_n578), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT122), .B1(new_n1008), .B2(new_n747), .ZN(new_n1071));
  XOR2_X1   g646(.A(KEYINPUT123), .B(G2078), .Z(new_n1072));
  NOR3_X1   g647(.A1(new_n1061), .A2(new_n1060), .A3(new_n1072), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n540), .B1(new_n1063), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1068), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1067), .A2(new_n578), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1063), .A2(new_n1074), .A3(G301), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT54), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1030), .A2(new_n996), .ZN(new_n1080));
  INV_X1    g655(.A(G1976), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(new_n586), .ZN(new_n1082));
  AOI211_X1 g657(.A(KEYINPUT52), .B(new_n1082), .C1(G288), .C2(new_n1081), .ZN(new_n1083));
  XOR2_X1   g658(.A(G305), .B(G1981), .Z(new_n1084));
  OR2_X1    g659(.A1(new_n1084), .A2(KEYINPUT49), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(KEYINPUT49), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(new_n1086), .A3(new_n1080), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1082), .A2(KEYINPUT52), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1083), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G303), .A2(G8), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1091), .B(KEYINPUT55), .ZN(new_n1092));
  XOR2_X1   g667(.A(new_n1092), .B(KEYINPUT113), .Z(new_n1093));
  OAI22_X1  g668(.A1(new_n1021), .A2(G1971), .B1(new_n1008), .B2(G2090), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G8), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1092), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1090), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1076), .A2(new_n1079), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1059), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1098), .A2(new_n1077), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1101), .B1(new_n1014), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1014), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1010), .A2(new_n996), .A3(G286), .ZN(new_n1105));
  XOR2_X1   g680(.A(new_n1105), .B(KEYINPUT115), .Z(new_n1106));
  INV_X1    g681(.A(new_n1098), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT63), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1101), .A2(KEYINPUT62), .A3(new_n1014), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT63), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1106), .A2(new_n1107), .A3(new_n1111), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1096), .A2(new_n1083), .A3(new_n1089), .ZN(new_n1113));
  NOR2_X1   g688(.A1(G288), .A2(G1976), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1087), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(G1981), .B2(G305), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1113), .B1(new_n1080), .B2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1109), .A2(new_n1110), .A3(new_n1112), .A4(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n995), .B1(new_n1104), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(KEYINPUT124), .A2(KEYINPUT46), .ZN(new_n1120));
  XOR2_X1   g695(.A(new_n977), .B(new_n1120), .Z(new_n1121));
  NAND2_X1  g696(.A1(new_n981), .A2(new_n771), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1122), .A2(new_n975), .B1(KEYINPUT124), .B2(KEYINPUT46), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(KEYINPUT47), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n980), .A2(new_n990), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1126), .B(KEYINPUT126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT125), .B(KEYINPUT48), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1127), .B(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1125), .B1(new_n989), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n985), .A2(new_n986), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n821), .A2(new_n823), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n980), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1119), .A2(new_n1134), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g710(.A1(new_n674), .A2(G319), .ZN(new_n1137));
  NOR2_X1   g711(.A1(G401), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g712(.A(new_n1138), .B1(new_n696), .B2(new_n699), .ZN(new_n1139));
  AOI21_X1  g713(.A(new_n1139), .B1(new_n903), .B2(new_n904), .ZN(new_n1140));
  AND3_X1   g714(.A1(new_n965), .A2(new_n1140), .A3(KEYINPUT127), .ZN(new_n1141));
  AOI21_X1  g715(.A(KEYINPUT127), .B1(new_n965), .B2(new_n1140), .ZN(new_n1142));
  NOR2_X1   g716(.A1(new_n1141), .A2(new_n1142), .ZN(G308));
  NAND2_X1  g717(.A1(new_n965), .A2(new_n1140), .ZN(new_n1144));
  INV_X1    g718(.A(KEYINPUT127), .ZN(new_n1145));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g720(.A1(new_n965), .A2(new_n1140), .A3(KEYINPUT127), .ZN(new_n1147));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n1147), .ZN(G225));
endmodule


