//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n865, new_n866, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT100), .ZN(new_n203));
  XOR2_X1   g002(.A(G134gat), .B(G162gat), .Z(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(KEYINPUT17), .ZN(new_n206));
  NOR2_X1   g005(.A1(G29gat), .A2(G36gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT14), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT87), .B(G36gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G29gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT15), .ZN(new_n213));
  OR2_X1    g012(.A1(G43gat), .A2(G50gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(G43gat), .A2(G50gat), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n216), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n214), .A2(new_n213), .A3(new_n215), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n218), .A2(new_n209), .A3(new_n211), .A4(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n206), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT88), .ZN(new_n222));
  AND4_X1   g021(.A1(new_n218), .A2(new_n209), .A3(new_n211), .A4(new_n219), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n218), .B1(new_n209), .B2(new_n211), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n217), .A2(KEYINPUT88), .A3(new_n220), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n221), .B1(new_n227), .B2(new_n206), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT98), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230));
  NAND2_X1  g029(.A1(G99gat), .A2(G106gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT97), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(new_n232), .B2(new_n231), .ZN(new_n234));
  OAI211_X1 g033(.A(KEYINPUT96), .B(KEYINPUT7), .C1(G85gat), .C2(G92gat), .ZN(new_n235));
  INV_X1    g034(.A(G85gat), .ZN(new_n236));
  INV_X1    g035(.A(G92gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND4_X1  g037(.A1(KEYINPUT96), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n234), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(G99gat), .B(G106gat), .Z(new_n241));
  AOI21_X1  g040(.A(new_n229), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n241), .ZN(new_n243));
  INV_X1    g042(.A(new_n241), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n244), .A2(new_n234), .A3(new_n238), .A4(new_n239), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n242), .B1(new_n246), .B2(new_n229), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n228), .A2(new_n247), .ZN(new_n248));
  NOR3_X1   g047(.A1(new_n223), .A2(new_n224), .A3(new_n222), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT88), .B1(new_n217), .B2(new_n220), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n247), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT41), .ZN(new_n253));
  INV_X1    g052(.A(G232gat), .ZN(new_n254));
  INV_X1    g053(.A(G233gat), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n252), .A2(KEYINPUT99), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT99), .B1(new_n252), .B2(new_n257), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n248), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n261), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n248), .B(new_n263), .C1(new_n258), .C2(new_n259), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n205), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n262), .A2(new_n264), .A3(new_n205), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(G71gat), .B(G78gat), .Z(new_n270));
  INV_X1    g069(.A(KEYINPUT92), .ZN(new_n271));
  NAND2_X1  g070(.A1(G71gat), .A2(G78gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT9), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n270), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G64gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G57gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT91), .B(G57gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n277), .B1(new_n278), .B2(new_n276), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n275), .B(new_n279), .C1(new_n271), .C2(new_n274), .ZN(new_n280));
  XNOR2_X1  g079(.A(G57gat), .B(G64gat), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n270), .B1(new_n273), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(KEYINPUT21), .ZN(new_n285));
  XNOR2_X1  g084(.A(G127gat), .B(G155gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G183gat), .B(G211gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G15gat), .B(G22gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT16), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n291), .B1(new_n292), .B2(G1gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(G1gat), .B2(new_n291), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n294), .A2(G8gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(G8gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT94), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT94), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n280), .A2(new_n300), .A3(new_n282), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n298), .B1(new_n302), .B2(KEYINPUT21), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT95), .ZN(new_n304));
  OR2_X1    g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n304), .ZN(new_n306));
  NAND2_X1  g105(.A1(G231gat), .A2(G233gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT93), .ZN(new_n308));
  XOR2_X1   g107(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n309));
  XOR2_X1   g108(.A(new_n308), .B(new_n309), .Z(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n305), .A2(new_n306), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n311), .B1(new_n305), .B2(new_n306), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n290), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n314), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(new_n289), .A3(new_n312), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n269), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G229gat), .A2(G233gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n251), .A2(new_n298), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n320), .B(new_n321), .C1(new_n228), .C2(new_n298), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT89), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n206), .B1(new_n249), .B2(new_n250), .ZN(new_n325));
  INV_X1    g124(.A(new_n221), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n297), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n328), .A2(KEYINPUT89), .A3(new_n320), .A4(new_n321), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n324), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n298), .B1(new_n325), .B2(new_n326), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n227), .A2(new_n297), .ZN(new_n333));
  INV_X1    g132(.A(new_n320), .ZN(new_n334));
  NOR3_X1   g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n227), .A2(new_n297), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n336), .ZN(new_n337));
  XOR2_X1   g136(.A(new_n320), .B(KEYINPUT13), .Z(new_n338));
  AOI22_X1  g137(.A1(new_n335), .A2(KEYINPUT18), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G113gat), .B(G141gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(G197gat), .ZN(new_n341));
  XOR2_X1   g140(.A(KEYINPUT11), .B(G169gat), .Z(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n331), .A2(new_n339), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n345), .B1(new_n331), .B2(new_n339), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT101), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT10), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n280), .A2(new_n243), .A3(new_n245), .A4(new_n282), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n350), .B(new_n351), .C1(new_n247), .C2(new_n284), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n299), .A2(new_n247), .A3(KEYINPUT10), .A4(new_n301), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G230gat), .A2(G233gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n351), .B1(new_n247), .B2(new_n284), .ZN(new_n357));
  INV_X1    g156(.A(new_n355), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G120gat), .B(G148gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(G176gat), .B(G204gat), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  NAND3_X1  g161(.A1(new_n356), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n362), .B1(new_n356), .B2(new_n359), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n349), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n365), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(KEYINPUT101), .A3(new_n363), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n319), .A2(new_n348), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT69), .ZN(new_n373));
  INV_X1    g172(.A(G127gat), .ZN(new_n374));
  OR2_X1    g173(.A1(new_n374), .A2(G134gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(G134gat), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(G120gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(G113gat), .ZN(new_n379));
  INV_X1    g178(.A(G113gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G120gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT66), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT1), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G113gat), .B(G120gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT66), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n377), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT1), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n375), .A2(new_n376), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT67), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(new_n378), .A3(G113gat), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n391), .A2(new_n381), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n379), .A2(KEYINPUT67), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n389), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n387), .A2(new_n394), .A3(KEYINPUT68), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT68), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n375), .A2(new_n376), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n388), .B1(new_n385), .B2(KEYINPUT66), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n379), .A2(new_n381), .A3(KEYINPUT66), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n393), .A2(new_n391), .A3(new_n381), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n377), .A2(new_n401), .A3(new_n388), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n396), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n373), .B1(new_n395), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT64), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT25), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(G169gat), .ZN(new_n408));
  INV_X1    g207(.A(G176gat), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT23), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT23), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(G169gat), .B2(G176gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(G169gat), .A2(G176gat), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n410), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(G183gat), .A2(G190gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AND2_X1   g217(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G190gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n414), .A2(new_n415), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n415), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n417), .A2(new_n416), .B1(new_n419), .B2(G190gat), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n410), .A2(new_n412), .A3(new_n413), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n407), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n413), .ZN(new_n429));
  NOR3_X1   g228(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n417), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  XOR2_X1   g230(.A(KEYINPUT27), .B(G183gat), .Z(new_n432));
  INV_X1    g231(.A(G190gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT28), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n437));
  AOI21_X1  g236(.A(G190gat), .B1(new_n437), .B2(KEYINPUT27), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT27), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n439), .A2(KEYINPUT65), .A3(G183gat), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT28), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n431), .B1(new_n436), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n427), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT68), .B1(new_n387), .B2(new_n394), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n400), .A2(new_n396), .A3(new_n402), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(KEYINPUT69), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n404), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(G227gat), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n450), .A2(new_n255), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n444), .B(new_n373), .C1(new_n403), .C2(new_n395), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT32), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT33), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g255(.A(G15gat), .B(G43gat), .Z(new_n457));
  XNOR2_X1  g256(.A(G71gat), .B(G99gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n454), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n459), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n453), .B(KEYINPUT32), .C1(new_n455), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n449), .A2(new_n452), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT34), .B1(new_n465), .B2(new_n451), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT34), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n464), .B(new_n467), .C1(new_n450), .C2(new_n255), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n463), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n460), .A2(new_n466), .A3(new_n468), .A4(new_n462), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT70), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(KEYINPUT70), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G197gat), .B(G204gat), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT22), .ZN(new_n477));
  INV_X1    g276(.A(G211gat), .ZN(new_n478));
  INV_X1    g277(.A(G218gat), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  XOR2_X1   g280(.A(G211gat), .B(G218gat), .Z(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  AND2_X1   g282(.A1(G155gat), .A2(G162gat), .ZN(new_n484));
  NOR2_X1   g283(.A1(G155gat), .A2(G162gat), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G141gat), .B(G148gat), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT2), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(G155gat), .B2(G162gat), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n486), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(G141gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(G148gat), .ZN(new_n492));
  INV_X1    g291(.A(G148gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(G141gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G155gat), .B(G162gat), .ZN(new_n496));
  INV_X1    g295(.A(G155gat), .ZN(new_n497));
  INV_X1    g296(.A(G162gat), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT2), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n495), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT3), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n490), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  XOR2_X1   g301(.A(KEYINPUT71), .B(KEYINPUT29), .Z(new_n503));
  AOI21_X1  g302(.A(new_n483), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n504), .B1(G228gat), .B2(G233gat), .ZN(new_n505));
  INV_X1    g304(.A(new_n483), .ZN(new_n506));
  INV_X1    g305(.A(new_n503), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n501), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n500), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n490), .A2(new_n500), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT29), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n483), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n512), .B1(new_n514), .B2(new_n501), .ZN(new_n515));
  OAI211_X1 g314(.A(G228gat), .B(G233gat), .C1(new_n515), .C2(new_n504), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(KEYINPUT31), .B(G50gat), .Z(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G78gat), .B(G106gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(G22gat), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n519), .B(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n524), .A2(KEYINPUT35), .ZN(new_n525));
  INV_X1    g324(.A(G226gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n526), .A2(new_n255), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(new_n427), .B2(new_n443), .ZN(new_n528));
  INV_X1    g327(.A(new_n407), .ZN(new_n529));
  NOR3_X1   g328(.A1(new_n424), .A2(new_n425), .A3(new_n423), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n415), .B1(new_n414), .B2(new_n421), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI221_X1 g331(.A(new_n417), .B1(new_n430), .B2(new_n429), .C1(new_n435), .C2(new_n441), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT29), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n483), .B(new_n528), .C1(new_n534), .C2(new_n527), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT72), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n527), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(new_n444), .B2(KEYINPUT29), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n539), .A2(KEYINPUT72), .A3(new_n483), .A4(new_n528), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n507), .B1(new_n532), .B2(new_n533), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n528), .B1(new_n541), .B2(new_n527), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n506), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n537), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G8gat), .B(G36gat), .Z(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT73), .ZN(new_n546));
  XNOR2_X1  g345(.A(G64gat), .B(G92gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n550), .A2(KEYINPUT74), .A3(KEYINPUT30), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n535), .A2(new_n536), .B1(new_n542), .B2(new_n506), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n552), .A2(KEYINPUT30), .A3(new_n540), .A4(new_n548), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n544), .A2(new_n549), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT74), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT30), .ZN(new_n557));
  INV_X1    g356(.A(new_n550), .ZN(new_n558));
  AOI22_X1  g357(.A1(new_n551), .A2(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G225gat), .A2(G233gat), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n490), .A2(new_n500), .A3(new_n501), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n501), .B1(new_n490), .B2(new_n500), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n400), .A2(new_n402), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n512), .A2(new_n400), .A3(new_n402), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT4), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n446), .A2(new_n512), .A3(new_n447), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n567), .B(new_n570), .C1(new_n571), .C2(new_n569), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT76), .B(KEYINPUT5), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n509), .B1(new_n387), .B2(new_n394), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n568), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n573), .B1(new_n575), .B2(new_n562), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n568), .A2(new_n569), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n577), .B1(new_n571), .B2(new_n569), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n495), .A2(new_n496), .A3(new_n499), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n496), .B1(new_n499), .B2(new_n495), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT3), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n581), .B(new_n502), .C1(new_n387), .C2(new_n394), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n582), .A2(new_n561), .A3(new_n573), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n572), .A2(new_n576), .B1(new_n578), .B2(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(G1gat), .B(G29gat), .Z(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G57gat), .B(G85gat), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n587), .B(new_n588), .Z(new_n589));
  AOI21_X1  g388(.A(KEYINPUT6), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n589), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n591), .B1(new_n584), .B2(KEYINPUT80), .ZN(new_n592));
  AND4_X1   g391(.A1(KEYINPUT4), .A2(new_n446), .A3(new_n512), .A4(new_n447), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n570), .A2(new_n561), .A3(new_n582), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n576), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n571), .A2(new_n569), .ZN(new_n596));
  INV_X1    g395(.A(new_n577), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n583), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT80), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n590), .B1(new_n592), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT79), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT6), .ZN(new_n604));
  NOR4_X1   g403(.A1(new_n584), .A2(new_n603), .A3(new_n604), .A4(new_n589), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n589), .B1(new_n595), .B2(new_n598), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT79), .B1(new_n607), .B2(KEYINPUT6), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n602), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n560), .A2(new_n610), .A3(KEYINPUT84), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT84), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n605), .A2(new_n608), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n602), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n612), .B1(new_n559), .B2(new_n614), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n475), .B(new_n525), .C1(new_n611), .C2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n470), .ZN(new_n617));
  INV_X1    g416(.A(new_n471), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n523), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n551), .A2(new_n556), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT75), .ZN(new_n622));
  OAI21_X1  g421(.A(KEYINPUT78), .B1(new_n584), .B2(new_n589), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT78), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n590), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n613), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT75), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n551), .A2(new_n556), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n558), .A2(new_n557), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n622), .A2(new_n627), .A3(new_n629), .A4(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT35), .B1(new_n620), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n524), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT36), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n635), .B1(new_n470), .B2(new_n471), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n636), .B1(new_n475), .B2(new_n635), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n561), .B1(new_n578), .B2(new_n582), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT39), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(KEYINPUT39), .B1(new_n575), .B2(new_n562), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n589), .B1(new_n639), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n638), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n639), .A2(new_n643), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n646), .A2(KEYINPUT40), .A3(new_n589), .A4(new_n641), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n645), .B(new_n647), .C1(new_n601), .C2(new_n592), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n523), .B1(new_n559), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT38), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT37), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n552), .A2(new_n651), .A3(new_n540), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n652), .A2(new_n549), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n544), .A2(KEYINPUT37), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n506), .B(new_n528), .C1(new_n534), .C2(new_n527), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(KEYINPUT37), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n538), .B1(new_n444), .B2(new_n507), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n506), .B1(new_n658), .B2(new_n528), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT38), .B1(new_n660), .B2(KEYINPUT81), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT81), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n657), .B2(new_n659), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n661), .A2(new_n549), .A3(new_n652), .A4(new_n663), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n664), .A2(new_n613), .A3(new_n558), .A4(new_n602), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n655), .B1(new_n665), .B2(KEYINPUT82), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT82), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n610), .A2(new_n667), .A3(new_n558), .A4(new_n664), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n649), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n634), .B(new_n637), .C1(new_n669), .C2(KEYINPUT83), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT83), .ZN(new_n671));
  AOI211_X1 g470(.A(new_n671), .B(new_n649), .C1(new_n668), .C2(new_n666), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n633), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT85), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n633), .B(KEYINPUT85), .C1(new_n670), .C2(new_n672), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n372), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n627), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g479(.A1(new_n677), .A2(new_n560), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(KEYINPUT103), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n677), .A2(new_n683), .A3(new_n560), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n682), .A2(G8gat), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT16), .B(G8gat), .Z(new_n686));
  NAND4_X1  g485(.A1(new_n677), .A2(KEYINPUT42), .A3(new_n560), .A4(new_n686), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n682), .A2(new_n684), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n686), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n689), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n686), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n695), .B1(new_n682), .B2(new_n684), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n696), .A2(KEYINPUT104), .A3(new_n692), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n688), .B1(new_n694), .B2(new_n697), .ZN(G1325gat));
  INV_X1    g497(.A(new_n677), .ZN(new_n699));
  OAI21_X1  g498(.A(G15gat), .B1(new_n699), .B2(new_n637), .ZN(new_n700));
  INV_X1    g499(.A(new_n475), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n701), .A2(G15gat), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n700), .B1(new_n699), .B2(new_n702), .ZN(G1326gat));
  NAND2_X1  g502(.A1(new_n677), .A2(new_n524), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT43), .B(G22gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  NAND2_X1  g505(.A1(new_n675), .A2(new_n676), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n318), .A2(new_n370), .A3(new_n348), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(new_n268), .A3(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(G29gat), .A3(new_n627), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT45), .Z(new_n711));
  OR2_X1    g510(.A1(new_n669), .A2(KEYINPUT83), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n637), .A2(new_n634), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n669), .A2(KEYINPUT83), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n269), .B1(new_n715), .B2(new_n633), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n269), .B1(new_n675), .B2(new_n676), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(new_n717), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n708), .ZN(new_n721));
  OAI21_X1  g520(.A(G29gat), .B1(new_n721), .B2(new_n627), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n711), .A2(new_n722), .ZN(G1328gat));
  NOR3_X1   g522(.A1(new_n709), .A2(new_n559), .A3(new_n210), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n210), .B1(new_n721), .B2(new_n559), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1329gat));
  INV_X1    g527(.A(new_n637), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(G43gat), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n709), .A2(new_n701), .ZN(new_n731));
  OAI22_X1  g530(.A1(new_n721), .A2(new_n730), .B1(new_n731), .B2(G43gat), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g532(.A(new_n717), .B1(new_n707), .B2(new_n268), .ZN(new_n734));
  INV_X1    g533(.A(new_n718), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n524), .B(new_n708), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT107), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n720), .A2(new_n738), .A3(new_n524), .A4(new_n708), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n737), .A2(G50gat), .A3(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT48), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n709), .A2(KEYINPUT106), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n719), .A2(new_n743), .A3(new_n708), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n523), .A2(G50gat), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n741), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n740), .A2(new_n747), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n736), .A2(G50gat), .ZN(new_n749));
  AOI211_X1 g548(.A(G50gat), .B(new_n523), .C1(new_n742), .C2(new_n744), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n741), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n751), .ZN(G1331gat));
  AOI21_X1  g551(.A(new_n268), .B1(new_n317), .B2(new_n315), .ZN(new_n753));
  AND4_X1   g552(.A1(new_n673), .A2(new_n348), .A3(new_n370), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n678), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(new_n278), .ZN(G1332gat));
  INV_X1    g555(.A(KEYINPUT49), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n560), .B1(new_n757), .B2(new_n276), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT108), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n754), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n276), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1333gat));
  NAND3_X1  g561(.A1(new_n754), .A2(G71gat), .A3(new_n729), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n475), .B(KEYINPUT109), .Z(new_n764));
  AND2_X1   g563(.A1(new_n754), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n765), .B2(G71gat), .ZN(new_n766));
  XOR2_X1   g565(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(G1334gat));
  NAND2_X1  g567(.A1(new_n754), .A2(new_n524), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT112), .ZN(new_n770));
  XNOR2_X1  g569(.A(KEYINPUT111), .B(G78gat), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1335gat));
  INV_X1    g571(.A(new_n348), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n773), .A2(new_n318), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n720), .A2(new_n370), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(G85gat), .B1(new_n775), .B2(new_n627), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n716), .A2(new_n777), .A3(new_n774), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n673), .A2(new_n268), .ZN(new_n779));
  INV_X1    g578(.A(new_n774), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT51), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n778), .A2(new_n781), .A3(new_n370), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n783), .A2(new_n236), .A3(new_n678), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n776), .A2(new_n784), .ZN(G1336gat));
  OAI21_X1  g584(.A(G92gat), .B1(new_n775), .B2(new_n559), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n560), .A2(new_n237), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n786), .B(new_n787), .C1(new_n782), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n370), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT85), .B1(new_n715), .B2(new_n633), .ZN(new_n791));
  INV_X1    g590(.A(new_n676), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n268), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT44), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n790), .B1(new_n794), .B2(new_n718), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n237), .B1(new_n795), .B2(new_n560), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n782), .A2(new_n788), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT52), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n789), .A2(new_n798), .ZN(G1337gat));
  OAI21_X1  g598(.A(G99gat), .B1(new_n775), .B2(new_n637), .ZN(new_n800));
  OR3_X1    g599(.A1(new_n782), .A2(G99gat), .A3(new_n701), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(G1338gat));
  INV_X1    g601(.A(G106gat), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(new_n782), .B2(new_n523), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n524), .A2(G106gat), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n775), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n806), .B(new_n807), .ZN(G1339gat));
  NAND3_X1  g607(.A1(new_n753), .A2(new_n348), .A3(new_n369), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n358), .B1(new_n352), .B2(new_n353), .ZN(new_n811));
  XNOR2_X1  g610(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n362), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n356), .A2(KEYINPUT54), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n354), .A2(new_n355), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n267), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n818), .B1(new_n819), .B2(new_n265), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n331), .A2(new_n339), .A3(new_n345), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n320), .B1(new_n328), .B2(new_n321), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n337), .A2(new_n338), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n343), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g624(.A(KEYINPUT55), .B(new_n813), .C1(new_n814), .C2(new_n815), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n363), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n820), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n366), .A2(new_n368), .A3(new_n821), .A4(new_n824), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n818), .B1(new_n346), .B2(new_n347), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n830), .B(KEYINPUT114), .C1(new_n831), .C2(new_n827), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n269), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n826), .A2(new_n363), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n834), .B(new_n818), .C1(new_n347), .C2(new_n346), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT114), .B1(new_n835), .B2(new_n830), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n829), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n318), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n810), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n839), .A2(new_n627), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n620), .A2(new_n560), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(new_n380), .A3(new_n773), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(new_n839), .B2(new_n524), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n830), .B1(new_n831), .B2(new_n827), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n269), .A3(new_n832), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n318), .B1(new_n851), .B2(new_n829), .ZN(new_n852));
  OAI211_X1 g651(.A(KEYINPUT115), .B(new_n523), .C1(new_n852), .C2(new_n810), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n847), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n560), .A2(new_n627), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(new_n475), .A3(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n773), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n845), .B1(new_n858), .B2(G113gat), .ZN(new_n859));
  AOI211_X1 g658(.A(KEYINPUT116), .B(new_n380), .C1(new_n857), .C2(new_n773), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n844), .B1(new_n859), .B2(new_n860), .ZN(G1340gat));
  AOI21_X1  g660(.A(G120gat), .B1(new_n843), .B2(new_n370), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n369), .A2(new_n378), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n857), .B2(new_n863), .ZN(G1341gat));
  OAI21_X1  g663(.A(G127gat), .B1(new_n856), .B2(new_n838), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n843), .A2(new_n374), .A3(new_n318), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1342gat));
  NOR3_X1   g666(.A1(new_n842), .A2(G134gat), .A3(new_n269), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT56), .ZN(new_n869));
  OAI21_X1  g668(.A(G134gat), .B1(new_n856), .B2(new_n269), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(G1343gat));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n839), .A2(KEYINPUT57), .A3(new_n523), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n637), .A2(new_n855), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n268), .B1(new_n835), .B2(new_n830), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n838), .B1(new_n877), .B2(new_n828), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n523), .B1(new_n878), .B2(new_n809), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n876), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n873), .B1(new_n874), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n878), .A2(new_n809), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n524), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n875), .B1(new_n884), .B2(KEYINPUT57), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n880), .B(new_n524), .C1(new_n852), .C2(new_n810), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT117), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n882), .A2(new_n773), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(G141gat), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n729), .A2(new_n523), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n559), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n839), .A2(new_n891), .A3(new_n627), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n348), .A2(G141gat), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n872), .B1(new_n889), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n885), .A2(new_n886), .A3(new_n773), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(G141gat), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT58), .B1(new_n892), .B2(new_n893), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n898), .B1(new_n897), .B2(new_n899), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT119), .B1(new_n895), .B2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n904));
  AOI22_X1  g703(.A1(new_n888), .A2(G141gat), .B1(new_n892), .B2(new_n893), .ZN(new_n905));
  OAI221_X1 g704(.A(new_n904), .B1(new_n900), .B2(new_n901), .C1(new_n905), .C2(new_n872), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n903), .A2(new_n906), .ZN(G1344gat));
  NAND3_X1  g706(.A1(new_n892), .A2(new_n493), .A3(new_n370), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n877), .A2(new_n828), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n318), .B1(new_n910), .B2(KEYINPUT120), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n911), .B1(KEYINPUT120), .B2(new_n910), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n809), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n880), .A3(new_n524), .ZN(new_n914));
  OAI21_X1  g713(.A(KEYINPUT57), .B1(new_n839), .B2(new_n523), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n370), .A3(new_n876), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n909), .B1(new_n917), .B2(G148gat), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n882), .A2(new_n887), .ZN(new_n919));
  AOI211_X1 g718(.A(KEYINPUT59), .B(new_n493), .C1(new_n919), .C2(new_n370), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n908), .B1(new_n918), .B2(new_n920), .ZN(G1345gat));
  NAND3_X1  g720(.A1(new_n892), .A2(new_n497), .A3(new_n318), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n919), .A2(new_n318), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(new_n497), .ZN(G1346gat));
  AOI21_X1  g723(.A(G162gat), .B1(new_n892), .B2(new_n268), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n269), .A2(new_n498), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n919), .B2(new_n926), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n839), .A2(new_n678), .ZN(new_n928));
  INV_X1    g727(.A(new_n620), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n560), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT121), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(G169gat), .B1(new_n932), .B2(new_n773), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n678), .A2(new_n559), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n764), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT122), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n854), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n348), .A2(new_n408), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n933), .B1(new_n937), .B2(new_n938), .ZN(G1348gat));
  NAND3_X1  g738(.A1(new_n932), .A2(new_n409), .A3(new_n370), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n937), .A2(new_n370), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(new_n409), .ZN(G1349gat));
  NOR2_X1   g741(.A1(new_n838), .A2(new_n432), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n932), .A2(new_n943), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n854), .A2(new_n318), .A3(new_n936), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n945), .A2(KEYINPUT123), .ZN(new_n946));
  OAI21_X1  g745(.A(G183gat), .B1(new_n945), .B2(KEYINPUT123), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT60), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT60), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n950), .B(new_n944), .C1(new_n946), .C2(new_n947), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1350gat));
  NAND3_X1  g751(.A1(new_n932), .A2(new_n433), .A3(new_n268), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n268), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(G190gat), .ZN(new_n956));
  AOI211_X1 g755(.A(KEYINPUT61), .B(new_n433), .C1(new_n937), .C2(new_n268), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n953), .B1(new_n956), .B2(new_n957), .ZN(G1351gat));
  NAND2_X1  g757(.A1(new_n890), .A2(new_n560), .ZN(new_n959));
  XOR2_X1   g758(.A(new_n959), .B(KEYINPUT124), .Z(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(new_n928), .ZN(new_n961));
  XNOR2_X1  g760(.A(KEYINPUT125), .B(G197gat), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n961), .A2(new_n348), .A3(new_n963), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT126), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n637), .A2(new_n934), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n916), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n963), .B1(new_n967), .B2(new_n348), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n965), .A2(new_n968), .ZN(G1352gat));
  NOR3_X1   g768(.A1(new_n961), .A2(G204gat), .A3(new_n369), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n970), .B(KEYINPUT62), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n916), .A2(new_n370), .A3(new_n966), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(G204gat), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n973), .ZN(G1353gat));
  NAND4_X1  g773(.A1(new_n914), .A2(new_n318), .A3(new_n915), .A4(new_n966), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(G211gat), .ZN(new_n976));
  OR2_X1    g775(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n977));
  NAND2_X1  g776(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(new_n961), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n980), .A2(new_n478), .A3(new_n318), .ZN(new_n981));
  OAI211_X1 g780(.A(new_n979), .B(new_n981), .C1(new_n976), .C2(new_n977), .ZN(G1354gat));
  OAI21_X1  g781(.A(G218gat), .B1(new_n967), .B2(new_n269), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n980), .A2(new_n479), .A3(new_n268), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(G1355gat));
endmodule


