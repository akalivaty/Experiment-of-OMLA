//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1272, new_n1273,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT64), .Z(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  NAND4_X1  g0017(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n210), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT65), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT1), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AND2_X1   g0022(.A1(new_n220), .A2(new_n221), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR3_X1   g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR4_X1   g0027(.A1(new_n213), .A2(new_n222), .A3(new_n223), .A4(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT66), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT67), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n233), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT69), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G351));
  NAND3_X1  g0048(.A1(new_n206), .A2(KEYINPUT6), .A3(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT82), .ZN(new_n250));
  AND2_X1   g0050(.A1(G97), .A2(G107), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G97), .A2(G107), .ZN(new_n252));
  OAI21_X1  g0052(.A(KEYINPUT83), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT83), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G97), .A2(G107), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n207), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT6), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n253), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n225), .B1(new_n250), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT7), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n260), .B1(new_n261), .B2(G20), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n206), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n225), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G77), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR3_X1   g0071(.A1(new_n259), .A2(new_n267), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT71), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g0075(.A1(KEYINPUT71), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(new_n226), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G1), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G13), .A3(G20), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n275), .A2(new_n226), .A3(new_n276), .A4(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n268), .A2(G1), .ZN(new_n282));
  OAI21_X1  g0082(.A(G97), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT84), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n280), .A2(new_n205), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n284), .B1(new_n283), .B2(new_n285), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n272), .A2(new_n278), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n290));
  OAI211_X1 g0090(.A(G250), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G283), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  OAI211_X1 g0093(.A(G244), .B(new_n293), .C1(new_n263), .C2(new_n264), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT4), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n291), .B(new_n292), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n294), .A2(new_n295), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n290), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G274), .ZN(new_n299));
  INV_X1    g0099(.A(new_n226), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G41), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G45), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(G1), .ZN(new_n304));
  XNOR2_X1  g0104(.A(KEYINPUT5), .B(G41), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AND2_X1   g0106(.A1(KEYINPUT5), .A2(G41), .ZN(new_n307));
  NOR2_X1   g0107(.A1(KEYINPUT5), .A2(G41), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n304), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n301), .A2(G1), .A3(G13), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n309), .A2(G257), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n298), .A2(new_n306), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G179), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n298), .A2(new_n316), .A3(new_n306), .A4(new_n312), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT86), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n294), .A2(new_n295), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n261), .A2(KEYINPUT4), .A3(G244), .A4(new_n293), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n319), .A2(new_n320), .A3(new_n291), .A4(new_n292), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n311), .B1(new_n321), .B2(new_n290), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT86), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n322), .A2(new_n323), .A3(new_n316), .A4(new_n306), .ZN(new_n324));
  AND4_X1   g0124(.A1(new_n289), .A2(new_n315), .A3(new_n318), .A4(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G190), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n298), .A2(new_n326), .A3(new_n306), .A4(new_n312), .ZN(new_n327));
  NOR3_X1   g0127(.A1(new_n309), .A2(new_n290), .A3(new_n299), .ZN(new_n328));
  AOI211_X1 g0128(.A(new_n328), .B(new_n311), .C1(new_n321), .C2(new_n290), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n327), .B1(new_n329), .B2(G200), .ZN(new_n330));
  INV_X1    g0130(.A(new_n271), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT7), .B1(new_n265), .B2(new_n225), .ZN(new_n332));
  NOR4_X1   g0132(.A1(new_n263), .A2(new_n264), .A3(new_n260), .A4(G20), .ZN(new_n333));
  OAI21_X1  g0133(.A(G107), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n250), .A2(new_n258), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n331), .B(new_n334), .C1(new_n335), .C2(new_n225), .ZN(new_n336));
  INV_X1    g0136(.A(new_n288), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n336), .A2(new_n277), .B1(new_n337), .B2(new_n286), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n330), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT85), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT85), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n330), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n325), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT73), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(KEYINPUT10), .ZN(new_n345));
  INV_X1    g0145(.A(G41), .ZN(new_n346));
  AOI21_X1  g0146(.A(G1), .B1(new_n346), .B2(new_n303), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(new_n310), .A3(G274), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n279), .B1(G41), .B2(G45), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n310), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G226), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n348), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n261), .A2(G222), .A3(new_n293), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n354), .A2(KEYINPUT70), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(KEYINPUT70), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n261), .A2(G1698), .ZN(new_n358));
  INV_X1    g0158(.A(G223), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n358), .A2(new_n359), .B1(new_n270), .B2(new_n261), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g0161(.A(G190), .B(new_n353), .C1(new_n361), .C2(new_n310), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n357), .A2(new_n360), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n352), .B1(new_n363), .B2(new_n290), .ZN(new_n364));
  INV_X1    g0164(.A(G200), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n367));
  INV_X1    g0167(.A(G150), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n225), .A2(G33), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT8), .B(G58), .ZN(new_n370));
  OAI221_X1 g0170(.A(new_n367), .B1(new_n368), .B2(new_n269), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n280), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n371), .A2(new_n277), .B1(new_n201), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n281), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n279), .A2(G20), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(G50), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT9), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT9), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n344), .A2(KEYINPUT10), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n345), .B1(new_n366), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n383), .ZN(new_n385));
  INV_X1    g0185(.A(new_n345), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n361), .A2(new_n310), .ZN(new_n387));
  OAI21_X1  g0187(.A(G200), .B1(new_n387), .B2(new_n352), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n385), .A2(new_n386), .A3(new_n388), .A4(new_n362), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n364), .A2(new_n316), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n314), .B1(new_n387), .B2(new_n352), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n377), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n384), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n370), .B1(new_n279), .B2(G20), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n374), .A2(new_n394), .B1(new_n372), .B2(new_n370), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(G68), .B1(new_n332), .B2(new_n333), .ZN(new_n397));
  INV_X1    g0197(.A(G159), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT80), .B1(new_n269), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(G20), .A2(G33), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT80), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(new_n401), .A3(G159), .ZN(new_n402));
  XNOR2_X1  g0202(.A(G58), .B(G68), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n399), .A2(new_n402), .B1(G20), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n397), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n278), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n397), .A2(KEYINPUT16), .A3(new_n404), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n396), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT81), .ZN(new_n410));
  NOR2_X1   g0210(.A1(G223), .A2(G1698), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(new_n351), .B2(G1698), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n412), .A2(new_n261), .B1(G33), .B2(G87), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n410), .B1(new_n413), .B2(new_n310), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n359), .A2(new_n293), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n351), .A2(G1698), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n415), .B(new_n416), .C1(new_n263), .C2(new_n264), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G87), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n310), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT81), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n310), .A2(G232), .A3(new_n349), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n348), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(G179), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n414), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n314), .B1(new_n419), .B2(new_n422), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT18), .B1(new_n409), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(G68), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(new_n262), .B2(new_n266), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n399), .A2(new_n402), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n403), .A2(G20), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n406), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n433), .A2(new_n408), .A3(new_n277), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n395), .ZN(new_n435));
  INV_X1    g0235(.A(new_n426), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT18), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n427), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n422), .A2(G190), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n414), .A2(new_n420), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n365), .B1(new_n419), .B2(new_n422), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n409), .A2(KEYINPUT17), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n434), .A3(new_n395), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT17), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n439), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n261), .A2(G232), .A3(new_n293), .ZN(new_n450));
  INV_X1    g0250(.A(G238), .ZN(new_n451));
  OAI221_X1 g0251(.A(new_n450), .B1(new_n206), .B2(new_n261), .C1(new_n451), .C2(new_n358), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n290), .ZN(new_n453));
  INV_X1    g0253(.A(new_n350), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n454), .A2(G244), .B1(new_n302), .B2(new_n347), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n314), .ZN(new_n457));
  INV_X1    g0257(.A(new_n370), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n458), .A2(new_n400), .B1(G20), .B2(G77), .ZN(new_n459));
  XNOR2_X1  g0259(.A(KEYINPUT15), .B(G87), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n460), .B2(new_n369), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n461), .A2(new_n277), .B1(new_n270), .B2(new_n372), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n374), .A2(G77), .A3(new_n375), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT72), .B1(new_n457), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n453), .A2(new_n316), .A3(new_n455), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n457), .A2(new_n464), .A3(KEYINPUT72), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n464), .B1(new_n456), .B2(G200), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n470), .B1(new_n326), .B2(new_n456), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n449), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n393), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n348), .B1(new_n350), .B2(new_n451), .ZN(new_n474));
  OAI211_X1 g0274(.A(G232), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT74), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n261), .A2(KEYINPUT74), .A3(G232), .A4(G1698), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G97), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n261), .A2(G226), .A3(new_n293), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n477), .A2(new_n478), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n474), .B1(new_n481), .B2(new_n290), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT13), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI211_X1 g0284(.A(KEYINPUT13), .B(new_n474), .C1(new_n481), .C2(new_n290), .ZN(new_n485));
  OAI21_X1  g0285(.A(G169), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT14), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n481), .A2(new_n290), .ZN(new_n488));
  INV_X1    g0288(.A(new_n474), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT13), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n488), .A2(new_n483), .A3(new_n489), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT14), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(new_n494), .A3(G169), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT79), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT75), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n482), .A2(new_n497), .A3(new_n483), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n497), .B1(new_n482), .B2(new_n483), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n316), .B1(new_n490), .B2(KEYINPUT13), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n496), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n492), .A2(KEYINPUT75), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n482), .A2(new_n497), .A3(new_n483), .ZN(new_n504));
  AND4_X1   g0304(.A1(new_n496), .A2(new_n501), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n487), .B(new_n495), .C1(new_n502), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n372), .A2(new_n428), .ZN(new_n507));
  XNOR2_X1  g0307(.A(new_n507), .B(KEYINPUT12), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n375), .A2(G68), .ZN(new_n509));
  OR2_X1    g0309(.A1(new_n281), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n400), .A2(G50), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT76), .ZN(new_n512));
  XNOR2_X1  g0312(.A(new_n511), .B(new_n512), .ZN(new_n513));
  OAI22_X1  g0313(.A1(new_n369), .A2(new_n270), .B1(new_n225), .B2(G68), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n277), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  XOR2_X1   g0315(.A(KEYINPUT77), .B(KEYINPUT11), .Z(new_n516));
  AND2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n515), .A2(new_n516), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n508), .B(new_n510), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n506), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n503), .A2(new_n491), .A3(G190), .A4(new_n504), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(G200), .B1(new_n484), .B2(new_n485), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n508), .A2(new_n510), .ZN(new_n524));
  INV_X1    g0324(.A(new_n518), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n515), .A2(new_n516), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT78), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT78), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n521), .A2(new_n530), .A3(new_n527), .A4(new_n523), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n473), .A2(new_n520), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT21), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT20), .ZN(new_n536));
  AOI21_X1  g0336(.A(G20), .B1(G33), .B2(G283), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n268), .A2(G97), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT88), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n539), .B1(new_n537), .B2(new_n538), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n225), .A2(G116), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n277), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n536), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n276), .A2(new_n226), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n543), .B1(new_n547), .B2(new_n275), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n292), .B(new_n225), .C1(G33), .C2(new_n205), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT88), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n548), .A2(new_n552), .A3(KEYINPUT20), .ZN(new_n553));
  OAI21_X1  g0353(.A(G116), .B1(new_n281), .B2(new_n282), .ZN(new_n554));
  INV_X1    g0354(.A(G116), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n280), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n546), .A2(new_n553), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(G264), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n558));
  OAI211_X1 g0358(.A(G257), .B(new_n293), .C1(new_n263), .C2(new_n264), .ZN(new_n559));
  OR2_X1    g0359(.A1(KEYINPUT3), .A2(G33), .ZN(new_n560));
  NAND2_X1  g0360(.A1(KEYINPUT3), .A2(G33), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(G303), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n558), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n563), .A2(new_n290), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n309), .A2(new_n310), .ZN(new_n565));
  INV_X1    g0365(.A(G270), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n306), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(G169), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n535), .B1(new_n557), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n554), .A2(new_n556), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n548), .A2(new_n552), .A3(KEYINPUT20), .ZN(new_n571));
  AOI21_X1  g0371(.A(KEYINPUT20), .B1(new_n548), .B2(new_n552), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR3_X1   g0373(.A1(new_n564), .A2(new_n567), .A3(new_n316), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n290), .B1(new_n304), .B2(new_n305), .ZN(new_n576));
  INV_X1    g0376(.A(new_n309), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n576), .A2(G270), .B1(new_n577), .B2(new_n302), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n563), .A2(new_n290), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n314), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n573), .A2(KEYINPUT21), .A3(new_n580), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n569), .A2(new_n575), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n564), .A2(new_n567), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G190), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n584), .B(new_n557), .C1(new_n365), .C2(new_n583), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n309), .A2(G264), .A3(new_n310), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n306), .A2(new_n588), .ZN(new_n589));
  OR2_X1    g0389(.A1(G250), .A2(G1698), .ZN(new_n590));
  INV_X1    g0390(.A(G257), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G1698), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n590), .B(new_n592), .C1(new_n263), .C2(new_n264), .ZN(new_n593));
  NAND2_X1  g0393(.A1(G33), .A2(G294), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n310), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n314), .B1(new_n589), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n593), .A2(new_n594), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n290), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n598), .A2(new_n316), .A3(new_n306), .A4(new_n588), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT23), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(new_n206), .A3(G20), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n225), .A2(G33), .A3(G116), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT23), .B1(new_n225), .B2(G107), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT90), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT90), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n608), .B(KEYINPUT23), .C1(new_n225), .C2(G107), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n605), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT22), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n225), .A2(KEYINPUT89), .A3(G87), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n261), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n611), .B1(new_n261), .B2(new_n612), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n610), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT24), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT24), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n610), .B(new_n617), .C1(new_n613), .C2(new_n614), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n278), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n372), .A2(new_n206), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n620), .B(KEYINPUT25), .ZN(new_n621));
  INV_X1    g0421(.A(new_n282), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n547), .A2(new_n275), .A3(new_n280), .A4(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n623), .A2(new_n206), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n601), .B1(new_n619), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT91), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n261), .A2(G244), .A3(G1698), .ZN(new_n629));
  NAND2_X1  g0429(.A1(G33), .A2(G116), .ZN(new_n630));
  OAI211_X1 g0430(.A(G238), .B(new_n293), .C1(new_n263), .C2(new_n264), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n290), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n302), .A2(new_n304), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT87), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n303), .B2(G1), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n279), .A2(KEYINPUT87), .A3(G45), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n310), .A2(new_n636), .A3(G250), .A4(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n633), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G200), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n639), .B1(new_n290), .B2(new_n632), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(G190), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT19), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n225), .B1(new_n479), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(G87), .B2(new_n207), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n645), .B1(new_n369), .B2(new_n205), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n225), .B(G68), .C1(new_n263), .C2(new_n264), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n277), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n374), .A2(G87), .A3(new_n622), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n460), .A2(new_n372), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n642), .A2(new_n644), .A3(new_n654), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n651), .B(new_n653), .C1(new_n623), .C2(new_n460), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n633), .A2(new_n640), .A3(new_n316), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n656), .B(new_n657), .C1(G169), .C2(new_n643), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT91), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n601), .B(new_n660), .C1(new_n619), .C2(new_n626), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n598), .A2(G190), .A3(new_n306), .A4(new_n588), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n589), .A2(new_n595), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n662), .B1(new_n663), .B2(new_n365), .ZN(new_n664));
  OR3_X1    g0464(.A1(new_n619), .A2(new_n664), .A3(new_n626), .ZN(new_n665));
  AND4_X1   g0465(.A1(new_n628), .A2(new_n659), .A3(new_n661), .A4(new_n665), .ZN(new_n666));
  AND4_X1   g0466(.A1(new_n343), .A2(new_n534), .A3(new_n587), .A4(new_n666), .ZN(G372));
  NOR2_X1   g0467(.A1(new_n522), .A2(new_n528), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n520), .B1(new_n668), .B2(new_n469), .ZN(new_n669));
  INV_X1    g0469(.A(new_n448), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n439), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n384), .A2(new_n389), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n392), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT92), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n582), .A2(new_n675), .A3(new_n627), .ZN(new_n676));
  INV_X1    g0476(.A(new_n627), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n569), .A2(new_n581), .A3(new_n575), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT92), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n655), .A2(new_n658), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n619), .A2(new_n664), .A3(new_n626), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n289), .A2(new_n318), .A3(new_n315), .A4(new_n324), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n330), .A2(new_n338), .A3(new_n341), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n341), .B1(new_n330), .B2(new_n338), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n683), .B(new_n684), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n680), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n684), .A2(new_n681), .ZN(new_n689));
  XOR2_X1   g0489(.A(KEYINPUT93), .B(KEYINPUT26), .Z(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT26), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n691), .B(new_n658), .C1(new_n692), .C2(new_n689), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n534), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n674), .A2(new_n695), .ZN(G369));
  NAND3_X1  g0496(.A1(new_n279), .A2(new_n225), .A3(G13), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n697), .A2(KEYINPUT27), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(KEYINPUT27), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(new_n699), .A3(G213), .ZN(new_n700));
  INV_X1    g0500(.A(G343), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n557), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT94), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n704), .B1(new_n586), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n705), .B2(new_n586), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n582), .A2(new_n704), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(G330), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n628), .A2(new_n665), .A3(new_n661), .ZN(new_n711));
  INV_X1    g0511(.A(new_n619), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n703), .B1(new_n712), .B2(new_n625), .ZN(new_n713));
  OAI22_X1  g0513(.A1(new_n711), .A2(new_n713), .B1(new_n627), .B2(new_n703), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n678), .A2(new_n703), .ZN(new_n716));
  OAI22_X1  g0516(.A1(new_n711), .A2(new_n716), .B1(new_n627), .B2(new_n702), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n715), .A2(new_n718), .ZN(G399));
  NAND2_X1  g0519(.A1(new_n211), .A2(new_n346), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G87), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n252), .A2(new_n722), .A3(new_n555), .ZN(new_n723));
  XOR2_X1   g0523(.A(new_n723), .B(KEYINPUT95), .Z(new_n724));
  NOR3_X1   g0524(.A1(new_n721), .A2(new_n279), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n224), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(new_n721), .ZN(new_n727));
  XOR2_X1   g0527(.A(new_n727), .B(KEYINPUT28), .Z(new_n728));
  NAND4_X1  g0528(.A1(new_n666), .A2(new_n343), .A3(new_n587), .A4(new_n703), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  INV_X1    g0530(.A(new_n574), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n322), .A2(new_n643), .A3(new_n663), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n643), .A2(new_n663), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n734), .A2(KEYINPUT30), .A3(new_n322), .A4(new_n574), .ZN(new_n735));
  INV_X1    g0535(.A(new_n583), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n663), .A2(G179), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n736), .A2(new_n737), .A3(new_n313), .A4(new_n641), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n733), .A2(new_n735), .A3(new_n738), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n702), .ZN(new_n740));
  AOI21_X1  g0540(.A(KEYINPUT31), .B1(new_n739), .B2(new_n702), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n729), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(KEYINPUT96), .A3(G330), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(KEYINPUT96), .B1(new_n743), .B2(G330), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT99), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n325), .A2(new_n692), .A3(new_n659), .ZN(new_n749));
  XOR2_X1   g0549(.A(new_n658), .B(KEYINPUT97), .Z(new_n750));
  INV_X1    g0550(.A(new_n690), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(new_n684), .B2(new_n681), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n340), .A2(new_n342), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n582), .A2(new_n628), .A3(new_n661), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n754), .A2(new_n755), .A3(new_n684), .A4(new_n683), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT98), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n343), .A2(KEYINPUT98), .A3(new_n683), .A4(new_n755), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n748), .B(new_n702), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n755), .A2(new_n683), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n757), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n753), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n763), .A2(new_n759), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(KEYINPUT99), .B1(new_n765), .B2(new_n703), .ZN(new_n766));
  OAI21_X1  g0566(.A(KEYINPUT29), .B1(new_n760), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n694), .A2(new_n703), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT29), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n747), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n728), .B1(new_n771), .B2(G1), .ZN(G364));
  AND2_X1   g0572(.A1(new_n225), .A2(G13), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n279), .B1(new_n773), .B2(G45), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n721), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n710), .A2(new_n776), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n707), .A2(new_n708), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G330), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G13), .A2(G33), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n778), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n776), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n226), .B1(G20), .B2(new_n314), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n211), .A2(new_n261), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT100), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G355), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(G116), .B2(new_n211), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n791), .A2(KEYINPUT101), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n247), .A2(G45), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n211), .A2(new_n265), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(new_n303), .B2(new_n726), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n791), .A2(KEYINPUT101), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n783), .B(new_n787), .C1(new_n792), .C2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n225), .A2(G179), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n798), .A2(new_n326), .A3(G200), .ZN(new_n799));
  INV_X1    g0599(.A(G283), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n225), .A2(new_n316), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G200), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(G190), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  XOR2_X1   g0605(.A(KEYINPUT33), .B(G317), .Z(new_n806));
  NAND3_X1  g0606(.A1(new_n798), .A2(G190), .A3(G200), .ZN(new_n807));
  INV_X1    g0607(.A(G303), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n805), .A2(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n803), .A2(new_n326), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n801), .B(new_n809), .C1(G326), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n365), .A2(G190), .ZN(new_n812));
  OAI21_X1  g0612(.A(G20), .B1(new_n812), .B2(G179), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT102), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(G294), .ZN(new_n819));
  NOR2_X1   g0619(.A1(G190), .A2(G200), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n798), .A2(new_n820), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n821), .A2(KEYINPUT103), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(KEYINPUT103), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(G329), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n812), .A2(new_n225), .A3(new_n316), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(G322), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n265), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n802), .A2(new_n820), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n830), .B1(G311), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n811), .A2(new_n819), .A3(new_n826), .A4(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n817), .A2(new_n205), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n261), .B1(new_n828), .B2(new_n202), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G77), .B2(new_n832), .ZN(new_n837));
  INV_X1    g0637(.A(new_n799), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n810), .A2(G50), .B1(new_n838), .B2(G107), .ZN(new_n839));
  INV_X1    g0639(.A(new_n807), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n804), .A2(G68), .B1(new_n840), .B2(G87), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n821), .A2(new_n398), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT32), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n837), .A2(new_n839), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n834), .B1(new_n835), .B2(new_n844), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n786), .B(new_n797), .C1(new_n787), .C2(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n777), .A2(new_n780), .B1(new_n785), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G396));
  NOR2_X1   g0648(.A1(new_n787), .A2(new_n781), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n261), .B1(new_n832), .B2(G116), .ZN(new_n851));
  INV_X1    g0651(.A(G294), .ZN(new_n852));
  INV_X1    g0652(.A(G311), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n851), .B1(new_n852), .B2(new_n828), .C1(new_n824), .C2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n810), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n855), .A2(new_n808), .B1(new_n799), .B2(new_n722), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n805), .A2(new_n800), .B1(new_n807), .B2(new_n206), .ZN(new_n857));
  NOR4_X1   g0657(.A1(new_n854), .A2(new_n835), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(G132), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n261), .B1(new_n824), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n799), .A2(new_n428), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(G50), .B2(new_n840), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT104), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n860), .B(new_n863), .C1(G58), .C2(new_n818), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n832), .A2(G159), .B1(new_n827), .B2(G143), .ZN(new_n865));
  INV_X1    g0665(.A(G137), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n865), .B1(new_n855), .B2(new_n866), .C1(new_n368), .C2(new_n805), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT34), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n858), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n787), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n776), .B1(G77), .B2(new_n850), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n871), .B(KEYINPUT105), .Z(new_n872));
  NAND2_X1  g0672(.A1(new_n464), .A2(new_n702), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n469), .A2(new_n471), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n468), .A2(new_n467), .ZN(new_n875));
  OR3_X1    g0675(.A1(new_n875), .A2(new_n465), .A3(new_n873), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n877), .A2(new_n782), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n877), .B(KEYINPUT106), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n768), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n703), .B(new_n877), .C1(new_n688), .C2(new_n693), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n747), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n883), .A2(new_n776), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n747), .A2(new_n881), .A3(new_n882), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n879), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(G384));
  AOI21_X1  g0687(.A(new_n533), .B1(new_n768), .B2(new_n769), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n673), .B1(new_n767), .B2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT109), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n439), .A2(new_n700), .ZN(new_n891));
  INV_X1    g0691(.A(new_n520), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n703), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n435), .A2(new_n436), .ZN(new_n894));
  INV_X1    g0694(.A(new_n700), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n435), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n894), .A2(new_n896), .A3(new_n445), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT37), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT37), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n894), .A2(new_n896), .A3(new_n899), .A4(new_n445), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n896), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n439), .B2(new_n448), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n901), .A2(new_n903), .A3(KEYINPUT38), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n901), .B2(new_n903), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT39), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n901), .A2(new_n903), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT38), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n901), .A2(new_n903), .A3(KEYINPUT38), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT39), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n907), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n495), .A2(new_n487), .ZN(new_n916));
  INV_X1    g0716(.A(new_n505), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n501), .A2(new_n503), .A3(new_n504), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT79), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n916), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n532), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n527), .A2(new_n703), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n922), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n522), .B2(new_n528), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n506), .B2(new_n519), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n469), .A2(new_n702), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT107), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT108), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n882), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n931), .B1(new_n882), .B2(new_n930), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n928), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n891), .B1(new_n893), .B2(new_n915), .C1(new_n934), .C2(new_n906), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n890), .B(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n743), .B1(new_n904), .B2(new_n905), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n924), .B1(new_n920), .B2(new_n532), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n877), .B1(new_n938), .B2(new_n926), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT110), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT40), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g0742(.A(KEYINPUT110), .B(KEYINPUT40), .C1(new_n937), .C2(new_n939), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n944), .A2(new_n534), .A3(new_n743), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n944), .B1(new_n534), .B2(new_n743), .ZN(new_n946));
  INV_X1    g0746(.A(G330), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n936), .A2(new_n948), .B1(new_n279), .B2(new_n773), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n936), .B2(new_n948), .ZN(new_n950));
  INV_X1    g0750(.A(new_n335), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(KEYINPUT35), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(KEYINPUT35), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n226), .A2(new_n225), .A3(new_n555), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT36), .Z(new_n956));
  OAI211_X1 g0756(.A(new_n726), .B(G77), .C1(new_n202), .C2(new_n428), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n201), .A2(G68), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n279), .B(G13), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  NOR3_X1   g0759(.A1(new_n950), .A2(new_n956), .A3(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT111), .Z(G367));
  AND3_X1   g0761(.A1(new_n232), .A2(new_n211), .A3(new_n265), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n783), .A2(new_n787), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n211), .B2(new_n460), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n831), .A2(new_n201), .B1(new_n821), .B2(new_n866), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n265), .B(new_n965), .C1(G150), .C2(new_n827), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n818), .A2(G68), .ZN(new_n967));
  AOI22_X1  g0767(.A1(G143), .A2(new_n810), .B1(new_n804), .B2(G159), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n799), .A2(new_n270), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(G58), .B2(new_n840), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n966), .A2(new_n967), .A3(new_n968), .A4(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n821), .ZN(new_n972));
  AOI22_X1  g0772(.A1(G283), .A2(new_n832), .B1(new_n972), .B2(G317), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n840), .A2(KEYINPUT46), .A3(G116), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT46), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n807), .B2(new_n555), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n261), .B1(new_n827), .B2(G303), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n973), .A2(new_n974), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n799), .A2(new_n205), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(G311), .B2(new_n810), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(new_n852), .B2(new_n805), .C1(new_n817), .C2(new_n206), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n971), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT47), .Z(new_n983));
  OAI221_X1 g0783(.A(new_n776), .B1(new_n962), .B2(new_n964), .C1(new_n983), .C2(new_n870), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT114), .Z(new_n985));
  OR2_X1    g0785(.A1(new_n654), .A2(new_n703), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n659), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT112), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n986), .A2(new_n658), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n659), .A2(KEYINPUT112), .A3(new_n986), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n783), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n985), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n715), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT45), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n338), .A2(new_n703), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n762), .A2(new_n998), .B1(new_n684), .B2(new_n703), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n997), .B1(new_n1000), .B2(new_n717), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n718), .A2(new_n999), .A3(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1000), .A2(KEYINPUT44), .A3(new_n717), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT44), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n718), .B2(new_n999), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n996), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n715), .A2(new_n1003), .A3(new_n1007), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n711), .A2(new_n716), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n716), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1013), .B1(new_n714), .B2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n709), .B(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n771), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n720), .B(KEYINPUT41), .Z(new_n1018));
  AOI21_X1  g0818(.A(new_n775), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n999), .A2(new_n1012), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT42), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n992), .A2(KEYINPUT113), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT43), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n992), .A2(KEYINPUT113), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n340), .A2(new_n342), .B1(new_n628), .B2(new_n661), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n703), .B1(new_n1028), .B2(new_n325), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1022), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1022), .A2(new_n1029), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1026), .B1(new_n1024), .B2(new_n993), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n996), .A2(new_n999), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1033), .B(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n995), .B1(new_n1019), .B2(new_n1035), .ZN(G387));
  INV_X1    g0836(.A(new_n1016), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n714), .A2(new_n784), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n238), .A2(new_n303), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n370), .A2(G50), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT50), .ZN(new_n1041));
  AOI211_X1 g0841(.A(G45), .B(new_n724), .C1(G68), .C2(G77), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n794), .B(new_n1039), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n789), .A2(new_n724), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(G107), .B2(new_n211), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n963), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n776), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n828), .A2(new_n201), .B1(new_n831), .B2(new_n428), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n265), .B(new_n1048), .C1(G150), .C2(new_n972), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n817), .A2(new_n460), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n979), .B1(G159), .B2(new_n810), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n804), .A2(new_n458), .B1(new_n840), .B2(G77), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n853), .A2(new_n805), .B1(new_n855), .B2(new_n829), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1054), .A2(KEYINPUT115), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(KEYINPUT115), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n832), .A2(G303), .B1(new_n827), .B2(G317), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT48), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n817), .A2(new_n800), .B1(new_n852), .B2(new_n807), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1060), .A2(KEYINPUT49), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n261), .B1(new_n972), .B2(G326), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(new_n555), .C2(new_n799), .ZN(new_n1065));
  AOI21_X1  g0865(.A(KEYINPUT49), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1053), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1047), .B1(new_n1067), .B2(new_n787), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1037), .A2(new_n775), .B1(new_n1038), .B2(new_n1068), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n771), .A2(new_n1037), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n720), .B1(new_n771), .B2(new_n1037), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT116), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1016), .B(new_n747), .C1(new_n767), .C2(new_n770), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n1074), .A2(KEYINPUT116), .A3(new_n720), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1069), .B1(new_n1073), .B2(new_n1075), .ZN(G393));
  INV_X1    g0876(.A(new_n1074), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n721), .B1(new_n1077), .B2(new_n1011), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1074), .B1(new_n1010), .B2(new_n1009), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1011), .A2(new_n774), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1000), .A2(new_n783), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n243), .A2(new_n211), .A3(new_n265), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n963), .B1(new_n211), .B2(new_n205), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n776), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n818), .A2(G77), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n832), .A2(new_n458), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n265), .B1(new_n972), .B2(G143), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n428), .A2(new_n807), .B1(new_n799), .B2(new_n722), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G50), .B2(new_n804), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .A4(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n810), .A2(G150), .B1(G159), .B2(new_n827), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT51), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n810), .A2(G317), .B1(G311), .B2(new_n827), .ZN(new_n1094));
  XOR2_X1   g0894(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n1095));
  XNOR2_X1  g0895(.A(new_n1094), .B(new_n1095), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n206), .A2(new_n799), .B1(new_n807), .B2(new_n800), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G303), .B2(new_n804), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n265), .B1(new_n831), .B2(new_n852), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(G322), .B2(new_n972), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1098), .B(new_n1100), .C1(new_n555), .C2(new_n817), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n1091), .A2(new_n1093), .B1(new_n1096), .B2(new_n1101), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT118), .Z(new_n1103));
  AOI21_X1  g0903(.A(new_n1085), .B1(new_n1103), .B2(new_n787), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1081), .B1(new_n1082), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1080), .A2(new_n1105), .ZN(G390));
  NAND2_X1  g0906(.A1(new_n743), .A2(G330), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n939), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n912), .A2(new_n893), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n877), .B1(new_n760), .B2(new_n766), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n929), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1109), .B1(new_n1112), .B2(new_n928), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n934), .A2(new_n893), .B1(new_n914), .B2(new_n907), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1108), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n928), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n882), .A2(new_n930), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(KEYINPUT108), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n882), .A2(new_n930), .A3(new_n931), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1116), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n893), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n915), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT96), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1107), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1124), .A2(new_n744), .A3(new_n877), .A4(new_n928), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1116), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1122), .B(new_n1125), .C1(new_n1126), .C2(new_n1109), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1115), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n767), .A2(new_n888), .ZN(new_n1129));
  OR2_X1    g0929(.A1(new_n533), .A2(new_n1107), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1129), .A2(new_n674), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(KEYINPUT119), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT119), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n889), .A2(new_n1133), .A3(new_n1130), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n932), .A2(new_n933), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1124), .A2(new_n744), .A3(new_n877), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1108), .B1(new_n1136), .B2(new_n1116), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1116), .B1(new_n880), .B2(new_n1107), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1125), .A2(new_n1138), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1135), .A2(new_n1137), .B1(new_n1112), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1132), .A2(new_n1134), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n720), .B1(new_n1128), .B2(new_n1141), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1132), .A2(new_n1134), .A3(new_n1140), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1143), .A2(new_n1127), .A3(new_n1115), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n915), .A2(new_n781), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n776), .B1(new_n458), .B2(new_n850), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n206), .A2(new_n805), .B1(new_n855), .B2(new_n800), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n861), .B(new_n1148), .C1(G87), .C2(new_n840), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n825), .A2(G294), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n265), .B1(new_n828), .B2(new_n555), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G97), .B2(new_n832), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1149), .A2(new_n1086), .A3(new_n1150), .A4(new_n1152), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n805), .A2(new_n866), .B1(new_n799), .B2(new_n201), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G128), .B2(new_n810), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n825), .A2(G125), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n827), .A2(G132), .ZN(new_n1157));
  XOR2_X1   g0957(.A(KEYINPUT54), .B(G143), .Z(new_n1158));
  AOI21_X1  g0958(.A(new_n265), .B1(new_n832), .B2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .A4(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n807), .A2(new_n368), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1161), .B(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n398), .B2(new_n817), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1153), .B1(new_n1160), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1147), .B1(new_n1165), .B2(new_n787), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1146), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1128), .B2(new_n774), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1145), .A2(new_n1169), .ZN(G378));
  NAND2_X1  g0970(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1115), .A2(new_n1127), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1171), .B1(new_n1172), .B2(new_n1143), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n378), .A2(new_n700), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n393), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1174), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n384), .A2(new_n389), .A3(new_n392), .A4(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1175), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1178), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n944), .B2(G330), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n947), .B(new_n1181), .C1(new_n942), .C2(new_n943), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n935), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n928), .A2(new_n912), .A3(new_n743), .A4(new_n877), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT40), .B1(new_n1186), .B2(KEYINPUT110), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n943), .ZN(new_n1188));
  OAI21_X1  g0988(.A(G330), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1181), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n891), .B1(new_n915), .B2(new_n893), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n1120), .B2(new_n912), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n944), .A2(G330), .A3(new_n1182), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1190), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT122), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1185), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n935), .B(KEYINPUT122), .C1(new_n1183), .C2(new_n1184), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(KEYINPUT57), .A3(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n721), .B1(new_n1173), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1112), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1139), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1136), .A2(new_n1116), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1108), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1135), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1200), .A2(new_n1201), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1134), .B(new_n1132), .C1(new_n1128), .C2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1185), .A2(new_n1194), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT57), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1199), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1181), .A2(new_n781), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n261), .A2(G41), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n460), .B2(new_n831), .C1(new_n828), .C2(new_n206), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G283), .B2(new_n825), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n804), .A2(G97), .B1(new_n840), .B2(G77), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n810), .A2(G116), .B1(new_n838), .B2(G58), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1214), .A2(new_n967), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT58), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n268), .A2(new_n346), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n201), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n827), .A2(G128), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n866), .B2(new_n831), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G132), .B2(new_n804), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n810), .A2(G125), .B1(new_n840), .B2(new_n1158), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(new_n368), .C2(new_n817), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1219), .B1(new_n972), .B2(G124), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1227), .B(new_n1228), .C1(new_n398), .C2(new_n799), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1218), .B1(new_n1212), .B2(new_n1220), .C1(new_n1226), .C2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT121), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n870), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n1231), .B2(new_n1230), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n849), .A2(new_n201), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1211), .A2(new_n776), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n1208), .B2(new_n775), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1210), .A2(new_n1237), .ZN(G375));
  OAI21_X1  g1038(.A(new_n776), .B1(G68), .B2(new_n850), .ZN(new_n1239));
  XOR2_X1   g1039(.A(new_n1239), .B(KEYINPUT123), .Z(new_n1240));
  NOR2_X1   g1040(.A1(new_n928), .A2(new_n782), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n855), .A2(new_n852), .B1(new_n807), .B2(new_n205), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n969), .B(new_n1242), .C1(G116), .C2(new_n804), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n825), .A2(G303), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n265), .B1(new_n831), .B2(new_n206), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G283), .B2(new_n827), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1243), .A2(new_n1050), .A3(new_n1244), .A4(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n825), .A2(G128), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n804), .A2(new_n1158), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n832), .A2(G150), .B1(new_n827), .B2(G137), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n810), .A2(G132), .B1(new_n840), .B2(G159), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n261), .B1(new_n799), .B2(new_n202), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1253), .A2(KEYINPUT124), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(KEYINPUT124), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1254), .B(new_n1255), .C1(new_n201), .C2(new_n817), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1247), .B1(new_n1252), .B2(new_n1256), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1240), .B(new_n1241), .C1(new_n787), .C2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1140), .B2(new_n775), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1141), .A2(new_n1018), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1140), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1259), .B1(new_n1260), .B2(new_n1261), .ZN(G381));
  NAND2_X1  g1062(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1263));
  OAI21_X1  g1063(.A(KEYINPUT116), .B1(new_n1074), .B2(new_n720), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n1264), .A3(new_n1070), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(new_n847), .A3(new_n1069), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(G381), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(G390), .ZN(new_n1268));
  INV_X1    g1068(.A(G387), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1267), .A2(new_n1268), .A3(new_n886), .A4(new_n1269), .ZN(new_n1270));
  OR3_X1    g1070(.A1(G375), .A2(G378), .A3(new_n1270), .ZN(G407));
  NAND2_X1  g1071(.A1(new_n701), .A2(G213), .ZN(new_n1272));
  OR3_X1    g1072(.A1(G375), .A2(G378), .A3(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(G407), .A2(new_n1273), .A3(G213), .ZN(G409));
  NOR2_X1   g1074(.A1(G393), .A2(G396), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n847), .B1(new_n1265), .B2(new_n1069), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1275), .A2(new_n1276), .A3(G387), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT125), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G387), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G393), .A2(G396), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1279), .B1(new_n1280), .B2(new_n1266), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1268), .B1(new_n1277), .B2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1280), .A2(new_n1269), .A3(new_n1266), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1284));
  OAI211_X1 g1084(.A(G390), .B(new_n1283), .C1(new_n1284), .C2(new_n1279), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1282), .A2(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(G378), .B(new_n1237), .C1(new_n1199), .C2(new_n1209), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1168), .B1(new_n1144), .B2(new_n1142), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1207), .A2(new_n1018), .A3(new_n1208), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1196), .A2(new_n775), .A3(new_n1197), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1235), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1288), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1287), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT62), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1141), .A2(KEYINPUT60), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1171), .A2(new_n1206), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1134), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1133), .B1(new_n889), .B2(new_n1130), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1206), .B(KEYINPUT60), .C1(new_n1298), .C2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1297), .A2(new_n721), .A3(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(G384), .B1(new_n1301), .B2(new_n1259), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1261), .B1(KEYINPUT60), .B2(new_n1141), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1300), .A2(new_n721), .ZN(new_n1304));
  OAI211_X1 g1104(.A(G384), .B(new_n1259), .C1(new_n1303), .C2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1302), .A2(new_n1306), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1293), .A2(new_n1294), .A3(new_n1272), .A4(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT61), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(new_n1287), .A2(new_n1292), .B1(G213), .B2(new_n701), .ZN(new_n1310));
  INV_X1    g1110(.A(G2897), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1272), .A2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1312), .B1(new_n1302), .B2(new_n1306), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1259), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n886), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1315), .B(new_n1305), .C1(new_n1311), .C2(new_n1272), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1313), .A2(new_n1316), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1308), .B(new_n1309), .C1(new_n1310), .C2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1294), .B1(new_n1310), .B2(new_n1307), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1286), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(KEYINPUT63), .B1(new_n1310), .B2(new_n1317), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1310), .A2(new_n1307), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1282), .A2(new_n1285), .A3(new_n1309), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(new_n1324), .B(KEYINPUT126), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1310), .A2(KEYINPUT63), .A3(new_n1307), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1323), .A2(new_n1325), .A3(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1320), .A2(new_n1327), .ZN(G405));
  NAND2_X1  g1128(.A1(G375), .A2(new_n1288), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1307), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1329), .A2(new_n1287), .A3(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(G378), .B1(new_n1210), .B2(new_n1237), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1287), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1307), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1331), .A2(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1335), .A2(KEYINPUT127), .A3(new_n1286), .ZN(new_n1336));
  OR2_X1    g1136(.A1(new_n1286), .A2(KEYINPUT127), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1286), .A2(KEYINPUT127), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1331), .A2(new_n1334), .A3(new_n1337), .A4(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1336), .A2(new_n1339), .ZN(G402));
endmodule


