//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G116), .A2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n206), .B(new_n207), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  AOI21_X1  g0010(.A(new_n210), .B1(G50), .B2(G226), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G107), .A2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G58), .ZN(new_n213));
  INV_X1    g0013(.A(G232), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n211), .B(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n205), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT65), .Z(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT64), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n224), .A2(G1), .A3(G13), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G20), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n205), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT0), .Z(new_n232));
  AND2_X1   g0032(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n233));
  NOR4_X1   g0033(.A1(new_n221), .A2(new_n229), .A3(new_n232), .A4(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n214), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT66), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G150), .ZN(new_n252));
  INV_X1    g0052(.A(G20), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT69), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XOR2_X1   g0056(.A(KEYINPUT8), .B(G58), .Z(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  OAI221_X1 g0058(.A(new_n252), .B1(new_n253), .B2(new_n201), .C1(new_n256), .C2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n223), .A2(new_n225), .A3(new_n260), .ZN(new_n261));
  AND3_X1   g0061(.A1(new_n223), .A2(new_n225), .A3(new_n260), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(G1), .B2(new_n253), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n259), .A2(new_n261), .B1(G50), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G13), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n266), .A2(new_n253), .A3(G1), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G50), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT3), .B(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G222), .A2(G1698), .ZN(new_n273));
  INV_X1    g0073(.A(G1698), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G223), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n272), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n277), .B1(new_n223), .B2(new_n225), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n276), .B(new_n278), .C1(G77), .C2(new_n272), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  INV_X1    g0080(.A(G45), .ZN(new_n281));
  AOI21_X1  g0081(.A(G1), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT68), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(new_n277), .B2(new_n222), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n285), .A2(KEYINPUT68), .A3(G1), .A4(G13), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n282), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G226), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n284), .A2(new_n286), .ZN(new_n289));
  INV_X1    g0089(.A(G274), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT67), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n290), .B1(new_n282), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G1), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(G41), .B2(G45), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT67), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n289), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n279), .A2(new_n288), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G179), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n271), .B(new_n300), .C1(G169), .C2(new_n298), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n265), .A2(KEYINPUT9), .A3(new_n270), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT70), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n303), .B(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n297), .A2(G200), .ZN(new_n306));
  XOR2_X1   g0106(.A(new_n306), .B(KEYINPUT71), .Z(new_n307));
  INV_X1    g0107(.A(KEYINPUT9), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n271), .A2(new_n308), .B1(G190), .B2(new_n298), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n305), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n305), .A2(new_n309), .A3(new_n312), .A4(new_n307), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n302), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(G58), .B(G68), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n315), .A2(G20), .B1(G159), .B2(new_n251), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT7), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n272), .A2(new_n317), .A3(G20), .ZN(new_n318));
  INV_X1    g0118(.A(G33), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT3), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G33), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT75), .ZN(new_n323));
  AND3_X1   g0123(.A1(new_n320), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n323), .B1(new_n320), .B2(new_n322), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n253), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n318), .B1(new_n326), .B2(new_n317), .ZN(new_n327));
  OAI211_X1 g0127(.A(KEYINPUT16), .B(new_n316), .C1(new_n327), .C2(new_n216), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT16), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n317), .B1(new_n272), .B2(G20), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n320), .A2(new_n322), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(KEYINPUT7), .A3(new_n253), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n216), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n316), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n329), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n328), .A2(new_n261), .A3(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n257), .A2(new_n267), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(new_n263), .B2(new_n257), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  OR2_X1    g0139(.A1(G223), .A2(G1698), .ZN(new_n340));
  INV_X1    g0140(.A(G226), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G1698), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n320), .A2(new_n340), .A3(new_n322), .A4(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G33), .A2(G87), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n278), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n289), .A2(G232), .A3(new_n294), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n296), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G200), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(G190), .B2(new_n348), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n336), .A2(new_n339), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT17), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n336), .A2(KEYINPUT17), .A3(new_n339), .A4(new_n351), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n348), .A2(G169), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n346), .A2(new_n296), .A3(new_n347), .A4(G179), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n358), .A2(KEYINPUT76), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT76), .B1(new_n358), .B2(new_n359), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n336), .A2(new_n339), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT77), .B(KEYINPUT18), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n362), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n362), .A2(new_n363), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n364), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n357), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  OR3_X1    g0170(.A1(new_n268), .A2(KEYINPUT12), .A3(G68), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT12), .B1(new_n268), .B2(G68), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n264), .A2(G68), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n251), .A2(G50), .ZN(new_n374));
  OAI221_X1 g0174(.A(new_n374), .B1(new_n253), .B2(G68), .C1(new_n256), .C2(new_n202), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT11), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n375), .A2(new_n376), .A3(new_n261), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n376), .B1(new_n375), .B2(new_n261), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n373), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT74), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n379), .B(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT14), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT72), .ZN(new_n383));
  NOR2_X1   g0183(.A1(G226), .A2(G1698), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n214), .B2(G1698), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n385), .A2(new_n272), .B1(G33), .B2(G97), .ZN(new_n386));
  INV_X1    g0186(.A(new_n278), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n383), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n214), .A2(G1698), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(G226), .B2(G1698), .ZN(new_n390));
  INV_X1    g0190(.A(G97), .ZN(new_n391));
  OAI22_X1  g0191(.A1(new_n390), .A2(new_n331), .B1(new_n319), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n392), .A2(KEYINPUT72), .A3(new_n278), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n287), .A2(G238), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n388), .A2(new_n296), .A3(new_n393), .A4(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT13), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n394), .A2(new_n296), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT13), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n397), .A2(new_n398), .A3(new_n388), .A4(new_n393), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n382), .B1(new_n400), .B2(G169), .ZN(new_n401));
  INV_X1    g0201(.A(G169), .ZN(new_n402));
  AOI211_X1 g0202(.A(KEYINPUT14), .B(new_n402), .C1(new_n396), .C2(new_n399), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n400), .A2(new_n299), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n381), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n400), .A2(G200), .ZN(new_n408));
  INV_X1    g0208(.A(new_n379), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n396), .A2(new_n399), .A3(G190), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT73), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT73), .A4(new_n410), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n407), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n272), .A2(G238), .A3(G1698), .ZN(new_n417));
  INV_X1    g0217(.A(G107), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n272), .A2(new_n274), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n417), .B1(new_n418), .B2(new_n272), .C1(new_n419), .C2(new_n214), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n278), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n287), .A2(G244), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(new_n296), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G200), .ZN(new_n424));
  INV_X1    g0224(.A(new_n251), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n258), .A2(new_n425), .B1(new_n253), .B2(new_n202), .ZN(new_n426));
  XOR2_X1   g0226(.A(KEYINPUT15), .B(G87), .Z(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(new_n254), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n261), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n264), .A2(G77), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n267), .A2(new_n202), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G190), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n424), .B(new_n434), .C1(new_n435), .C2(new_n423), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n423), .A2(new_n402), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n437), .B(new_n433), .C1(G179), .C2(new_n423), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n314), .A2(new_n370), .A3(new_n416), .A4(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT5), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT80), .B1(new_n441), .B2(G41), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT80), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(new_n280), .A3(KEYINPUT5), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n441), .A2(G41), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n281), .A2(G1), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n442), .A2(new_n444), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n283), .A2(G274), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n272), .A2(G257), .A3(new_n274), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n272), .A2(G264), .A3(G1698), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n331), .A2(G303), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n449), .B1(new_n453), .B2(new_n278), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n442), .A2(new_n444), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n293), .A2(G45), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(new_n441), .B2(G41), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n455), .A2(new_n457), .B1(new_n284), .B2(new_n286), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G270), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G200), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(new_n435), .B2(new_n460), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT20), .ZN(new_n463));
  INV_X1    g0263(.A(G116), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G20), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n261), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G283), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n253), .ZN(new_n468));
  XNOR2_X1  g0268(.A(KEYINPUT78), .B(G97), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(new_n319), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n463), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n468), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n391), .A2(KEYINPUT78), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT78), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G97), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n472), .B1(new_n476), .B2(G33), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n477), .A2(KEYINPUT20), .A3(new_n261), .A4(new_n465), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n268), .A2(G116), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n319), .A2(G1), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n261), .A2(new_n267), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n480), .B1(new_n482), .B2(G116), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT84), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT84), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n479), .A2(new_n486), .A3(new_n483), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n462), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n418), .A2(G20), .ZN(new_n490));
  XNOR2_X1  g0290(.A(new_n490), .B(KEYINPUT23), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n272), .A2(new_n253), .A3(G87), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT22), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT22), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n272), .A2(new_n494), .A3(new_n253), .A4(G87), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n254), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G116), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT24), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n496), .A2(KEYINPUT24), .A3(new_n498), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n261), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n482), .A2(G107), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n267), .A2(new_n418), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n505), .B(KEYINPUT25), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n503), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n289), .A2(G264), .A3(new_n447), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT85), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT85), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n289), .A2(new_n511), .A3(new_n447), .A4(G264), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n272), .A2(G257), .A3(G1698), .ZN(new_n514));
  INV_X1    g0314(.A(G294), .ZN(new_n515));
  OAI221_X1 g0315(.A(new_n514), .B1(new_n319), .B2(new_n515), .C1(new_n419), .C2(new_n209), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n278), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n518), .A2(new_n449), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n299), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n510), .A2(new_n512), .B1(new_n516), .B2(new_n278), .ZN(new_n521));
  OR2_X1    g0321(.A1(new_n447), .A2(new_n448), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n402), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n508), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT21), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n479), .A2(new_n486), .A3(new_n483), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n486), .B1(new_n479), .B2(new_n483), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n460), .A2(G169), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI211_X1 g0331(.A(new_n526), .B(new_n402), .C1(new_n454), .C2(new_n459), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n454), .A2(G179), .A3(new_n459), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  OAI22_X1  g0334(.A1(new_n532), .A2(new_n534), .B1(new_n527), .B2(new_n528), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n525), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT6), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(new_n473), .B2(new_n475), .ZN(new_n538));
  OAI21_X1  g0338(.A(G107), .B1(new_n391), .B2(KEYINPUT6), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n418), .A3(G97), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n542), .A2(G20), .B1(G77), .B2(new_n251), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT7), .B1(new_n331), .B2(new_n253), .ZN(new_n544));
  OAI21_X1  g0344(.A(G107), .B1(new_n318), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n262), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n268), .A2(G97), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n482), .B2(G97), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(KEYINPUT81), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n539), .B(new_n540), .C1(new_n469), .C2(new_n537), .ZN(new_n551));
  OAI22_X1  g0351(.A1(new_n551), .A2(new_n253), .B1(new_n202), .B2(new_n425), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n418), .B1(new_n330), .B2(new_n332), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n261), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT81), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n555), .A3(new_n548), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n320), .A2(new_n322), .A3(G244), .A4(new_n274), .ZN(new_n558));
  NOR2_X1   g0358(.A1(KEYINPUT79), .A2(KEYINPUT4), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n559), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n272), .A2(G244), .A3(new_n274), .A4(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n272), .A2(G250), .A3(G1698), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n560), .A2(new_n562), .A3(new_n467), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n278), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n449), .B1(new_n458), .B2(G257), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n565), .A2(new_n566), .A3(G179), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n402), .B1(new_n565), .B2(new_n566), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(KEYINPUT82), .B1(new_n557), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n565), .A2(new_n566), .A3(G179), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n289), .A2(G257), .A3(new_n447), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n522), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n278), .B2(new_n564), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n571), .B1(new_n574), .B2(new_n402), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT82), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n575), .A2(new_n576), .A3(new_n550), .A4(new_n556), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n570), .A2(new_n577), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n496), .A2(KEYINPUT24), .A3(new_n498), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT24), .B1(new_n496), .B2(new_n498), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n506), .B1(new_n581), .B2(new_n261), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n519), .A2(G190), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n523), .A2(G200), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n582), .A2(new_n504), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n482), .A2(new_n427), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n428), .A2(new_n267), .ZN(new_n587));
  NAND3_X1  g0387(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n588), .A2(new_n253), .ZN(new_n589));
  AOI21_X1  g0389(.A(G87), .B1(new_n473), .B2(new_n475), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n589), .B1(new_n590), .B2(new_n418), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n331), .A2(G20), .A3(new_n216), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT19), .B1(new_n469), .B2(new_n497), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n586), .B(new_n587), .C1(new_n594), .C2(new_n262), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n217), .A2(new_n274), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(G244), .B2(new_n274), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n597), .A2(new_n331), .B1(new_n319), .B2(new_n464), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n278), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n289), .A2(G250), .A3(new_n456), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n446), .A2(new_n283), .A3(G274), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n599), .A2(new_n299), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n601), .A3(new_n600), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n402), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n595), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(G200), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n272), .A2(new_n253), .A3(G68), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT19), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n476), .B2(new_n254), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n469), .A2(G87), .A3(G107), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n607), .B(new_n609), .C1(new_n610), .C2(new_n589), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n611), .A2(new_n261), .B1(new_n267), .B2(new_n428), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT83), .ZN(new_n613));
  INV_X1    g0413(.A(new_n481), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n262), .A2(new_n268), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n613), .B1(new_n615), .B2(new_n208), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n482), .A2(KEYINPUT83), .A3(G87), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n599), .A2(G190), .A3(new_n600), .A4(new_n601), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n606), .A2(new_n612), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n605), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n565), .A2(new_n566), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n622), .A2(new_n435), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(G200), .B2(new_n622), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n554), .A2(new_n548), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n578), .A2(new_n585), .A3(new_n621), .A4(new_n627), .ZN(new_n628));
  NOR4_X1   g0428(.A1(new_n440), .A2(new_n489), .A3(new_n536), .A4(new_n628), .ZN(G372));
  INV_X1    g0429(.A(new_n411), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n630), .A2(new_n438), .ZN(new_n631));
  OR3_X1    g0431(.A1(new_n407), .A2(new_n631), .A3(KEYINPUT87), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT87), .B1(new_n407), .B2(new_n631), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(new_n357), .A3(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n358), .A2(new_n359), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT18), .B1(new_n363), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT18), .ZN(new_n638));
  AOI221_X4 g0438(.A(new_n638), .B1(new_n358), .B2(new_n359), .C1(new_n336), .C2(new_n339), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n634), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n311), .A2(new_n313), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n302), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n440), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n575), .A2(new_n605), .A3(new_n620), .A4(new_n625), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n644), .A2(KEYINPUT26), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n605), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n570), .A2(new_n621), .A3(new_n577), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n647), .B1(new_n648), .B2(KEYINPUT26), .ZN(new_n649));
  INV_X1    g0449(.A(new_n530), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT21), .B1(new_n488), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n460), .A2(KEYINPUT21), .A3(G169), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n533), .A2(new_n652), .B1(new_n485), .B2(new_n487), .ZN(new_n653));
  OAI21_X1  g0453(.A(KEYINPUT86), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT86), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n530), .B1(new_n485), .B2(new_n487), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n535), .B(new_n655), .C1(new_n656), .C2(KEYINPUT21), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n654), .A2(new_n525), .A3(new_n657), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n646), .B(new_n649), .C1(new_n658), .C2(new_n628), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n643), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n642), .A2(new_n660), .ZN(G369));
  NOR2_X1   g0461(.A1(new_n266), .A2(G20), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n293), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G213), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n529), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n654), .A2(new_n657), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n489), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n531), .A2(new_n535), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n529), .B2(new_n669), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n671), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT88), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G330), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n508), .A2(new_n668), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n585), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n525), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n508), .A2(new_n524), .A3(new_n520), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n669), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n668), .B1(new_n531), .B2(new_n535), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT89), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(new_n682), .A3(new_n680), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n691), .A2(new_n682), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n685), .A2(new_n692), .ZN(G399));
  INV_X1    g0493(.A(new_n230), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G1), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n610), .A2(new_n464), .ZN(new_n698));
  OAI22_X1  g0498(.A1(new_n697), .A2(new_n698), .B1(new_n228), .B2(new_n696), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT28), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT91), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n654), .A2(new_n525), .A3(new_n657), .ZN(new_n702));
  AOI22_X1  g0502(.A1(new_n570), .A2(new_n577), .B1(new_n624), .B2(new_n626), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n702), .A2(new_n621), .A3(new_n703), .A4(new_n585), .ZN(new_n704));
  AOI211_X1 g0504(.A(new_n647), .B(new_n645), .C1(new_n648), .C2(KEYINPUT26), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n668), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(KEYINPUT29), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT26), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n570), .A2(new_n708), .A3(new_n621), .A4(new_n577), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n647), .B1(new_n644), .B2(KEYINPUT26), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n681), .A2(new_n673), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n709), .B(new_n710), .C1(new_n628), .C2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n669), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT90), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT90), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n712), .A2(new_n715), .A3(new_n669), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n707), .B1(new_n717), .B2(KEYINPUT29), .ZN(new_n718));
  NOR4_X1   g0518(.A1(new_n628), .A2(new_n536), .A3(new_n489), .A4(new_n668), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n574), .B1(new_n521), .B2(new_n522), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n720), .A2(new_n299), .A3(new_n460), .A4(new_n603), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  INV_X1    g0522(.A(new_n603), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n574), .A2(new_n521), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n722), .B1(new_n724), .B2(new_n533), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n518), .A2(new_n622), .A3(new_n603), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(KEYINPUT30), .A3(new_n534), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n721), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n668), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT31), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n728), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n719), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G330), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n701), .B1(new_n718), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n716), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n715), .B1(new_n712), .B2(new_n669), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT29), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n707), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n736), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n742), .A2(KEYINPUT91), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n737), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n700), .B1(new_n745), .B2(G1), .ZN(G364));
  INV_X1    g0546(.A(new_n677), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n662), .A2(G45), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n696), .A2(G1), .A3(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(G330), .B2(new_n676), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OR3_X1    g0554(.A1(new_n676), .A2(G20), .A3(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT94), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n253), .A2(new_n435), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G179), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n756), .B1(new_n758), .B2(G200), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n758), .A2(new_n756), .A3(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n272), .B1(new_n763), .B2(G322), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G179), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G190), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G311), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n253), .A2(G190), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(G179), .A3(new_n349), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n764), .B1(new_n515), .B2(new_n768), .C1(new_n769), .C2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n349), .A2(G179), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n772), .B1(G283), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n758), .A2(new_n349), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G326), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n770), .A2(new_n765), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT96), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G329), .ZN(new_n782));
  XNOR2_X1  g0582(.A(KEYINPUT97), .B(KEYINPUT33), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(G317), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n770), .A2(G179), .A3(G200), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n757), .A2(new_n773), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n784), .A2(new_n786), .B1(G303), .B2(new_n788), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n776), .A2(new_n778), .A3(new_n782), .A4(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n777), .ZN(new_n791));
  INV_X1    g0591(.A(G50), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n791), .A2(new_n792), .B1(new_n771), .B2(new_n202), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(new_n763), .B2(G58), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT95), .Z(new_n795));
  NAND2_X1  g0595(.A1(new_n788), .A2(G87), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n775), .A2(G107), .ZN(new_n797));
  INV_X1    g0597(.A(G159), .ZN(new_n798));
  OAI21_X1  g0598(.A(KEYINPUT32), .B1(new_n779), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n796), .A2(new_n797), .A3(new_n272), .A4(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n767), .A2(G97), .ZN(new_n802));
  INV_X1    g0602(.A(new_n779), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G159), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n801), .B(new_n802), .C1(KEYINPUT32), .C2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n785), .A2(new_n216), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n790), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n226), .B1(new_n253), .B2(G169), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n694), .A2(new_n331), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT92), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G355), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n324), .A2(new_n325), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n230), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT93), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n246), .B2(new_n281), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n228), .A2(G45), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n813), .B1(G116), .B2(new_n230), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n754), .A2(G20), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n809), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n755), .A2(new_n810), .A3(new_n823), .A4(new_n750), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n752), .A2(new_n824), .ZN(G396));
  NAND2_X1  g0625(.A1(new_n433), .A2(new_n668), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n436), .A2(new_n438), .A3(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT99), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n827), .B(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n438), .B2(new_n669), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n830), .A2(new_n754), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n802), .B1(new_n762), .B2(new_n515), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT98), .Z(new_n833));
  NAND2_X1  g0633(.A1(new_n781), .A2(G311), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G107), .A2(new_n788), .B1(new_n775), .B2(G87), .ZN(new_n835));
  INV_X1    g0635(.A(G303), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n791), .A2(new_n836), .B1(new_n771), .B2(new_n464), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n272), .B(new_n837), .C1(G283), .C2(new_n786), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n833), .A2(new_n834), .A3(new_n835), .A4(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n771), .A2(new_n798), .ZN(new_n840));
  INV_X1    g0640(.A(G137), .ZN(new_n841));
  INV_X1    g0641(.A(G150), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n791), .A2(new_n841), .B1(new_n785), .B2(new_n842), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n840), .B(new_n843), .C1(new_n763), .C2(G143), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT34), .Z(new_n845));
  NAND2_X1  g0645(.A1(new_n767), .A2(G58), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n775), .A2(G68), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n815), .B1(G50), .B2(new_n788), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(G132), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n780), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n839), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n809), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n809), .A2(new_n753), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n202), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n831), .A2(new_n750), .A3(new_n853), .A4(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n829), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n659), .A2(new_n669), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n706), .B2(new_n830), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n743), .B(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n856), .B1(new_n860), .B2(new_n750), .ZN(G384));
  OAI21_X1  g0661(.A(new_n316), .B1(new_n327), .B2(new_n216), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n329), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(new_n261), .A3(new_n328), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n635), .B1(new_n864), .B2(new_n339), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n336), .A2(new_n339), .A3(new_n351), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT102), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n331), .A2(KEYINPUT75), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n272), .A2(new_n323), .ZN(new_n869));
  AOI21_X1  g0669(.A(G20), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n332), .B1(new_n870), .B2(KEYINPUT7), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n334), .B1(new_n871), .B2(G68), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n262), .B1(new_n872), .B2(KEYINPUT16), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n338), .B1(new_n873), .B2(new_n863), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n666), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT102), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n878), .B(new_n352), .C1(new_n874), .C2(new_n635), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n867), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT37), .ZN(new_n881));
  XOR2_X1   g0681(.A(new_n666), .B(KEYINPUT103), .Z(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n363), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n367), .A2(new_n884), .A3(new_n885), .A4(new_n352), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n369), .A2(new_n876), .A3(new_n875), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(KEYINPUT38), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n635), .B1(new_n336), .B2(new_n339), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(new_n884), .A3(new_n352), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT37), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n354), .B(new_n355), .C1(new_n639), .C2(new_n637), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n882), .B1(new_n336), .B2(new_n339), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n886), .A2(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT104), .B1(new_n896), .B2(KEYINPUT38), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n639), .A2(new_n637), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n895), .B1(new_n898), .B2(new_n356), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n866), .A2(new_n890), .A3(new_n895), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n886), .B1(new_n900), .B2(new_n885), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT104), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT38), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n889), .A2(new_n897), .A3(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n407), .A2(new_n669), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n866), .A2(new_n895), .A3(KEYINPUT37), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n880), .A2(KEYINPUT37), .B1(new_n367), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n368), .A2(new_n366), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n877), .B1(new_n913), .B2(new_n357), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n904), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n889), .A2(new_n915), .A3(KEYINPUT39), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n908), .A2(new_n910), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n379), .B(KEYINPUT74), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n668), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n407), .B2(new_n415), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n401), .A2(new_n403), .A3(new_n405), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n919), .B(new_n411), .C1(new_n922), .C2(new_n381), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n889), .A2(new_n915), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT101), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n438), .A2(new_n668), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n926), .B(new_n927), .C1(new_n706), .C2(new_n857), .ZN(new_n928));
  INV_X1    g0728(.A(new_n927), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT101), .B1(new_n858), .B2(new_n929), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n924), .B(new_n925), .C1(new_n928), .C2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n898), .A2(new_n882), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n917), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n718), .A2(new_n643), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n642), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n933), .B(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n924), .B(new_n830), .C1(new_n719), .C2(new_n733), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n906), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT40), .B1(new_n889), .B2(new_n915), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n939), .A2(KEYINPUT40), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n734), .A2(new_n440), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT105), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n941), .B(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(G330), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n936), .B(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n293), .B2(new_n662), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT35), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n227), .B1(new_n551), .B2(new_n948), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n949), .B(G116), .C1(new_n948), .C2(new_n551), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT36), .ZN(new_n951));
  OAI21_X1  g0751(.A(G77), .B1(new_n213), .B2(new_n216), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n952), .A2(new_n228), .B1(G50), .B2(new_n216), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(G1), .A3(new_n266), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT100), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n947), .A2(new_n951), .A3(new_n955), .ZN(G367));
  OAI21_X1  g0756(.A(new_n703), .B1(new_n626), .B2(new_n669), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n575), .A2(new_n625), .A3(new_n668), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(KEYINPUT107), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n958), .A2(KEYINPUT107), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n957), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n685), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT108), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n691), .A2(new_n962), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT42), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n578), .B1(new_n962), .B2(new_n525), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n669), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n612), .A2(new_n618), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n668), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n621), .A2(new_n972), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n972), .A2(new_n605), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n976));
  NOR2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(KEYINPUT43), .B2(new_n975), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n970), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n967), .A2(new_n977), .A3(new_n969), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n963), .A2(new_n964), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n965), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n979), .A2(new_n964), .A3(new_n963), .A4(new_n980), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n695), .B(KEYINPUT41), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n692), .A2(new_n961), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT45), .Z(new_n990));
  NOR2_X1   g0790(.A1(new_n692), .A2(new_n961), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT44), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(new_n685), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n683), .A2(new_n689), .A3(new_n688), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n691), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n677), .B(new_n996), .ZN(new_n997));
  AOI211_X1 g0797(.A(KEYINPUT109), .B(new_n997), .C1(new_n737), .C2(new_n744), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT109), .ZN(new_n999));
  INV_X1    g0799(.A(new_n997), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n999), .B1(new_n745), .B2(new_n1000), .ZN(new_n1001));
  NOR3_X1   g0801(.A1(new_n998), .A2(new_n1001), .A3(KEYINPUT110), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT110), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n745), .A2(new_n1000), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(KEYINPUT109), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n745), .A2(new_n999), .A3(new_n1000), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1003), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n994), .B1(new_n1002), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n988), .B1(new_n1008), .B2(new_n745), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n748), .A2(G1), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n986), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n768), .A2(new_n216), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n763), .B2(G150), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT112), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n777), .A2(G143), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n774), .A2(new_n202), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G137), .B2(new_n803), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n792), .A2(new_n771), .B1(new_n785), .B2(new_n798), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n272), .B1(new_n213), .B2(new_n787), .C1(new_n1018), .C2(KEYINPUT113), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(KEYINPUT113), .B2(new_n1018), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .A4(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(G283), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n771), .A2(new_n1022), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n762), .A2(new_n836), .B1(new_n476), .B2(new_n774), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1023), .B(new_n1024), .C1(G294), .C2(new_n786), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n788), .A2(G116), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT46), .ZN(new_n1027));
  XOR2_X1   g0827(.A(KEYINPUT111), .B(G317), .Z(new_n1028));
  AOI22_X1  g0828(.A1(new_n777), .A2(G311), .B1(new_n803), .B2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1025), .A2(new_n815), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n768), .A2(new_n418), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1021), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT47), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n809), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n973), .A2(new_n821), .A3(new_n974), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n817), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n822), .B1(new_n230), .B2(new_n428), .C1(new_n1036), .C2(new_n241), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n750), .A3(new_n1035), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1011), .A2(new_n1038), .ZN(G387));
  AOI22_X1  g0839(.A1(new_n812), .A2(new_n698), .B1(new_n418), .B2(new_n694), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT114), .Z(new_n1041));
  OAI21_X1  g0841(.A(new_n817), .B1(new_n281), .B2(new_n238), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT50), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n258), .A2(G50), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n698), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1045), .B(new_n281), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(G68), .B2(G77), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1041), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n749), .B1(new_n1048), .B2(new_n822), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n763), .A2(new_n1028), .B1(G322), .B2(new_n777), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n836), .B2(new_n771), .C1(new_n769), .C2(new_n785), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT48), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n1022), .B2(new_n768), .C1(new_n515), .C2(new_n787), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT49), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n814), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n803), .A2(G326), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n1055), .C2(new_n1054), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G116), .B2(new_n775), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n777), .A2(G159), .B1(new_n427), .B2(new_n767), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n258), .B2(new_n785), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n774), .A2(new_n391), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n771), .A2(new_n216), .ZN(new_n1064));
  NOR4_X1   g0864(.A1(new_n1062), .A2(new_n815), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n788), .A2(G77), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n792), .B2(new_n762), .C1(new_n842), .C2(new_n779), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n808), .B1(new_n1060), .B2(new_n1068), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1050), .B(new_n1069), .C1(new_n683), .C2(new_n821), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n1000), .B2(new_n1010), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n695), .B1(new_n745), .B2(new_n1000), .C1(new_n998), .C2(new_n1001), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(G393));
  XNOR2_X1  g0873(.A(new_n993), .B(new_n684), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n998), .B2(new_n1001), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1008), .A2(new_n695), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n994), .A2(new_n1010), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n762), .A2(new_n798), .B1(new_n842), .B2(new_n791), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT51), .Z(new_n1079));
  NAND2_X1  g0879(.A1(new_n803), .A2(G143), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n767), .A2(G77), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1080), .B(new_n1081), .C1(new_n792), .C2(new_n785), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n787), .A2(new_n216), .B1(new_n774), .B2(new_n208), .ZN(new_n1083));
  OR4_X1    g0883(.A1(new_n815), .A2(new_n1079), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n771), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1084), .B1(new_n257), .B2(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n763), .A2(G311), .B1(G317), .B2(new_n777), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT52), .Z(new_n1088));
  AOI22_X1  g0888(.A1(new_n1085), .A2(G294), .B1(new_n767), .B2(G116), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n272), .B1(new_n803), .B2(G322), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1090), .B(new_n797), .C1(new_n1022), .C2(new_n787), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT116), .Z(new_n1092));
  NAND3_X1  g0892(.A1(new_n1088), .A2(new_n1089), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G303), .B2(new_n786), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n809), .B1(new_n1086), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n822), .B1(new_n230), .B2(new_n476), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n817), .B2(new_n249), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT115), .Z(new_n1098));
  NAND3_X1  g0898(.A1(new_n1095), .A2(new_n750), .A3(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1099), .A2(KEYINPUT117), .B1(new_n821), .B2(new_n962), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(KEYINPUT117), .B2(new_n1099), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1076), .A2(new_n1077), .A3(new_n1101), .ZN(G390));
  INV_X1    g0902(.A(new_n628), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1103), .A2(new_n672), .A3(new_n711), .A4(new_n669), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1104), .A2(new_n731), .A3(new_n732), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1105), .A2(G330), .A3(new_n830), .A4(new_n924), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n924), .B1(new_n928), .B2(new_n930), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1108), .A2(new_n909), .B1(new_n908), .B2(new_n916), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n906), .A2(new_n909), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n830), .B1(new_n738), .B2(new_n739), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n929), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1110), .B1(new_n1112), .B2(new_n924), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1107), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n908), .A2(new_n916), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n924), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n668), .B(new_n829), .C1(new_n704), .C2(new_n705), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n926), .B1(new_n1117), .B2(new_n927), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n858), .A2(KEYINPUT101), .A3(new_n929), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1116), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1115), .B1(new_n1120), .B2(new_n910), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n927), .B1(new_n717), .B2(new_n830), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n906), .B(new_n909), .C1(new_n1122), .C2(new_n1116), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(new_n1123), .A3(new_n1106), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n830), .B(G330), .C1(new_n719), .C2(new_n733), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n1116), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1106), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(KEYINPUT118), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1122), .A2(new_n1106), .A3(new_n1127), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT118), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1125), .A2(new_n1132), .A3(new_n1128), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1130), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n942), .A2(G330), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n934), .A2(new_n642), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1114), .A2(new_n1124), .A3(new_n1134), .A4(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n695), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT119), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n1109), .A2(new_n1113), .A3(new_n1107), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1106), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1138), .A2(KEYINPUT119), .A3(new_n695), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1141), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1144), .A2(new_n1010), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1115), .A2(new_n753), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n272), .B1(new_n788), .B2(G87), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(KEYINPUT120), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n777), .A2(G283), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1153), .A2(new_n847), .A3(new_n1081), .A4(new_n1154), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n763), .A2(G116), .B1(G107), .B2(new_n786), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1156), .B1(KEYINPUT120), .B2(new_n1152), .C1(new_n476), .C2(new_n771), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1155), .B(new_n1157), .C1(G294), .C2(new_n781), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n272), .B1(new_n785), .B2(new_n841), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G128), .B2(new_n777), .ZN(new_n1160));
  INV_X1    g0960(.A(G125), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1160), .B1(new_n1161), .B2(new_n780), .C1(new_n762), .C2(new_n850), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n787), .A2(new_n842), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT53), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT54), .B(G143), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1164), .B1(new_n798), .B2(new_n768), .C1(new_n771), .C2(new_n1165), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1162), .B(new_n1166), .C1(G50), .C2(new_n775), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n809), .B1(new_n1158), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n854), .A2(new_n258), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1151), .A2(new_n750), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1150), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1149), .A2(new_n1172), .ZN(G378));
  NAND3_X1  g0973(.A1(new_n917), .A2(new_n931), .A3(new_n932), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n271), .A2(new_n876), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n314), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n314), .A2(new_n1175), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1178), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n641), .A2(new_n301), .A3(new_n1175), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n314), .A2(new_n1175), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1179), .A2(new_n1183), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n889), .A2(new_n897), .A3(new_n905), .ZN(new_n1185));
  OAI21_X1  g0985(.A(KEYINPUT40), .B1(new_n1185), .B2(new_n937), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n940), .A2(new_n938), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n735), .B(new_n1184), .C1(new_n1186), .C2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1184), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n903), .B1(new_n902), .B2(new_n904), .ZN(new_n1190));
  AOI211_X1 g0990(.A(KEYINPUT104), .B(KEYINPUT38), .C1(new_n899), .C2(new_n901), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n937), .B1(new_n1192), .B2(new_n889), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT40), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1187), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1189), .B1(new_n1195), .B2(G330), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1174), .B1(new_n1188), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1184), .B1(new_n941), .B2(new_n735), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(G330), .A3(new_n1189), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1198), .A2(new_n933), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n1010), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1184), .A2(new_n753), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n786), .A2(G97), .B1(new_n1085), .B2(new_n427), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n1022), .B2(new_n780), .C1(new_n762), .C2(new_n418), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1012), .B(new_n1205), .C1(G58), .C2(new_n775), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n815), .A2(new_n280), .A3(new_n1066), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1206), .B(new_n1208), .C1(new_n464), .C2(new_n791), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT58), .Z(new_n1210));
  OAI22_X1  g1010(.A1(new_n841), .A2(new_n771), .B1(new_n787), .B2(new_n1165), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n791), .A2(new_n1161), .B1(new_n785), .B2(new_n850), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(G150), .C2(new_n767), .ZN(new_n1213));
  INV_X1    g1013(.A(G128), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1213), .B1(new_n1214), .B2(new_n762), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT59), .Z(new_n1216));
  AOI211_X1 g1016(.A(G33), .B(G41), .C1(new_n775), .C2(G159), .ZN(new_n1217));
  INV_X1    g1017(.A(G124), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1217), .B1(new_n1218), .B2(new_n779), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT121), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1216), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(G50), .B1(new_n319), .B2(new_n280), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n814), .B2(G41), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n809), .B1(new_n1210), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n854), .A2(new_n792), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1203), .A2(new_n750), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1202), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1138), .A2(new_n1137), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT57), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1231), .A2(new_n1233), .A3(KEYINPUT122), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT122), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1231), .A2(new_n1201), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n696), .B1(new_n1237), .B2(new_n1232), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1230), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(G375));
  NOR2_X1   g1040(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1241), .A2(new_n988), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n854), .A2(new_n216), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n924), .B2(new_n754), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n814), .B1(new_n785), .B2(new_n1165), .C1(new_n762), .C2(new_n841), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G50), .B2(new_n767), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n788), .A2(G159), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n781), .A2(G128), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n791), .A2(new_n850), .B1(new_n774), .B2(new_n213), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(G150), .B2(new_n1085), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .A4(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n787), .A2(new_n391), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n780), .A2(new_n836), .B1(new_n418), .B2(new_n771), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n1016), .B(new_n1255), .C1(G294), .C2(new_n777), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n763), .A2(G283), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n786), .A2(G116), .B1(new_n767), .B2(new_n427), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1256), .A2(new_n331), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1253), .B1(new_n1254), .B2(new_n1259), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n749), .B(new_n1246), .C1(new_n809), .C2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(new_n1134), .B2(new_n1010), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1244), .A2(new_n1262), .ZN(G381));
  OR2_X1    g1063(.A1(G393), .A2(G396), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1264), .A2(G384), .ZN(new_n1265));
  XOR2_X1   g1065(.A(new_n1265), .B(KEYINPUT123), .Z(new_n1266));
  INV_X1    g1066(.A(G381), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1076), .A2(new_n1077), .A3(new_n1101), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1268), .A2(new_n1011), .A3(new_n1038), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT124), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1138), .A2(KEYINPUT119), .A3(new_n695), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT119), .B1(new_n1138), .B2(new_n695), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1272), .A2(new_n1273), .A3(new_n1146), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1271), .B1(new_n1274), .B2(new_n1171), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1149), .A2(KEYINPUT124), .A3(new_n1172), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1277), .A2(new_n1239), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1266), .A2(new_n1267), .A3(new_n1270), .A4(new_n1278), .ZN(G407));
  INV_X1    g1079(.A(G213), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n1278), .B2(new_n667), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G407), .A2(new_n1281), .ZN(G409));
  INV_X1    g1082(.A(new_n1230), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1231), .A2(new_n987), .A3(new_n1201), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1277), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT125), .B1(new_n1239), .B2(G378), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1237), .A2(new_n1232), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT122), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1136), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1198), .A2(new_n933), .A3(new_n1199), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n933), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT57), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1289), .B1(new_n1290), .B2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1231), .A2(new_n1233), .A3(KEYINPUT122), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1288), .A2(new_n1294), .A3(new_n695), .A4(new_n1295), .ZN(new_n1296));
  AND4_X1   g1096(.A1(KEYINPUT125), .A2(new_n1296), .A3(G378), .A4(new_n1283), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1286), .B1(new_n1287), .B2(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1280), .A2(G343), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT60), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1243), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT126), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1241), .A2(KEYINPUT60), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1302), .A2(KEYINPUT126), .A3(new_n1243), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1305), .A2(new_n695), .A3(new_n1306), .A4(new_n1307), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1308), .A2(G384), .A3(new_n1262), .ZN(new_n1309));
  AOI21_X1  g1109(.A(G384), .B1(new_n1308), .B2(new_n1262), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1298), .A2(new_n1300), .A3(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(KEYINPUT62), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT61), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT127), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1299), .A2(G2897), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1315), .B(new_n1317), .C1(new_n1309), .C2(new_n1310), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1311), .A2(KEYINPUT127), .ZN(new_n1322));
  AOI22_X1  g1122(.A1(new_n1275), .A2(new_n1276), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1296), .A2(G378), .A3(new_n1283), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT125), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1296), .A2(G378), .A3(KEYINPUT125), .A4(new_n1283), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1323), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  OAI211_X1 g1128(.A(new_n1321), .B(new_n1322), .C1(new_n1328), .C2(new_n1299), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT62), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1298), .A2(new_n1330), .A3(new_n1300), .A4(new_n1311), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1313), .A2(new_n1314), .A3(new_n1329), .A4(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(KEYINPUT110), .B1(new_n998), .B2(new_n1001), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1005), .A2(new_n1006), .A3(new_n1003), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1074), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n745), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n987), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1010), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n985), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1038), .ZN(new_n1340));
  OAI21_X1  g1140(.A(G390), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  XNOR2_X1  g1141(.A(G393), .B(G396), .ZN(new_n1342));
  AND3_X1   g1142(.A1(new_n1269), .A2(new_n1341), .A3(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1342), .B1(new_n1269), .B2(new_n1341), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1332), .A2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1329), .A2(KEYINPUT63), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(new_n1312), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1298), .A2(KEYINPUT63), .A3(new_n1300), .A4(new_n1311), .ZN(new_n1350));
  AND3_X1   g1150(.A1(new_n1345), .A2(new_n1350), .A3(new_n1314), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1349), .A2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1347), .A2(new_n1352), .ZN(G405));
  AOI22_X1  g1153(.A1(new_n1326), .A2(new_n1327), .B1(G375), .B2(new_n1277), .ZN(new_n1354));
  OR3_X1    g1154(.A1(new_n1343), .A2(new_n1344), .A3(new_n1354), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1354), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1311), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1355), .A2(new_n1311), .A3(new_n1356), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1359), .A2(new_n1360), .ZN(G402));
endmodule


