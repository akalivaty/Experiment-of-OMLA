

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751;

  XOR2_X1 U367 ( .A(n475), .B(n474), .Z(n741) );
  INV_X2 U368 ( .A(G953), .ZN(n482) );
  NOR2_X2 U369 ( .A1(n556), .A2(n547), .ZN(n617) );
  AND2_X2 U370 ( .A1(n639), .A2(n429), .ZN(n408) );
  OR2_X2 U371 ( .A1(n642), .A2(G902), .ZN(n520) );
  XNOR2_X2 U372 ( .A(n603), .B(KEYINPUT1), .ZN(n677) );
  AND2_X1 U373 ( .A1(n398), .A2(n358), .ZN(n396) );
  NAND2_X1 U374 ( .A1(n396), .A2(n393), .ZN(n400) );
  NAND2_X1 U375 ( .A1(n395), .A2(n394), .ZN(n393) );
  NAND2_X1 U376 ( .A1(n374), .A2(n604), .ZN(n622) );
  XNOR2_X1 U377 ( .A(n375), .B(n602), .ZN(n374) );
  OR2_X1 U378 ( .A1(n605), .A2(n348), .ZN(n415) );
  XNOR2_X1 U379 ( .A(n491), .B(n490), .ZN(n670) );
  XNOR2_X1 U380 ( .A(n460), .B(n459), .ZN(n605) );
  XNOR2_X1 U381 ( .A(n486), .B(G134), .ZN(n508) );
  XNOR2_X1 U382 ( .A(KEYINPUT65), .B(KEYINPUT8), .ZN(n411) );
  XNOR2_X2 U383 ( .A(n740), .B(G146), .ZN(n519) );
  XNOR2_X2 U384 ( .A(n508), .B(n507), .ZN(n740) );
  XNOR2_X1 U385 ( .A(n615), .B(n386), .ZN(n385) );
  INV_X1 U386 ( .A(KEYINPUT73), .ZN(n386) );
  AND2_X1 U387 ( .A1(n611), .A2(n383), .ZN(n382) );
  AND2_X1 U388 ( .A1(n413), .A2(n587), .ZN(n491) );
  INV_X1 U389 ( .A(KEYINPUT72), .ZN(n383) );
  INV_X1 U390 ( .A(n352), .ZN(n416) );
  XNOR2_X1 U391 ( .A(KEYINPUT67), .B(KEYINPUT4), .ZN(n504) );
  XNOR2_X1 U392 ( .A(G101), .B(KEYINPUT69), .ZN(n442) );
  XNOR2_X1 U393 ( .A(n498), .B(n497), .ZN(n499) );
  INV_X1 U394 ( .A(G140), .ZN(n501) );
  INV_X1 U395 ( .A(KEYINPUT44), .ZN(n427) );
  NOR2_X1 U396 ( .A1(n382), .A2(n380), .ZN(n379) );
  XNOR2_X1 U397 ( .A(n454), .B(n453), .ZN(n549) );
  XNOR2_X1 U398 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U399 ( .A(n457), .B(n456), .ZN(n666) );
  INV_X1 U400 ( .A(KEYINPUT30), .ZN(n543) );
  XNOR2_X1 U401 ( .A(n440), .B(n439), .ZN(n733) );
  INV_X1 U402 ( .A(G110), .ZN(n439) );
  XNOR2_X1 U403 ( .A(G104), .B(G107), .ZN(n440) );
  XNOR2_X1 U404 ( .A(G119), .B(G110), .ZN(n522) );
  XNOR2_X1 U405 ( .A(G140), .B(KEYINPUT10), .ZN(n475) );
  AND2_X1 U406 ( .A1(n617), .A2(n667), .ZN(n618) );
  XNOR2_X1 U407 ( .A(n606), .B(KEYINPUT79), .ZN(n613) );
  NAND2_X1 U408 ( .A1(n373), .A2(n372), .ZN(n606) );
  INV_X1 U409 ( .A(n605), .ZN(n372) );
  INV_X1 U410 ( .A(n622), .ZN(n373) );
  OR2_X1 U411 ( .A1(n723), .A2(G902), .ZN(n371) );
  XNOR2_X1 U412 ( .A(n480), .B(n479), .ZN(n586) );
  XNOR2_X1 U413 ( .A(n412), .B(G478), .ZN(n587) );
  NOR2_X1 U414 ( .A1(n718), .A2(G902), .ZN(n412) );
  INV_X1 U415 ( .A(KEYINPUT85), .ZN(n361) );
  XNOR2_X1 U416 ( .A(G116), .B(G113), .ZN(n443) );
  INV_X1 U417 ( .A(KEYINPUT66), .ZN(n468) );
  NOR2_X1 U418 ( .A1(n610), .A2(n383), .ZN(n378) );
  AND2_X1 U419 ( .A1(n381), .A2(n383), .ZN(n380) );
  NAND2_X1 U420 ( .A1(n482), .A2(G234), .ZN(n410) );
  XOR2_X1 U421 ( .A(G104), .B(G122), .Z(n471) );
  XNOR2_X1 U422 ( .A(G113), .B(G143), .ZN(n470) );
  XOR2_X1 U423 ( .A(KEYINPUT87), .B(KEYINPUT17), .Z(n433) );
  AND2_X1 U424 ( .A1(n419), .A2(n345), .ZN(n365) );
  INV_X1 U425 ( .A(KEYINPUT0), .ZN(n418) );
  XNOR2_X1 U426 ( .A(KEYINPUT16), .B(G122), .ZN(n447) );
  XNOR2_X1 U427 ( .A(n503), .B(n502), .ZN(n509) );
  XNOR2_X1 U428 ( .A(n501), .B(G101), .ZN(n502) );
  XNOR2_X1 U429 ( .A(KEYINPUT83), .B(KEYINPUT45), .ZN(n598) );
  NOR2_X1 U430 ( .A1(n409), .A2(n670), .ZN(n621) );
  BUF_X1 U431 ( .A(n549), .Z(n627) );
  XNOR2_X1 U432 ( .A(n544), .B(n543), .ZN(n545) );
  INV_X1 U433 ( .A(KEYINPUT102), .ZN(n392) );
  INV_X1 U434 ( .A(n643), .ZN(n394) );
  OR2_X1 U435 ( .A1(n643), .A2(G472), .ZN(n397) );
  XNOR2_X1 U436 ( .A(G128), .B(G137), .ZN(n521) );
  AND2_X1 U437 ( .A1(n640), .A2(G210), .ZN(n402) );
  NAND2_X1 U438 ( .A1(n406), .A2(n405), .ZN(n639) );
  INV_X1 U439 ( .A(n637), .ZN(n405) );
  AND2_X1 U440 ( .A1(n728), .A2(n600), .ZN(n406) );
  NOR2_X1 U441 ( .A1(n607), .A2(n655), .ZN(n646) );
  XNOR2_X1 U442 ( .A(n388), .B(n387), .ZN(G60) );
  INV_X1 U443 ( .A(KEYINPUT60), .ZN(n387) );
  NAND2_X1 U444 ( .A1(n389), .A2(n644), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n390), .B(n359), .ZN(n389) );
  XNOR2_X1 U446 ( .A(n368), .B(n367), .ZN(G51) );
  INV_X1 U447 ( .A(KEYINPUT56), .ZN(n367) );
  NAND2_X1 U448 ( .A1(n369), .A2(n644), .ZN(n368) );
  XNOR2_X1 U449 ( .A(n370), .B(n346), .ZN(n369) );
  XNOR2_X1 U450 ( .A(n401), .B(n357), .ZN(n571) );
  AND2_X1 U451 ( .A1(n415), .A2(n419), .ZN(n343) );
  NOR2_X1 U452 ( .A1(n681), .A2(n416), .ZN(n344) );
  AND2_X1 U453 ( .A1(n344), .A2(KEYINPUT22), .ZN(n345) );
  XOR2_X1 U454 ( .A(n708), .B(n710), .Z(n346) );
  XOR2_X1 U455 ( .A(n532), .B(n531), .Z(n347) );
  OR2_X1 U456 ( .A1(n417), .A2(KEYINPUT0), .ZN(n348) );
  AND2_X1 U457 ( .A1(n422), .A2(n361), .ZN(n349) );
  INV_X1 U458 ( .A(n610), .ZN(n384) );
  AND2_X1 U459 ( .A1(n366), .A2(n344), .ZN(n350) );
  AND2_X1 U460 ( .A1(n365), .A2(n415), .ZN(n351) );
  OR2_X1 U461 ( .A1(n431), .A2(n418), .ZN(n352) );
  AND2_X1 U462 ( .A1(n677), .A2(n555), .ZN(n353) );
  NOR2_X1 U463 ( .A1(n409), .A2(n671), .ZN(n354) );
  AND2_X1 U464 ( .A1(n553), .A2(n559), .ZN(n355) );
  AND2_X1 U465 ( .A1(n419), .A2(n352), .ZN(n356) );
  XOR2_X1 U466 ( .A(KEYINPUT64), .B(KEYINPUT32), .Z(n357) );
  AND2_X1 U467 ( .A1(n397), .A2(n644), .ZN(n358) );
  XNOR2_X1 U468 ( .A(n717), .B(KEYINPUT59), .ZN(n359) );
  NOR2_X1 U469 ( .A1(n482), .A2(G952), .ZN(n725) );
  INV_X1 U470 ( .A(KEYINPUT84), .ZN(n600) );
  XOR2_X1 U471 ( .A(G110), .B(KEYINPUT111), .Z(n360) );
  XNOR2_X1 U472 ( .A(n422), .B(n360), .ZN(G12) );
  NAND2_X1 U473 ( .A1(n391), .A2(n355), .ZN(n422) );
  NAND2_X1 U474 ( .A1(n364), .A2(n362), .ZN(n554) );
  NAND2_X1 U475 ( .A1(n363), .A2(n496), .ZN(n362) );
  NAND2_X1 U476 ( .A1(n350), .A2(n343), .ZN(n363) );
  NAND2_X1 U477 ( .A1(n351), .A2(n366), .ZN(n364) );
  INV_X1 U478 ( .A(n670), .ZN(n366) );
  NAND2_X1 U479 ( .A1(n402), .A2(n408), .ZN(n370) );
  NAND2_X1 U480 ( .A1(n559), .A2(n558), .ZN(n561) );
  XNOR2_X2 U481 ( .A(n371), .B(n347), .ZN(n559) );
  XNOR2_X1 U482 ( .A(n527), .B(n528), .ZN(n723) );
  NAND2_X1 U483 ( .A1(n601), .A2(n685), .ZN(n375) );
  NAND2_X1 U484 ( .A1(n379), .A2(n376), .ZN(n631) );
  OR2_X1 U485 ( .A1(n611), .A2(n377), .ZN(n376) );
  NAND2_X1 U486 ( .A1(n385), .A2(n378), .ZN(n377) );
  NAND2_X1 U487 ( .A1(n385), .A2(n384), .ZN(n381) );
  NAND2_X1 U488 ( .A1(n554), .A2(n565), .ZN(n552) );
  NAND2_X1 U489 ( .A1(n403), .A2(n408), .ZN(n390) );
  XNOR2_X1 U490 ( .A(n552), .B(n392), .ZN(n391) );
  XNOR2_X1 U491 ( .A(n425), .B(n427), .ZN(n597) );
  NAND2_X1 U492 ( .A1(n549), .A2(n666), .ZN(n460) );
  INV_X1 U493 ( .A(n721), .ZN(n395) );
  NAND2_X1 U494 ( .A1(n721), .A2(n399), .ZN(n398) );
  AND2_X1 U495 ( .A1(n643), .A2(G472), .ZN(n399) );
  XNOR2_X1 U496 ( .A(n400), .B(n645), .ZN(G57) );
  INV_X1 U497 ( .A(n571), .ZN(n421) );
  NAND2_X1 U498 ( .A1(n554), .A2(n353), .ZN(n401) );
  AND2_X2 U499 ( .A1(n408), .A2(n640), .ZN(n721) );
  AND2_X1 U500 ( .A1(n640), .A2(G475), .ZN(n403) );
  NAND2_X1 U501 ( .A1(n404), .A2(n637), .ZN(n407) );
  NOR2_X1 U502 ( .A1(n638), .A2(n600), .ZN(n404) );
  XNOR2_X2 U503 ( .A(n407), .B(KEYINPUT2), .ZN(n640) );
  NAND2_X1 U504 ( .A1(n605), .A2(KEYINPUT0), .ZN(n419) );
  NAND2_X1 U505 ( .A1(n667), .A2(n666), .ZN(n409) );
  XNOR2_X2 U506 ( .A(n411), .B(n410), .ZN(n483) );
  INV_X1 U507 ( .A(n587), .ZN(n548) );
  INV_X1 U508 ( .A(n586), .ZN(n413) );
  NOR2_X2 U509 ( .A1(n749), .A2(n751), .ZN(n624) );
  NOR2_X2 U510 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X2 U511 ( .A(n414), .B(G143), .ZN(n486) );
  XNOR2_X2 U512 ( .A(G128), .B(KEYINPUT80), .ZN(n414) );
  NAND2_X1 U513 ( .A1(n356), .A2(n415), .ZN(n582) );
  INV_X1 U514 ( .A(n431), .ZN(n417) );
  NAND2_X1 U515 ( .A1(n349), .A2(n421), .ZN(n423) );
  NAND2_X1 U516 ( .A1(n420), .A2(KEYINPUT85), .ZN(n424) );
  NAND2_X1 U517 ( .A1(n422), .A2(n421), .ZN(n420) );
  NAND2_X1 U518 ( .A1(n424), .A2(n423), .ZN(n426) );
  NAND2_X1 U519 ( .A1(n426), .A2(n428), .ZN(n425) );
  INV_X1 U520 ( .A(n750), .ZN(n428) );
  NAND2_X1 U521 ( .A1(n640), .A2(n639), .ZN(n430) );
  INV_X1 U522 ( .A(n641), .ZN(n429) );
  AND2_X1 U523 ( .A1(n706), .A2(n430), .ZN(n707) );
  XNOR2_X1 U524 ( .A(n485), .B(n484), .ZN(n487) );
  XNOR2_X1 U525 ( .A(n508), .B(n487), .ZN(n488) );
  AND2_X1 U526 ( .A1(n467), .A2(n466), .ZN(n431) );
  AND2_X1 U527 ( .A1(n630), .A2(n663), .ZN(n432) );
  INV_X1 U528 ( .A(KEYINPUT92), .ZN(n497) );
  XNOR2_X1 U529 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n505), .B(n469), .ZN(n473) );
  XNOR2_X1 U531 ( .A(n530), .B(KEYINPUT77), .ZN(n531) );
  XNOR2_X1 U532 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U533 ( .A(n526), .B(n741), .ZN(n527) );
  XOR2_X1 U534 ( .A(G101), .B(KEYINPUT109), .Z(n536) );
  XNOR2_X1 U535 ( .A(n486), .B(n433), .ZN(n438) );
  NAND2_X1 U536 ( .A1(G224), .A2(n482), .ZN(n435) );
  XNOR2_X1 U537 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n434) );
  XNOR2_X1 U538 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X2 U539 ( .A(G146), .B(G125), .Z(n474) );
  XNOR2_X1 U540 ( .A(n436), .B(n474), .ZN(n437) );
  XNOR2_X1 U541 ( .A(n438), .B(n437), .ZN(n441) );
  XNOR2_X1 U542 ( .A(n733), .B(KEYINPUT70), .ZN(n500) );
  XNOR2_X1 U543 ( .A(n441), .B(n500), .ZN(n449) );
  XNOR2_X1 U544 ( .A(n443), .B(n442), .ZN(n445) );
  XNOR2_X1 U545 ( .A(KEYINPUT3), .B(G119), .ZN(n444) );
  XNOR2_X1 U546 ( .A(n445), .B(n444), .ZN(n517) );
  INV_X1 U547 ( .A(KEYINPUT71), .ZN(n446) );
  XNOR2_X1 U548 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U549 ( .A(n517), .B(n448), .ZN(n732) );
  XNOR2_X1 U550 ( .A(n449), .B(n732), .ZN(n708) );
  XNOR2_X1 U551 ( .A(KEYINPUT15), .B(G902), .ZN(n641) );
  NAND2_X1 U552 ( .A1(n708), .A2(n641), .ZN(n454) );
  NOR2_X1 U553 ( .A1(G902), .A2(G237), .ZN(n450) );
  XNOR2_X1 U554 ( .A(n450), .B(KEYINPUT75), .ZN(n455) );
  NAND2_X1 U555 ( .A1(n455), .A2(G210), .ZN(n452) );
  INV_X1 U556 ( .A(KEYINPUT88), .ZN(n451) );
  NAND2_X1 U557 ( .A1(n455), .A2(G214), .ZN(n457) );
  INV_X1 U558 ( .A(KEYINPUT89), .ZN(n456) );
  INV_X1 U559 ( .A(KEYINPUT76), .ZN(n458) );
  XNOR2_X1 U560 ( .A(n458), .B(KEYINPUT19), .ZN(n459) );
  XOR2_X1 U561 ( .A(KEYINPUT90), .B(KEYINPUT14), .Z(n463) );
  NAND2_X1 U562 ( .A1(G234), .A2(G237), .ZN(n461) );
  XNOR2_X1 U563 ( .A(n461), .B(KEYINPUT74), .ZN(n462) );
  XNOR2_X1 U564 ( .A(n463), .B(n462), .ZN(n700) );
  INV_X1 U565 ( .A(n700), .ZN(n467) );
  XNOR2_X1 U566 ( .A(G898), .B(KEYINPUT91), .ZN(n734) );
  NAND2_X1 U567 ( .A1(G953), .A2(G902), .ZN(n537) );
  INV_X1 U568 ( .A(n537), .ZN(n464) );
  NAND2_X1 U569 ( .A1(n734), .A2(n464), .ZN(n465) );
  NAND2_X1 U570 ( .A1(n482), .A2(G952), .ZN(n540) );
  NAND2_X1 U571 ( .A1(n465), .A2(n540), .ZN(n466) );
  XNOR2_X1 U572 ( .A(KEYINPUT13), .B(G475), .ZN(n480) );
  XNOR2_X1 U573 ( .A(n468), .B(G131), .ZN(n505) );
  XNOR2_X1 U574 ( .A(n471), .B(n470), .ZN(n472) );
  XOR2_X1 U575 ( .A(n473), .B(n472), .Z(n478) );
  NOR2_X1 U576 ( .A1(G953), .A2(G237), .ZN(n512) );
  NAND2_X1 U577 ( .A1(G214), .A2(n512), .ZN(n476) );
  XNOR2_X1 U578 ( .A(n741), .B(n476), .ZN(n477) );
  XNOR2_X1 U579 ( .A(n478), .B(n477), .ZN(n717) );
  NOR2_X1 U580 ( .A1(G902), .A2(n717), .ZN(n479) );
  XNOR2_X1 U581 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n489) );
  XOR2_X1 U582 ( .A(G107), .B(G122), .Z(n481) );
  XOR2_X1 U583 ( .A(n481), .B(G116), .Z(n485) );
  NAND2_X1 U584 ( .A1(n483), .A2(G217), .ZN(n484) );
  XNOR2_X1 U585 ( .A(n489), .B(n488), .ZN(n718) );
  INV_X1 U586 ( .A(KEYINPUT100), .ZN(n490) );
  NAND2_X1 U587 ( .A1(G234), .A2(n641), .ZN(n492) );
  XNOR2_X1 U588 ( .A(KEYINPUT20), .B(n492), .ZN(n529) );
  NAND2_X1 U589 ( .A1(n529), .A2(G221), .ZN(n494) );
  XOR2_X1 U590 ( .A(KEYINPUT95), .B(KEYINPUT21), .Z(n493) );
  XNOR2_X1 U591 ( .A(n494), .B(n493), .ZN(n681) );
  INV_X1 U592 ( .A(n681), .ZN(n495) );
  INV_X1 U593 ( .A(KEYINPUT22), .ZN(n496) );
  NAND2_X1 U594 ( .A1(G227), .A2(n482), .ZN(n498) );
  XNOR2_X1 U595 ( .A(n500), .B(n499), .ZN(n503) );
  XNOR2_X1 U596 ( .A(n504), .B(G137), .ZN(n506) );
  XNOR2_X1 U597 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U598 ( .A(n519), .B(n509), .ZN(n711) );
  NOR2_X1 U599 ( .A1(n711), .A2(G902), .ZN(n511) );
  INV_X1 U600 ( .A(G469), .ZN(n510) );
  XNOR2_X2 U601 ( .A(n511), .B(n510), .ZN(n603) );
  INV_X1 U602 ( .A(n677), .ZN(n565) );
  NAND2_X1 U603 ( .A1(n512), .A2(G210), .ZN(n513) );
  XNOR2_X1 U604 ( .A(n513), .B(KEYINPUT5), .ZN(n515) );
  XNOR2_X1 U605 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n514) );
  XNOR2_X1 U606 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U607 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U608 ( .A(n519), .B(n518), .ZN(n642) );
  XNOR2_X2 U609 ( .A(n520), .B(G472), .ZN(n685) );
  XNOR2_X1 U610 ( .A(n685), .B(KEYINPUT6), .ZN(n572) );
  XNOR2_X1 U611 ( .A(n521), .B(KEYINPUT23), .ZN(n528) );
  NAND2_X1 U612 ( .A1(n483), .A2(G221), .ZN(n525) );
  XOR2_X1 U613 ( .A(KEYINPUT93), .B(KEYINPUT24), .Z(n523) );
  XNOR2_X1 U614 ( .A(n523), .B(n522), .ZN(n524) );
  NAND2_X1 U615 ( .A1(n529), .A2(G217), .ZN(n532) );
  XNOR2_X1 U616 ( .A(KEYINPUT25), .B(KEYINPUT94), .ZN(n530) );
  INV_X1 U617 ( .A(KEYINPUT101), .ZN(n533) );
  XNOR2_X1 U618 ( .A(n559), .B(n533), .ZN(n682) );
  INV_X1 U619 ( .A(n682), .ZN(n534) );
  NAND2_X1 U620 ( .A1(n572), .A2(n534), .ZN(n535) );
  NOR2_X1 U621 ( .A1(n552), .A2(n535), .ZN(n594) );
  XOR2_X1 U622 ( .A(n536), .B(n594), .Z(G3) );
  XNOR2_X1 U623 ( .A(G143), .B(KEYINPUT112), .ZN(n551) );
  NOR2_X1 U624 ( .A1(n700), .A2(n537), .ZN(n538) );
  XNOR2_X1 U625 ( .A(n538), .B(KEYINPUT103), .ZN(n539) );
  NOR2_X1 U626 ( .A1(G900), .A2(n539), .ZN(n542) );
  NOR2_X1 U627 ( .A1(n700), .A2(n540), .ZN(n541) );
  NOR2_X1 U628 ( .A1(n542), .A2(n541), .ZN(n556) );
  NOR2_X1 U629 ( .A1(n681), .A2(n559), .ZN(n678) );
  NAND2_X1 U630 ( .A1(n603), .A2(n678), .ZN(n583) );
  XNOR2_X1 U631 ( .A(n583), .B(KEYINPUT105), .ZN(n546) );
  NAND2_X1 U632 ( .A1(n685), .A2(n666), .ZN(n544) );
  NAND2_X1 U633 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U634 ( .A1(n586), .A2(n548), .ZN(n575) );
  INV_X1 U635 ( .A(n627), .ZN(n568) );
  NOR2_X1 U636 ( .A1(n575), .A2(n568), .ZN(n550) );
  AND2_X1 U637 ( .A1(n617), .A2(n550), .ZN(n610) );
  XOR2_X1 U638 ( .A(n551), .B(n610), .Z(G45) );
  INV_X1 U639 ( .A(n685), .ZN(n553) );
  AND2_X1 U640 ( .A1(n572), .A2(n682), .ZN(n555) );
  XOR2_X1 U641 ( .A(G119), .B(n571), .Z(G21) );
  NAND2_X1 U642 ( .A1(n587), .A2(n586), .ZN(n655) );
  INV_X1 U643 ( .A(n572), .ZN(n562) );
  INV_X1 U644 ( .A(n556), .ZN(n557) );
  AND2_X1 U645 ( .A1(n557), .A2(n495), .ZN(n558) );
  INV_X1 U646 ( .A(KEYINPUT68), .ZN(n560) );
  XNOR2_X1 U647 ( .A(n561), .B(n560), .ZN(n601) );
  NAND2_X1 U648 ( .A1(n562), .A2(n601), .ZN(n563) );
  NOR2_X1 U649 ( .A1(n655), .A2(n563), .ZN(n564) );
  NAND2_X1 U650 ( .A1(n666), .A2(n564), .ZN(n625) );
  XOR2_X1 U651 ( .A(n625), .B(KEYINPUT104), .Z(n566) );
  NAND2_X1 U652 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U653 ( .A(n567), .B(KEYINPUT43), .ZN(n569) );
  NAND2_X1 U654 ( .A1(n569), .A2(n568), .ZN(n634) );
  XOR2_X1 U655 ( .A(G140), .B(KEYINPUT115), .Z(n570) );
  XNOR2_X1 U656 ( .A(n634), .B(n570), .ZN(G42) );
  NAND2_X1 U657 ( .A1(n677), .A2(n678), .ZN(n579) );
  NOR2_X1 U658 ( .A1(n579), .A2(n572), .ZN(n573) );
  XNOR2_X1 U659 ( .A(n573), .B(KEYINPUT33), .ZN(n676) );
  NOR2_X1 U660 ( .A1(n676), .A2(n582), .ZN(n574) );
  XNOR2_X1 U661 ( .A(n574), .B(KEYINPUT34), .ZN(n577) );
  XOR2_X1 U662 ( .A(n575), .B(KEYINPUT78), .Z(n576) );
  NAND2_X1 U663 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U664 ( .A(n578), .B(KEYINPUT35), .ZN(n750) );
  INV_X1 U665 ( .A(n579), .ZN(n580) );
  NAND2_X1 U666 ( .A1(n580), .A2(n685), .ZN(n690) );
  NOR2_X1 U667 ( .A1(n690), .A2(n582), .ZN(n581) );
  XNOR2_X1 U668 ( .A(n581), .B(KEYINPUT31), .ZN(n658) );
  INV_X1 U669 ( .A(n582), .ZN(n585) );
  NOR2_X1 U670 ( .A1(n583), .A2(n685), .ZN(n584) );
  NAND2_X1 U671 ( .A1(n585), .A2(n584), .ZN(n652) );
  NAND2_X1 U672 ( .A1(n658), .A2(n652), .ZN(n592) );
  NOR2_X1 U673 ( .A1(n587), .A2(n586), .ZN(n589) );
  INV_X1 U674 ( .A(KEYINPUT98), .ZN(n588) );
  XNOR2_X1 U675 ( .A(n589), .B(n588), .ZN(n659) );
  INV_X1 U676 ( .A(n659), .ZN(n608) );
  INV_X1 U677 ( .A(n655), .ZN(n590) );
  NOR2_X1 U678 ( .A1(n608), .A2(n590), .ZN(n671) );
  XNOR2_X1 U679 ( .A(n671), .B(KEYINPUT82), .ZN(n612) );
  INV_X1 U680 ( .A(n612), .ZN(n591) );
  NAND2_X1 U681 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U682 ( .A(n593), .B(KEYINPUT99), .ZN(n595) );
  NOR2_X1 U683 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U684 ( .A1(n597), .A2(n596), .ZN(n599) );
  XNOR2_X1 U685 ( .A(n599), .B(n598), .ZN(n638) );
  XNOR2_X1 U686 ( .A(KEYINPUT107), .B(KEYINPUT28), .ZN(n602) );
  XNOR2_X1 U687 ( .A(n603), .B(KEYINPUT106), .ZN(n604) );
  INV_X1 U688 ( .A(n613), .ZN(n607) );
  NAND2_X1 U689 ( .A1(n613), .A2(n608), .ZN(n648) );
  NAND2_X1 U690 ( .A1(n648), .A2(KEYINPUT47), .ZN(n609) );
  NOR2_X1 U691 ( .A1(n646), .A2(n609), .ZN(n611) );
  NOR2_X1 U692 ( .A1(n612), .A2(KEYINPUT47), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n614), .A2(n613), .ZN(n615) );
  INV_X1 U694 ( .A(KEYINPUT38), .ZN(n616) );
  XNOR2_X1 U695 ( .A(n627), .B(n616), .ZN(n667) );
  XNOR2_X1 U696 ( .A(n618), .B(KEYINPUT39), .ZN(n633) );
  NOR2_X1 U697 ( .A1(n655), .A2(n633), .ZN(n620) );
  XNOR2_X1 U698 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n619) );
  XNOR2_X1 U699 ( .A(n620), .B(n619), .ZN(n749) );
  XNOR2_X1 U700 ( .A(KEYINPUT41), .B(n621), .ZN(n694) );
  NOR2_X1 U701 ( .A1(n694), .A2(n622), .ZN(n623) );
  XNOR2_X1 U702 ( .A(n623), .B(KEYINPUT42), .ZN(n751) );
  XNOR2_X1 U703 ( .A(n624), .B(KEYINPUT46), .ZN(n630) );
  INV_X1 U704 ( .A(n625), .ZN(n626) );
  AND2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U706 ( .A(n628), .B(KEYINPUT36), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n677), .A2(n629), .ZN(n663) );
  NAND2_X1 U708 ( .A1(n631), .A2(n432), .ZN(n632) );
  XNOR2_X1 U709 ( .A(n632), .B(KEYINPUT48), .ZN(n636) );
  OR2_X1 U710 ( .A1(n633), .A2(n659), .ZN(n664) );
  NAND2_X1 U711 ( .A1(n634), .A2(n664), .ZN(n635) );
  INV_X1 U712 ( .A(n638), .ZN(n728) );
  XOR2_X1 U713 ( .A(KEYINPUT62), .B(n642), .Z(n643) );
  INV_X1 U714 ( .A(n725), .ZN(n644) );
  XNOR2_X1 U715 ( .A(KEYINPUT86), .B(KEYINPUT63), .ZN(n645) );
  XOR2_X1 U716 ( .A(n646), .B(G146), .Z(G48) );
  XOR2_X1 U717 ( .A(G128), .B(KEYINPUT29), .Z(n647) );
  XNOR2_X1 U718 ( .A(n648), .B(n647), .ZN(G30) );
  NOR2_X1 U719 ( .A1(n652), .A2(n655), .ZN(n649) );
  XOR2_X1 U720 ( .A(G104), .B(n649), .Z(G6) );
  XOR2_X1 U721 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n651) );
  XNOR2_X1 U722 ( .A(G107), .B(KEYINPUT110), .ZN(n650) );
  XNOR2_X1 U723 ( .A(n651), .B(n650), .ZN(n654) );
  NOR2_X1 U724 ( .A1(n652), .A2(n659), .ZN(n653) );
  XOR2_X1 U725 ( .A(n654), .B(n653), .Z(G9) );
  NOR2_X1 U726 ( .A1(n655), .A2(n658), .ZN(n657) );
  XNOR2_X1 U727 ( .A(G113), .B(KEYINPUT113), .ZN(n656) );
  XNOR2_X1 U728 ( .A(n657), .B(n656), .ZN(G15) );
  NOR2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U730 ( .A(KEYINPUT114), .B(n660), .Z(n661) );
  XNOR2_X1 U731 ( .A(G116), .B(n661), .ZN(G18) );
  XOR2_X1 U732 ( .A(G125), .B(KEYINPUT37), .Z(n662) );
  XNOR2_X1 U733 ( .A(n663), .B(n662), .ZN(G27) );
  INV_X1 U734 ( .A(n664), .ZN(n665) );
  XOR2_X1 U735 ( .A(G134), .B(n665), .Z(G36) );
  NOR2_X1 U736 ( .A1(n694), .A2(n676), .ZN(n703) );
  NOR2_X1 U737 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U738 ( .A(KEYINPUT119), .B(n668), .Z(n669) );
  NOR2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n673) );
  XNOR2_X1 U740 ( .A(n354), .B(KEYINPUT120), .ZN(n672) );
  NOR2_X1 U741 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U742 ( .A(KEYINPUT121), .B(n674), .Z(n675) );
  NOR2_X1 U743 ( .A1(n676), .A2(n675), .ZN(n696) );
  OR2_X1 U744 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U745 ( .A(n679), .B(KEYINPUT118), .ZN(n680) );
  XNOR2_X1 U746 ( .A(KEYINPUT50), .B(n680), .ZN(n689) );
  NAND2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U748 ( .A(n683), .B(KEYINPUT49), .ZN(n684) );
  XNOR2_X1 U749 ( .A(n684), .B(KEYINPUT116), .ZN(n686) );
  NOR2_X1 U750 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U751 ( .A(KEYINPUT117), .B(n687), .Z(n688) );
  NAND2_X1 U752 ( .A1(n689), .A2(n688), .ZN(n691) );
  NAND2_X1 U753 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U754 ( .A(KEYINPUT51), .B(n692), .ZN(n693) );
  NOR2_X1 U755 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U756 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U757 ( .A(n697), .B(KEYINPUT122), .Z(n698) );
  XNOR2_X1 U758 ( .A(KEYINPUT52), .B(n698), .ZN(n699) );
  NAND2_X1 U759 ( .A1(G952), .A2(n699), .ZN(n701) );
  NOR2_X1 U760 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U761 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U762 ( .A(n704), .B(KEYINPUT123), .ZN(n705) );
  NOR2_X1 U763 ( .A1(n705), .A2(G953), .ZN(n706) );
  XNOR2_X1 U764 ( .A(KEYINPUT53), .B(n707), .ZN(G75) );
  XOR2_X1 U765 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n709) );
  XNOR2_X1 U766 ( .A(n709), .B(KEYINPUT81), .ZN(n710) );
  NAND2_X1 U767 ( .A1(n721), .A2(G469), .ZN(n715) );
  XOR2_X1 U768 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n713) );
  XNOR2_X1 U769 ( .A(n711), .B(KEYINPUT124), .ZN(n712) );
  XNOR2_X1 U770 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X1 U771 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U772 ( .A1(n725), .A2(n716), .ZN(G54) );
  NAND2_X1 U773 ( .A1(n721), .A2(G478), .ZN(n719) );
  XNOR2_X1 U774 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U775 ( .A1(n725), .A2(n720), .ZN(G63) );
  NAND2_X1 U776 ( .A1(n721), .A2(G217), .ZN(n722) );
  XNOR2_X1 U777 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U778 ( .A1(n725), .A2(n724), .ZN(G66) );
  NAND2_X1 U779 ( .A1(G953), .A2(G224), .ZN(n726) );
  XOR2_X1 U780 ( .A(KEYINPUT61), .B(n726), .Z(n727) );
  NOR2_X1 U781 ( .A1(n734), .A2(n727), .ZN(n731) );
  NAND2_X1 U782 ( .A1(n728), .A2(n482), .ZN(n729) );
  XNOR2_X1 U783 ( .A(n729), .B(KEYINPUT125), .ZN(n730) );
  NOR2_X1 U784 ( .A1(n731), .A2(n730), .ZN(n738) );
  XOR2_X1 U785 ( .A(n733), .B(n732), .Z(n736) );
  NAND2_X1 U786 ( .A1(G953), .A2(n734), .ZN(n735) );
  NAND2_X1 U787 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U788 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U789 ( .A(KEYINPUT126), .B(n739), .ZN(G69) );
  XNOR2_X1 U790 ( .A(n741), .B(n740), .ZN(n743) );
  XNOR2_X1 U791 ( .A(n637), .B(n743), .ZN(n742) );
  NAND2_X1 U792 ( .A1(n742), .A2(n482), .ZN(n748) );
  XOR2_X1 U793 ( .A(G227), .B(n743), .Z(n744) );
  NAND2_X1 U794 ( .A1(n744), .A2(G900), .ZN(n745) );
  NAND2_X1 U795 ( .A1(n745), .A2(G953), .ZN(n746) );
  XOR2_X1 U796 ( .A(KEYINPUT127), .B(n746), .Z(n747) );
  NAND2_X1 U797 ( .A1(n748), .A2(n747), .ZN(G72) );
  XOR2_X1 U798 ( .A(n749), .B(G131), .Z(G33) );
  XOR2_X1 U799 ( .A(n750), .B(G122), .Z(G24) );
  XOR2_X1 U800 ( .A(G137), .B(n751), .Z(G39) );
endmodule

