//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n778, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n996, new_n997, new_n998;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT85), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT85), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G29gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  AOI21_X1  g005(.A(KEYINPUT86), .B1(new_n206), .B2(G36gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT86), .ZN(new_n208));
  INV_X1    g007(.A(G36gat), .ZN(new_n209));
  AOI211_X1 g008(.A(new_n208), .B(new_n209), .C1(new_n203), .C2(new_n205), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT88), .B1(new_n207), .B2(new_n210), .ZN(new_n211));
  AND2_X1   g010(.A1(G43gat), .A2(G50gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(G43gat), .A2(G50gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT15), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G43gat), .ZN(new_n215));
  INV_X1    g014(.A(G50gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218));
  NAND2_X1  g017(.A1(G43gat), .A2(G50gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT14), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(new_n202), .A3(new_n209), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n223), .A2(KEYINPUT87), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n227), .B1(KEYINPUT87), .B2(new_n223), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n221), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT85), .B(G29gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n208), .B1(new_n230), .B2(new_n209), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n206), .A2(KEYINPUT86), .A3(G36gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT88), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n211), .A2(new_n229), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT84), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n223), .A2(new_n236), .ZN(new_n237));
  NOR3_X1   g036(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT84), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n226), .A2(KEYINPUT83), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT83), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n241), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n237), .A2(new_n239), .A3(new_n240), .A4(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n243), .A2(new_n232), .A3(new_n231), .ZN(new_n244));
  INV_X1    g043(.A(new_n214), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n235), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G15gat), .B(G22gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT90), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G8gat), .ZN(new_n251));
  INV_X1    g050(.A(G8gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n248), .A2(new_n249), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT16), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n248), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G1gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n251), .A2(new_n257), .A3(new_n256), .A4(new_n253), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n247), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT17), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n233), .B1(new_n231), .B2(new_n232), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT87), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n226), .B1(new_n238), .B2(new_n266), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n214), .B(new_n220), .C1(new_n267), .C2(new_n224), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n269), .A2(new_n234), .B1(new_n245), .B2(new_n244), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n264), .B1(new_n270), .B2(KEYINPUT89), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT89), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n247), .A2(new_n272), .A3(KEYINPUT17), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n261), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n263), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G229gat), .A2(G233gat), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n276), .A2(KEYINPUT91), .A3(KEYINPUT18), .A4(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT17), .B1(new_n247), .B2(new_n272), .ZN(new_n279));
  AOI211_X1 g078(.A(KEYINPUT89), .B(new_n264), .C1(new_n235), .C2(new_n246), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n275), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n281), .A2(KEYINPUT18), .A3(new_n277), .A4(new_n262), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT91), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G113gat), .B(G141gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(G197gat), .ZN(new_n287));
  XOR2_X1   g086(.A(KEYINPUT11), .B(G169gat), .Z(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n290));
  XOR2_X1   g089(.A(new_n289), .B(new_n290), .Z(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n281), .A2(new_n277), .A3(new_n262), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT18), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT92), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(new_n247), .B2(new_n261), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(new_n262), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n277), .B(KEYINPUT13), .Z(new_n298));
  AOI22_X1  g097(.A1(new_n293), .A2(new_n294), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n285), .A2(new_n292), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n292), .B1(new_n285), .B2(new_n299), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G204gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G197gat), .ZN(new_n304));
  INV_X1    g103(.A(G197gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G204gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n304), .A2(new_n306), .A3(KEYINPUT70), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n312), .A2(KEYINPUT71), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(KEYINPUT71), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  XOR2_X1   g115(.A(G211gat), .B(G218gat), .Z(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n316), .A2(KEYINPUT72), .A3(new_n318), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n309), .A2(new_n310), .B1(new_n313), .B2(new_n314), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n317), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G169gat), .ZN(new_n324));
  INV_X1    g123(.A(G176gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327));
  OR3_X1    g126(.A1(new_n326), .A2(KEYINPUT26), .A3(new_n327), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n327), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT27), .B(G183gat), .ZN(new_n330));
  INV_X1    g129(.A(G190gat), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n330), .A2(KEYINPUT28), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT28), .B1(new_n330), .B2(new_n331), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n328), .B(new_n329), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n335), .A2(KEYINPUT24), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n336), .A2(new_n326), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n327), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G183gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n331), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n343), .A2(KEYINPUT24), .A3(new_n335), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n337), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT64), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT25), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n334), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n345), .A2(new_n347), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n337), .A2(new_n341), .A3(KEYINPUT25), .A4(new_n344), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(KEYINPUT64), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT29), .ZN(new_n353));
  NAND2_X1  g152(.A1(G226gat), .A2(G233gat), .ZN(new_n354));
  AOI22_X1  g153(.A1(new_n349), .A2(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n350), .A2(KEYINPUT64), .A3(new_n351), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n334), .A2(new_n348), .ZN(new_n357));
  INV_X1    g156(.A(new_n354), .ZN(new_n358));
  NOR3_X1   g157(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n323), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT73), .ZN(new_n361));
  OAI22_X1  g160(.A1(new_n356), .A2(new_n357), .B1(KEYINPUT29), .B2(new_n358), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n349), .A2(new_n354), .A3(new_n352), .ZN(new_n363));
  INV_X1    g162(.A(new_n323), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n360), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n364), .B1(new_n362), .B2(new_n363), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT73), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G8gat), .B(G36gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(G64gat), .B(G92gat), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n370), .B(new_n371), .Z(new_n372));
  NAND2_X1  g171(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT74), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT30), .ZN(new_n376));
  INV_X1    g175(.A(new_n372), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n377), .B1(new_n366), .B2(new_n368), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT74), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n375), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n369), .A2(new_n372), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n381), .B1(KEYINPUT30), .B2(new_n378), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(G155gat), .ZN(new_n384));
  INV_X1    g183(.A(G162gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G155gat), .A2(G162gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT75), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT75), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n390), .A3(new_n387), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n387), .A2(KEYINPUT2), .ZN(new_n392));
  INV_X1    g191(.A(G141gat), .ZN(new_n393));
  INV_X1    g192(.A(G148gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(G141gat), .A2(G148gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n392), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n389), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n388), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n395), .A2(new_n396), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n399), .A2(new_n400), .A3(new_n390), .A4(new_n392), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(G113gat), .ZN(new_n405));
  INV_X1    g204(.A(G120gat), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT1), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n407), .B1(new_n405), .B2(new_n406), .ZN(new_n408));
  INV_X1    g207(.A(G127gat), .ZN(new_n409));
  INV_X1    g208(.A(G134gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  XOR2_X1   g210(.A(KEYINPUT65), .B(G127gat), .Z(new_n412));
  OAI211_X1 g211(.A(new_n408), .B(new_n411), .C1(new_n410), .C2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G127gat), .B(G134gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT66), .B(G113gat), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n407), .B(new_n414), .C1(new_n415), .C2(new_n406), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n398), .A2(new_n401), .A3(KEYINPUT3), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n404), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT4), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n398), .A2(new_n401), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n420), .B1(new_n421), .B2(new_n417), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n413), .A2(new_n416), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n423), .A2(KEYINPUT4), .A3(new_n402), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n419), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G225gat), .A2(G233gat), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n423), .A2(new_n402), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n421), .A2(new_n417), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n426), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT5), .ZN(new_n431));
  OAI22_X1  g230(.A1(new_n425), .A2(new_n427), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n422), .A2(new_n424), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n433), .A2(KEYINPUT5), .A3(new_n426), .A4(new_n419), .ZN(new_n434));
  XNOR2_X1  g233(.A(G1gat), .B(G29gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n435), .B(KEYINPUT0), .ZN(new_n436));
  XNOR2_X1  g235(.A(G57gat), .B(G85gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n432), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT40), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT39), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n428), .A2(new_n426), .A3(new_n429), .ZN(new_n442));
  AOI211_X1 g241(.A(new_n441), .B(new_n442), .C1(new_n427), .C2(new_n425), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n425), .A2(new_n441), .A3(new_n427), .ZN(new_n444));
  INV_X1    g243(.A(new_n438), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n440), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT81), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  OR3_X1    g248(.A1(new_n443), .A2(new_n440), .A3(new_n446), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n383), .A2(new_n439), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT37), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n372), .B1(new_n369), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n453), .B1(new_n452), .B2(new_n369), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT38), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n438), .B1(new_n432), .B2(new_n434), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT76), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n456), .B(new_n439), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n457), .A2(new_n458), .ZN(new_n460));
  OAI22_X1  g259(.A1(new_n459), .A2(new_n460), .B1(new_n456), .B2(new_n439), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n375), .A2(new_n379), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT38), .ZN(new_n464));
  INV_X1    g263(.A(new_n365), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT37), .B1(new_n465), .B2(new_n367), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n453), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n455), .A2(new_n462), .A3(new_n463), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(G228gat), .A2(G233gat), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n316), .A2(new_n318), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n353), .B1(new_n320), .B2(new_n317), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n403), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n472), .A2(new_n421), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n404), .A2(new_n353), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n474), .A2(new_n323), .ZN(new_n475));
  OAI211_X1 g274(.A(KEYINPUT77), .B(new_n469), .C1(new_n473), .C2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT77), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n472), .A2(new_n421), .B1(new_n474), .B2(new_n323), .ZN(new_n478));
  INV_X1    g277(.A(new_n469), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n403), .B1(new_n323), .B2(KEYINPUT29), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n421), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n475), .A2(new_n469), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n476), .A2(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT78), .B(G22gat), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G78gat), .B(G106gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT31), .B(G50gat), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n487), .B(new_n488), .Z(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT79), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n490), .B1(new_n484), .B2(new_n485), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n480), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n483), .A2(new_n482), .ZN(new_n493));
  AND4_X1   g292(.A1(new_n492), .A2(new_n493), .A3(new_n485), .A4(new_n490), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n486), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n492), .A2(new_n493), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n496), .A2(KEYINPUT80), .A3(G22gat), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT80), .ZN(new_n498));
  INV_X1    g297(.A(G22gat), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n498), .B1(new_n484), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n489), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n497), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n495), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n451), .A2(new_n468), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT34), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n423), .B1(new_n356), .B2(new_n357), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n349), .A2(new_n417), .A3(new_n352), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G227gat), .A2(G233gat), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n510), .ZN(new_n512));
  AOI211_X1 g311(.A(KEYINPUT34), .B(new_n512), .C1(new_n507), .C2(new_n508), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n507), .A2(new_n508), .A3(new_n512), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT32), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT33), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(G15gat), .B(G43gat), .Z(new_n519));
  XNOR2_X1  g318(.A(G71gat), .B(G99gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n516), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n521), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n515), .B(KEYINPUT32), .C1(new_n517), .C2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n514), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n525), .A2(KEYINPUT68), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(KEYINPUT68), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n522), .A2(new_n524), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n511), .A2(new_n513), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT69), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT69), .B1(new_n528), .B2(new_n529), .ZN(new_n531));
  OAI22_X1  g330(.A1(new_n526), .A2(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT36), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT67), .B1(new_n511), .B2(new_n513), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n528), .B(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT36), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n380), .A2(new_n461), .A3(new_n382), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n534), .A2(new_n537), .B1(new_n503), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n505), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT35), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n495), .A2(new_n541), .A3(new_n502), .ZN(new_n542));
  INV_X1    g341(.A(new_n532), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n380), .A2(new_n461), .A3(new_n382), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n495), .A2(new_n502), .A3(new_n536), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT35), .B1(new_n546), .B2(new_n538), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n302), .B1(new_n540), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(new_n384), .ZN(new_n551));
  XNOR2_X1  g350(.A(G183gat), .B(G211gat), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n551), .B(new_n552), .Z(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G57gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(G64gat), .ZN(new_n556));
  INV_X1    g355(.A(G64gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(G57gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT93), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT93), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n556), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G71gat), .A2(G78gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n560), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  OR2_X1    g365(.A1(G71gat), .A2(G78gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n563), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n558), .A2(KEYINPUT94), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT94), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n571), .A2(new_n557), .A3(G57gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n556), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n563), .B1(new_n567), .B2(new_n564), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n566), .A2(new_n569), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT21), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(G127gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n409), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n275), .B1(new_n576), .B2(new_n577), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n584), .B1(new_n582), .B2(new_n583), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n554), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n582), .A2(new_n583), .ZN(new_n588));
  INV_X1    g387(.A(new_n584), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n590), .A2(new_n591), .A3(new_n553), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  AND3_X1   g392(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT97), .B1(G85gat), .B2(G92gat), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT7), .ZN(new_n596));
  OAI22_X1  g395(.A1(new_n594), .A2(new_n595), .B1(KEYINPUT96), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G85gat), .A2(G92gat), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT97), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n596), .A2(KEYINPUT96), .ZN(new_n601));
  NAND3_X1  g400(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G99gat), .A2(G106gat), .ZN(new_n604));
  INV_X1    g403(.A(G85gat), .ZN(new_n605));
  INV_X1    g404(.A(G92gat), .ZN(new_n606));
  AOI22_X1  g405(.A1(KEYINPUT8), .A2(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n597), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT100), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G99gat), .B(G106gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n611), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n608), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(new_n575), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n604), .A2(KEYINPUT8), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n605), .A2(new_n606), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n601), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n600), .A2(new_n602), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n621), .A2(new_n622), .A3(new_n613), .A4(new_n603), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n613), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n611), .A2(KEYINPUT98), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n608), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AOI22_X1  g425(.A1(new_n559), .A2(KEYINPUT93), .B1(new_n564), .B2(new_n563), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n568), .B1(new_n627), .B2(new_n562), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n573), .A2(new_n574), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n623), .B(new_n626), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT10), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n623), .A2(new_n626), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n633), .A2(KEYINPUT10), .A3(new_n575), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G230gat), .A2(G233gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n615), .A2(new_n630), .ZN(new_n638));
  INV_X1    g437(.A(new_n636), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G120gat), .B(G148gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(G176gat), .B(G204gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n642), .B(new_n643), .Z(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n637), .A2(new_n640), .A3(new_n644), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G190gat), .B(G218gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT99), .ZN(new_n651));
  NAND3_X1  g450(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n653), .B1(new_n247), .B2(new_n633), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n279), .A2(new_n280), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n654), .B1(new_n655), .B2(new_n633), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n650), .A2(KEYINPUT99), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT95), .ZN(new_n662));
  XNOR2_X1  g461(.A(G134gat), .B(G162gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n659), .A2(new_n660), .A3(new_n665), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n656), .A2(new_n657), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n664), .B1(new_n667), .B2(new_n658), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n593), .B(new_n649), .C1(new_n666), .C2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT101), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n666), .A2(new_n668), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n673), .A2(KEYINPUT101), .A3(new_n593), .A4(new_n649), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n549), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n461), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(new_n257), .ZN(G1324gat));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n679));
  INV_X1    g478(.A(new_n383), .ZN(new_n680));
  OAI21_X1  g479(.A(G8gat), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT16), .B(G8gat), .Z(new_n682));
  NAND4_X1  g481(.A1(new_n549), .A2(new_n383), .A3(new_n675), .A4(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n679), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n683), .A2(new_n679), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT102), .ZN(G1325gat));
  NAND2_X1  g486(.A1(new_n534), .A2(new_n537), .ZN(new_n688));
  OAI21_X1  g487(.A(G15gat), .B1(new_n676), .B2(new_n688), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n532), .A2(G15gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n689), .B1(new_n676), .B2(new_n690), .ZN(G1326gat));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n504), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT43), .B(G22gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  NOR3_X1   g493(.A1(new_n673), .A2(new_n593), .A3(new_n648), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n549), .A2(new_n695), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n696), .A2(new_n461), .A3(new_n206), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT45), .Z(new_n698));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699));
  AOI211_X1 g498(.A(new_n699), .B(new_n673), .C1(new_n540), .C2(new_n548), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n545), .A2(new_n701), .A3(new_n547), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n545), .B2(new_n547), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n540), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n672), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n700), .B1(new_n705), .B2(new_n699), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(new_n300), .B2(new_n301), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n282), .A2(new_n283), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n282), .A2(new_n283), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n299), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n291), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n285), .A2(new_n292), .A3(new_n299), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(KEYINPUT103), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n708), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n593), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n715), .A2(new_n716), .A3(new_n649), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT104), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n706), .A2(new_n718), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n719), .A2(new_n462), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n698), .B1(new_n720), .B2(new_n230), .ZN(G1328gat));
  NOR3_X1   g520(.A1(new_n696), .A2(G36gat), .A3(new_n680), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT46), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n706), .A2(new_n383), .A3(new_n718), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G36gat), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT106), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n723), .A2(KEYINPUT106), .A3(new_n725), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(G1329gat));
  INV_X1    g529(.A(new_n688), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n719), .A2(G43gat), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n215), .B1(new_n696), .B2(new_n532), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT47), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n732), .A2(new_n736), .A3(new_n733), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n737), .ZN(G1330gat));
  AND3_X1   g537(.A1(new_n495), .A2(new_n536), .A3(new_n502), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n541), .B1(new_n739), .B2(new_n544), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n495), .A2(new_n502), .A3(new_n541), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n741), .A2(new_n538), .A3(new_n532), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT105), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n545), .A2(new_n701), .A3(new_n547), .ZN(new_n744));
  AOI22_X1  g543(.A1(new_n743), .A2(new_n744), .B1(new_n505), .B2(new_n539), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n699), .B1(new_n745), .B2(new_n673), .ZN(new_n746));
  INV_X1    g545(.A(new_n700), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n746), .A2(new_n747), .A3(new_n503), .A4(new_n718), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G50gat), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n549), .A2(new_n216), .A3(new_n503), .A4(new_n695), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n748), .A2(KEYINPUT108), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n706), .A2(new_n755), .A3(new_n503), .A4(new_n718), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n754), .A2(new_n756), .A3(G50gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n750), .A2(KEYINPUT48), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT109), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT109), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n216), .B1(new_n748), .B2(KEYINPUT108), .ZN(new_n762));
  AOI211_X1 g561(.A(new_n761), .B(new_n758), .C1(new_n762), .C2(new_n756), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n753), .B1(new_n760), .B2(new_n763), .ZN(G1331gat));
  NOR4_X1   g563(.A1(new_n715), .A2(new_n716), .A3(new_n672), .A4(new_n649), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT110), .Z(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(new_n745), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n462), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n383), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n771));
  XOR2_X1   g570(.A(KEYINPUT49), .B(G64gat), .Z(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n770), .B2(new_n772), .ZN(G1333gat));
  NAND2_X1  g572(.A1(new_n767), .A2(new_n731), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n532), .A2(G71gat), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n774), .A2(G71gat), .B1(new_n767), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g576(.A1(new_n767), .A2(new_n503), .ZN(new_n778));
  XOR2_X1   g577(.A(KEYINPUT111), .B(G78gat), .Z(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(G1335gat));
  NOR2_X1   g579(.A1(new_n715), .A2(new_n593), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(new_n649), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n706), .A2(new_n462), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n704), .A2(new_n672), .A3(new_n781), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n462), .A2(new_n605), .A3(new_n648), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n790), .B(KEYINPUT112), .Z(new_n791));
  OAI22_X1  g590(.A1(new_n784), .A2(new_n605), .B1(new_n789), .B2(new_n791), .ZN(G1336gat));
  XNOR2_X1  g591(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n785), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n785), .A2(KEYINPUT114), .A3(new_n793), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n796), .B(new_n797), .C1(new_n786), .C2(new_n785), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n680), .A2(G92gat), .A3(new_n649), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n706), .A2(new_n383), .A3(new_n783), .ZN(new_n800));
  AOI22_X1  g599(.A1(new_n798), .A2(new_n799), .B1(G92gat), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802));
  INV_X1    g601(.A(new_n799), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n789), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n800), .A2(G92gat), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n801), .A2(new_n802), .B1(new_n804), .B2(new_n805), .ZN(G1337gat));
  NAND3_X1  g605(.A1(new_n706), .A2(new_n731), .A3(new_n783), .ZN(new_n807));
  XOR2_X1   g606(.A(KEYINPUT115), .B(G99gat), .Z(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n532), .A2(new_n649), .A3(new_n808), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n787), .B2(new_n788), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT116), .ZN(G1338gat));
  NOR3_X1   g612(.A1(new_n504), .A2(G106gat), .A3(new_n649), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n706), .A2(new_n503), .A3(new_n783), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n798), .A2(new_n814), .B1(G106gat), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n817));
  INV_X1    g616(.A(new_n814), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n789), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n815), .A2(G106gat), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n816), .A2(new_n817), .B1(new_n819), .B2(new_n820), .ZN(G1339gat));
  NOR2_X1   g620(.A1(new_n715), .A2(new_n669), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n632), .A2(new_n639), .A3(new_n634), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n639), .B1(new_n632), .B2(new_n634), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n635), .A2(new_n826), .A3(new_n636), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n645), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n823), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g631(.A(KEYINPUT117), .B(new_n823), .C1(new_n827), .C2(new_n829), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n632), .A2(new_n639), .A3(new_n634), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n637), .A2(KEYINPUT54), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n644), .B1(new_n825), .B2(new_n826), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n836), .A2(KEYINPUT55), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n647), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT118), .B1(new_n834), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842));
  AOI211_X1 g641(.A(new_n842), .B(new_n839), .C1(new_n832), .C2(new_n833), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n297), .A2(new_n298), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n276), .A2(new_n277), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n289), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n672), .A2(new_n713), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n713), .A2(new_n648), .A3(new_n847), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n850), .B1(new_n715), .B2(new_n844), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n849), .B1(new_n851), .B2(new_n672), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n822), .B1(new_n852), .B2(new_n716), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n853), .A2(new_n461), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n680), .A3(new_n739), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n855), .B(KEYINPUT119), .Z(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n415), .A3(new_n715), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n680), .A2(new_n462), .ZN(new_n858));
  OR4_X1    g657(.A1(new_n503), .A2(new_n853), .A3(new_n532), .A4(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(G113gat), .B1(new_n859), .B2(new_n302), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n857), .A2(new_n860), .ZN(G1340gat));
  NAND3_X1  g660(.A1(new_n856), .A2(new_n406), .A3(new_n648), .ZN(new_n862));
  OAI21_X1  g661(.A(G120gat), .B1(new_n859), .B2(new_n649), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(G1341gat));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n716), .A2(new_n412), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n865), .B1(new_n859), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n412), .B1(new_n855), .B2(new_n716), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n859), .A2(new_n865), .A3(new_n866), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n869), .A2(new_n870), .ZN(G1342gat));
  OR3_X1    g670(.A1(new_n855), .A2(G134gat), .A3(new_n673), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n873));
  OAI21_X1  g672(.A(G134gat), .B1(new_n859), .B2(new_n673), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(G1343gat));
  NOR3_X1   g675(.A1(new_n731), .A2(new_n383), .A3(new_n504), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n854), .A2(new_n877), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n878), .A2(G141gat), .A3(new_n302), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(KEYINPUT58), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n731), .A2(new_n858), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n883), .B1(new_n853), .B2(new_n504), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n504), .A2(new_n883), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n840), .A2(new_n830), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n886), .B1(new_n712), .B2(new_n713), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n673), .B1(new_n887), .B2(new_n850), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n593), .B1(new_n849), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n885), .B1(new_n889), .B2(new_n822), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n882), .B1(new_n884), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n302), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n880), .B1(new_n893), .B2(new_n393), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n891), .A2(new_n715), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n879), .B1(new_n895), .B2(G141gat), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT58), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(G1344gat));
  INV_X1    g697(.A(new_n878), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(new_n394), .A3(new_n648), .ZN(new_n900));
  AOI211_X1 g699(.A(KEYINPUT59), .B(new_n394), .C1(new_n891), .C2(new_n648), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n839), .B1(new_n832), .B2(new_n833), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n848), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n593), .B1(new_n904), .B2(new_n888), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n671), .A2(new_n674), .A3(new_n302), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n503), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n883), .ZN(new_n908));
  INV_X1    g707(.A(new_n885), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n853), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n648), .A3(new_n881), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n902), .B1(new_n911), .B2(G148gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n900), .B1(new_n901), .B2(new_n912), .ZN(G1345gat));
  NAND3_X1  g712(.A1(new_n899), .A2(new_n384), .A3(new_n593), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n891), .A2(new_n593), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n915), .B2(new_n384), .ZN(G1346gat));
  NOR3_X1   g715(.A1(new_n878), .A2(G162gat), .A3(new_n673), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT121), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n891), .A2(new_n672), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n385), .ZN(G1347gat));
  NAND2_X1  g719(.A1(new_n715), .A2(new_n844), .ZN(new_n921));
  INV_X1    g720(.A(new_n850), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n672), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(new_n849), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n716), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n822), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n680), .A2(new_n462), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n543), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n927), .A2(new_n504), .A3(new_n930), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n931), .A2(new_n324), .A3(new_n302), .ZN(new_n932));
  INV_X1    g731(.A(new_n928), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n853), .A2(new_n546), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(G169gat), .B1(new_n934), .B2(new_n715), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n932), .A2(new_n935), .ZN(G1348gat));
  OAI21_X1  g735(.A(G176gat), .B1(new_n931), .B2(new_n649), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n934), .A2(new_n325), .A3(new_n648), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1349gat));
  OAI21_X1  g738(.A(G183gat), .B1(new_n931), .B2(new_n716), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n934), .A2(new_n330), .A3(new_n593), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT60), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n943), .A2(KEYINPUT122), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n942), .B(new_n944), .ZN(G1350gat));
  NOR4_X1   g744(.A1(new_n853), .A2(new_n503), .A3(new_n673), .A4(new_n929), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT123), .B1(new_n946), .B2(new_n331), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n927), .A2(new_n504), .A3(new_n672), .A4(new_n930), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT123), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n948), .A2(new_n949), .A3(G190gat), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n947), .A2(KEYINPUT61), .A3(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n952));
  OAI211_X1 g751(.A(KEYINPUT123), .B(new_n952), .C1(new_n946), .C2(new_n331), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n934), .A2(new_n331), .A3(new_n672), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(KEYINPUT124), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n947), .A2(KEYINPUT61), .A3(new_n950), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n957), .A2(new_n958), .A3(new_n953), .A4(new_n954), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n956), .A2(new_n959), .ZN(G1351gat));
  AOI21_X1  g759(.A(new_n909), .B1(new_n925), .B2(new_n926), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n904), .A2(new_n888), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(new_n716), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n671), .A2(new_n674), .A3(new_n302), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT57), .B1(new_n965), .B2(new_n503), .ZN(new_n966));
  OAI21_X1  g765(.A(KEYINPUT126), .B1(new_n961), .B2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n908), .B(new_n968), .C1(new_n853), .C2(new_n909), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n731), .A2(new_n933), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n967), .A2(new_n892), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(G197gat), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n853), .A2(new_n933), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n731), .A2(new_n504), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n973), .A2(KEYINPUT125), .A3(new_n974), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n977), .A2(new_n305), .A3(new_n715), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n972), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(KEYINPUT127), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n972), .A2(new_n982), .A3(new_n979), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n981), .A2(new_n983), .ZN(G1352gat));
  NOR3_X1   g783(.A1(new_n975), .A2(G204gat), .A3(new_n649), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT62), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n967), .A2(new_n969), .A3(new_n970), .ZN(new_n987));
  AND2_X1   g786(.A1(new_n987), .A2(new_n648), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n986), .B1(new_n988), .B2(new_n303), .ZN(G1353gat));
  NOR2_X1   g788(.A1(new_n716), .A2(G211gat), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n977), .A2(new_n978), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n910), .A2(new_n593), .A3(new_n970), .ZN(new_n992));
  AND3_X1   g791(.A1(new_n992), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n993));
  AOI21_X1  g792(.A(KEYINPUT63), .B1(new_n992), .B2(G211gat), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(G1354gat));
  INV_X1    g794(.A(G218gat), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n977), .A2(new_n672), .A3(new_n978), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n673), .A2(new_n996), .ZN(new_n998));
  AOI22_X1  g797(.A1(new_n996), .A2(new_n997), .B1(new_n987), .B2(new_n998), .ZN(G1355gat));
endmodule


