//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1211, new_n1212, new_n1213,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT65), .Z(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n223), .A2(new_n224), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n209), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(new_n207), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT64), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n229), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  AND3_X1   g0034(.A1(new_n225), .A2(new_n226), .A3(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G226), .B(G232), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  INV_X1    g0047(.A(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT68), .B(G50), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  INV_X1    g0055(.A(new_n230), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT3), .B(G33), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(G222), .A3(new_n260), .ZN(new_n261));
  XOR2_X1   g0061(.A(new_n261), .B(KEYINPUT70), .Z(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(G1698), .ZN(new_n263));
  INV_X1    g0063(.A(G223), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n265), .B1(G77), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n258), .B1(new_n262), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n257), .A2(KEYINPUT69), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT69), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G33), .A3(G41), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(new_n275), .A3(new_n256), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  INV_X1    g0077(.A(G45), .ZN(new_n278));
  AOI21_X1  g0078(.A(G1), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n276), .A2(G274), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n279), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G226), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n280), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n272), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G169), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n230), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n206), .A2(G20), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(G50), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT8), .B(G58), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n207), .A2(G33), .ZN(new_n297));
  INV_X1    g0097(.A(G150), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G20), .A2(G33), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n296), .A2(new_n297), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(G20), .B2(new_n203), .ZN(new_n302));
  INV_X1    g0102(.A(new_n292), .ZN(new_n303));
  OAI221_X1 g0103(.A(new_n295), .B1(G50), .B2(new_n289), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G179), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n285), .A2(new_n305), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n288), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n285), .A2(G190), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT72), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n286), .A2(G200), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n304), .B(KEYINPUT9), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n311), .B(KEYINPUT71), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT10), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n314), .A2(new_n309), .A3(new_n315), .A4(new_n310), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n307), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n293), .A2(G68), .A3(new_n294), .ZN(new_n318));
  XOR2_X1   g0118(.A(new_n318), .B(KEYINPUT74), .Z(new_n319));
  NAND2_X1  g0119(.A1(new_n299), .A2(G50), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT73), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n320), .B(new_n321), .ZN(new_n322));
  OAI22_X1  g0122(.A1(new_n297), .A2(new_n217), .B1(new_n207), .B2(G68), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n292), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT11), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n324), .A2(new_n325), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n289), .A2(G68), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT12), .ZN(new_n329));
  NOR4_X1   g0129(.A1(new_n319), .A2(new_n326), .A3(new_n327), .A4(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G190), .ZN(new_n331));
  MUX2_X1   g0131(.A(G226), .B(G232), .S(G1698), .Z(new_n332));
  AOI22_X1  g0132(.A1(new_n332), .A2(new_n259), .B1(G33), .B2(G97), .ZN(new_n333));
  OAI221_X1 g0133(.A(new_n280), .B1(new_n282), .B2(new_n212), .C1(new_n333), .C2(new_n258), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n334), .A2(KEYINPUT13), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(KEYINPUT13), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n330), .B1(new_n331), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G200), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n339), .B1(new_n335), .B2(new_n336), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT75), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n337), .B2(new_n305), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n335), .A2(KEYINPUT75), .A3(G179), .A4(new_n336), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n337), .A2(G169), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT14), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT14), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n337), .A2(new_n348), .A3(G169), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n345), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n330), .B(KEYINPUT76), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n341), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n259), .A2(G232), .A3(new_n260), .ZN(new_n353));
  OAI221_X1 g0153(.A(new_n353), .B1(new_n219), .B2(new_n259), .C1(new_n263), .C2(new_n212), .ZN(new_n354));
  INV_X1    g0154(.A(new_n258), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n356), .B(new_n280), .C1(new_n218), .C2(new_n282), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G200), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n293), .A2(G77), .A3(new_n294), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(G77), .B2(new_n289), .ZN(new_n360));
  INV_X1    g0160(.A(new_n296), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n361), .A2(new_n299), .B1(G20), .B2(G77), .ZN(new_n362));
  XNOR2_X1  g0162(.A(KEYINPUT15), .B(G87), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n362), .B1(new_n297), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n360), .B1(new_n292), .B2(new_n364), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n358), .B(new_n365), .C1(new_n331), .C2(new_n357), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n365), .B1(new_n357), .B2(new_n287), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(G179), .B2(new_n357), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n317), .A2(new_n352), .A3(new_n366), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n283), .A2(G1698), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(G223), .B2(G1698), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n266), .A2(KEYINPUT77), .A3(G33), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT77), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n267), .A2(new_n269), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n371), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n268), .A2(new_n213), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n355), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n276), .A2(G232), .A3(new_n281), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n280), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(new_n379), .A3(new_n331), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n380), .A2(KEYINPUT80), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT80), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n280), .A2(new_n378), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n266), .A2(KEYINPUT77), .A3(G33), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n259), .B2(new_n373), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n385), .A2(new_n371), .B1(new_n268), .B2(new_n213), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n383), .B1(new_n386), .B2(new_n355), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n382), .B1(new_n387), .B2(new_n331), .ZN(new_n388));
  AOI21_X1  g0188(.A(G200), .B1(new_n377), .B2(new_n379), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n381), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n248), .A2(new_n211), .ZN(new_n392));
  OAI21_X1  g0192(.A(G20), .B1(new_n392), .B2(new_n201), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n299), .A2(G159), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(new_n385), .B2(new_n207), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n374), .A2(new_n397), .A3(new_n207), .A4(new_n372), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G68), .ZN(new_n400));
  OAI211_X1 g0200(.A(KEYINPUT16), .B(new_n396), .C1(new_n398), .C2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT16), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n397), .B1(new_n259), .B2(G20), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n270), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n211), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n402), .B1(new_n405), .B2(new_n395), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n401), .A2(new_n406), .A3(new_n292), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n361), .A2(new_n294), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n303), .A2(new_n289), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n408), .A2(new_n409), .B1(new_n289), .B2(new_n361), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT78), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n410), .B(new_n411), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT17), .B1(new_n391), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n387), .A2(new_n382), .A3(new_n331), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n380), .A2(KEYINPUT80), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n415), .B1(new_n416), .B2(new_n389), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n407), .A2(new_n412), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT17), .ZN(new_n419));
  NOR3_X1   g0219(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n414), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n377), .A2(new_n379), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(G169), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n305), .B2(new_n422), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT18), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n418), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(new_n418), .B2(new_n424), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT79), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n418), .A2(new_n424), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT18), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT79), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n418), .A2(new_n424), .A3(new_n425), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n421), .A2(new_n428), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n369), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n206), .A2(G45), .ZN(new_n436));
  OR2_X1    g0236(.A1(KEYINPUT5), .A2(G41), .ZN(new_n437));
  NAND2_X1  g0237(.A1(KEYINPUT5), .A2(G41), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n439), .A2(new_n276), .A3(G274), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n278), .A2(G1), .ZN(new_n441));
  INV_X1    g0241(.A(new_n438), .ZN(new_n442));
  NOR2_X1   g0242(.A1(KEYINPUT5), .A2(G41), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n276), .A2(new_n444), .A3(G257), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n259), .A2(KEYINPUT4), .A3(G244), .A4(new_n260), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n259), .A2(G250), .A3(G1698), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G283), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n260), .A2(G244), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(new_n374), .B2(new_n372), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT4), .B1(new_n453), .B2(KEYINPUT83), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT83), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(new_n385), .B2(new_n452), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n451), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n447), .B1(new_n457), .B2(new_n258), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT84), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(KEYINPUT84), .B(new_n447), .C1(new_n457), .C2(new_n258), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(G200), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n206), .A2(G33), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n289), .A2(new_n463), .A3(new_n230), .A4(new_n291), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  OR3_X1    g0265(.A1(new_n289), .A2(KEYINPUT82), .A3(G97), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT82), .B1(new_n289), .B2(G97), .ZN(new_n467));
  AOI22_X1  g0267(.A1(G97), .A2(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n219), .B1(new_n403), .B2(new_n404), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT6), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n470), .A2(KEYINPUT81), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n470), .A2(KEYINPUT81), .ZN(new_n472));
  INV_X1    g0272(.A(G97), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(new_n219), .ZN(new_n474));
  NOR2_X1   g0274(.A1(G97), .A2(G107), .ZN(new_n475));
  OAI22_X1  g0275(.A1(new_n471), .A2(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(G97), .A3(new_n219), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n207), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n300), .A2(new_n217), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n469), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n468), .B1(new_n481), .B2(new_n303), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n454), .A2(new_n456), .ZN(new_n483));
  INV_X1    g0283(.A(new_n451), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n446), .B1(new_n485), .B2(new_n355), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n482), .B1(new_n486), .B2(G190), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n462), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n458), .A2(new_n287), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n305), .B(new_n447), .C1(new_n457), .C2(new_n258), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(new_n482), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n212), .A2(new_n260), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n218), .A2(G1698), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n374), .B2(new_n372), .ZN(new_n495));
  INV_X1    g0295(.A(G116), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n268), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT85), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT85), .ZN(new_n499));
  INV_X1    g0299(.A(new_n497), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n499), .B(new_n500), .C1(new_n385), .C2(new_n494), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n498), .A2(new_n501), .A3(new_n355), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n436), .A2(G274), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n214), .B2(new_n436), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n276), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n502), .A2(new_n305), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(G169), .B1(new_n502), .B2(new_n505), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT86), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n502), .A2(new_n305), .A3(new_n505), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT86), .ZN(new_n510));
  INV_X1    g0310(.A(new_n505), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n374), .A2(new_n372), .ZN(new_n512));
  INV_X1    g0312(.A(new_n494), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n497), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n258), .B1(new_n514), .B2(new_n499), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n511), .B1(new_n515), .B2(new_n498), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n509), .B(new_n510), .C1(new_n516), .C2(G169), .ZN(new_n517));
  XNOR2_X1  g0317(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n518), .A2(new_n207), .A3(G33), .A4(G97), .ZN(new_n519));
  NOR3_X1   g0319(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n520));
  AOI21_X1  g0320(.A(G20), .B1(G33), .B2(G97), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n519), .B1(new_n522), .B2(new_n518), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n512), .A2(new_n207), .A3(G68), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n292), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n363), .A2(new_n290), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n526), .B(new_n527), .C1(new_n363), .C2(new_n464), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n508), .A2(new_n517), .A3(new_n528), .ZN(new_n529));
  OR3_X1    g0329(.A1(new_n464), .A2(KEYINPUT88), .A3(new_n213), .ZN(new_n530));
  OAI21_X1  g0330(.A(KEYINPUT88), .B1(new_n464), .B2(new_n213), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n526), .A2(new_n527), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n533), .B1(G190), .B2(new_n516), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n339), .B2(new_n516), .ZN(new_n535));
  AND4_X1   g0335(.A1(new_n488), .A2(new_n491), .A3(new_n529), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n214), .A2(new_n260), .ZN(new_n537));
  INV_X1    g0337(.A(G257), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G1698), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n374), .B2(new_n372), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G294), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n355), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n276), .A2(new_n444), .A3(G264), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(new_n440), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n287), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(G179), .B2(new_n546), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n290), .A2(KEYINPUT25), .A3(new_n219), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT25), .B1(new_n290), .B2(new_n219), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n549), .A2(new_n550), .B1(new_n219), .B2(new_n464), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n512), .A2(KEYINPUT22), .A3(new_n207), .A4(G87), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT24), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT22), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n207), .A2(G87), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n554), .B1(new_n270), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT23), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n207), .B2(G107), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n219), .A2(KEYINPUT23), .A3(G20), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n558), .A2(new_n559), .B1(new_n497), .B2(new_n207), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n552), .A2(new_n553), .A3(new_n556), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(KEYINPUT22), .A2(G87), .ZN(new_n562));
  AOI211_X1 g0362(.A(G20), .B(new_n562), .C1(new_n374), .C2(new_n372), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n556), .A2(new_n560), .ZN(new_n564));
  OAI21_X1  g0364(.A(KEYINPUT24), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n551), .B1(new_n566), .B2(new_n292), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n548), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n545), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n542), .B1(new_n385), .B2(new_n540), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n570), .B1(new_n571), .B2(new_n355), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT90), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n572), .A2(new_n573), .A3(new_n331), .A4(new_n440), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n544), .A2(new_n331), .A3(new_n440), .A4(new_n545), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT90), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n546), .A2(new_n339), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n578), .A2(KEYINPUT91), .A3(new_n567), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT91), .B1(new_n578), .B2(new_n567), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n569), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT21), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n276), .A2(new_n444), .A3(G270), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n440), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n538), .A2(new_n260), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n220), .A2(G1698), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n374), .B2(new_n372), .ZN(new_n588));
  INV_X1    g0388(.A(G303), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n259), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n355), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n584), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G169), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n290), .A2(new_n496), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n464), .B2(new_n496), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n450), .B(new_n207), .C1(G33), .C2(new_n473), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n596), .B(new_n292), .C1(new_n207), .C2(G116), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT20), .ZN(new_n598));
  OR2_X1    g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n598), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n595), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n582), .B1(new_n593), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n592), .A2(G200), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n603), .B(new_n601), .C1(new_n331), .C2(new_n592), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n592), .A2(KEYINPUT21), .A3(G169), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n584), .A2(G179), .A3(new_n591), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n601), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(KEYINPUT89), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT89), .ZN(new_n609));
  AOI211_X1 g0409(.A(new_n609), .B(new_n601), .C1(new_n605), .C2(new_n606), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n602), .B(new_n604), .C1(new_n608), .C2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n581), .A2(new_n611), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n435), .A2(new_n536), .A3(new_n612), .ZN(G372));
  INV_X1    g0413(.A(new_n491), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT92), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n502), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n515), .A2(KEYINPUT92), .A3(new_n498), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n511), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n534), .B1(new_n618), .B2(new_n339), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n509), .B(new_n528), .C1(new_n618), .C2(G169), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n614), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT26), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n614), .A2(new_n529), .A3(new_n535), .A4(KEYINPUT26), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n607), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n602), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n488), .B(new_n491), .C1(new_n628), .C2(new_n568), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n619), .B1(new_n579), .B2(new_n580), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n620), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n435), .B1(new_n626), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n430), .A2(new_n432), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n341), .A2(new_n368), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n635), .B1(new_n351), .B2(new_n350), .ZN(new_n636));
  INV_X1    g0436(.A(new_n421), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n313), .A2(new_n316), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n307), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n632), .A2(new_n640), .ZN(G369));
  INV_X1    g0441(.A(new_n581), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n645), .A3(G213), .ZN(new_n646));
  INV_X1    g0446(.A(G343), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n642), .B1(new_n567), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(new_n569), .B2(new_n649), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n601), .A2(new_n649), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n628), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n611), .B2(new_n652), .ZN(new_n654));
  XNOR2_X1  g0454(.A(KEYINPUT93), .B(G330), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n608), .A2(new_n610), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n648), .B1(new_n659), .B2(new_n602), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n660), .A2(new_n642), .B1(new_n568), .B2(new_n649), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n658), .A2(new_n661), .ZN(G399));
  INV_X1    g0462(.A(new_n227), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(G41), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n520), .A2(new_n496), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n664), .A2(new_n665), .A3(new_n206), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n666), .B1(new_n233), .B2(new_n664), .ZN(new_n667));
  XOR2_X1   g0467(.A(new_n667), .B(KEYINPUT28), .Z(new_n668));
  NAND3_X1  g0468(.A1(new_n612), .A2(new_n536), .A3(new_n649), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT31), .ZN(new_n670));
  AOI21_X1  g0470(.A(KEYINPUT92), .B1(new_n515), .B2(new_n498), .ZN(new_n671));
  AND4_X1   g0471(.A1(KEYINPUT92), .A2(new_n498), .A3(new_n501), .A4(new_n355), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n505), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n592), .A2(new_n546), .A3(new_n305), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n458), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT30), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n584), .A2(G179), .A3(new_n591), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n677), .A2(new_n502), .A3(new_n505), .A4(new_n572), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n676), .B1(new_n678), .B2(new_n458), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n678), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT95), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n681), .A2(new_n682), .A3(KEYINPUT30), .A4(new_n486), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n544), .A2(new_n545), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n606), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n486), .A2(KEYINPUT30), .A3(new_n516), .A4(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT95), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n680), .B1(new_n683), .B2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n670), .B1(new_n688), .B2(new_n649), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n680), .A2(KEYINPUT94), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n683), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT94), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n675), .A2(new_n679), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n690), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n649), .A2(new_n670), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n669), .A2(new_n689), .A3(new_n696), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n697), .A2(KEYINPUT96), .A3(new_n655), .ZN(new_n698));
  AOI21_X1  g0498(.A(KEYINPUT96), .B1(new_n697), .B2(new_n655), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n620), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(new_n621), .B2(KEYINPUT26), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n614), .A2(new_n529), .A3(new_n535), .A4(new_n622), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n614), .B1(new_n462), .B2(new_n487), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n569), .B(new_n602), .C1(new_n608), .C2(new_n610), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI211_X1 g0506(.A(new_n702), .B(new_n703), .C1(new_n706), .C2(new_n630), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n707), .A2(KEYINPUT29), .A3(new_n649), .ZN(new_n708));
  INV_X1    g0508(.A(new_n631), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n648), .B1(new_n709), .B2(new_n625), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n708), .B1(new_n710), .B2(KEYINPUT29), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n700), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n668), .B1(new_n713), .B2(G1), .ZN(G364));
  INV_X1    g0514(.A(new_n664), .ZN(new_n715));
  INV_X1    g0515(.A(G13), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G20), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n206), .B1(new_n717), .B2(G45), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n715), .A2(KEYINPUT97), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT97), .ZN(new_n720));
  INV_X1    g0520(.A(new_n718), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n720), .B1(new_n664), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n657), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(new_n655), .B2(new_n654), .ZN(new_n726));
  NOR2_X1   g0526(.A1(G13), .A2(G33), .ZN(new_n727));
  XOR2_X1   g0527(.A(new_n727), .B(KEYINPUT98), .Z(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G20), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n230), .B1(G20), .B2(new_n287), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n233), .A2(new_n278), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n385), .A2(new_n227), .ZN(new_n733));
  AOI211_X1 g0533(.A(new_n732), .B(new_n733), .C1(new_n251), .C2(G45), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n663), .A2(new_n270), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G355), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(G116), .B2(new_n227), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n731), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n207), .A2(new_n305), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n339), .A2(G190), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G190), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n211), .A2(new_n741), .B1(new_n743), .B2(new_n217), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n739), .A2(G190), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n339), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(G200), .ZN(new_n747));
  AOI22_X1  g0547(.A1(G50), .A2(new_n746), .B1(new_n747), .B2(G58), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n207), .A2(G179), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n742), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G159), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n331), .A2(G179), .A3(G200), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n207), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n748), .B1(KEYINPUT32), .B2(new_n752), .C1(new_n473), .C2(new_n754), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n744), .B(new_n755), .C1(KEYINPUT32), .C2(new_n752), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n740), .A2(new_n749), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n219), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n749), .A2(G190), .A3(G200), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n270), .B(new_n758), .C1(G87), .C2(new_n760), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT99), .Z(new_n762));
  INV_X1    g0562(.A(new_n741), .ZN(new_n763));
  INV_X1    g0563(.A(G317), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(KEYINPUT33), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n764), .A2(KEYINPUT33), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n763), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n747), .ZN(new_n768));
  INV_X1    g0568(.A(G322), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT100), .Z(new_n771));
  INV_X1    g0571(.A(G283), .ZN(new_n772));
  INV_X1    g0572(.A(G294), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n270), .B1(new_n757), .B2(new_n772), .C1(new_n754), .C2(new_n773), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n760), .A2(G303), .B1(new_n751), .B2(G329), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n775), .B1(new_n776), .B2(new_n743), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n774), .B(new_n777), .C1(G326), .C2(new_n746), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n756), .A2(new_n762), .B1(new_n771), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n730), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n738), .B(new_n724), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT101), .ZN(new_n782));
  INV_X1    g0582(.A(new_n729), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n782), .B1(new_n654), .B2(new_n783), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n726), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(G396));
  OAI21_X1  g0586(.A(new_n366), .B1(new_n365), .B2(new_n649), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n368), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n368), .A2(new_n648), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n710), .B(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n724), .B1(new_n792), .B2(new_n700), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n700), .B2(new_n792), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n730), .A2(new_n727), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n723), .B1(new_n217), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n743), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G116), .A2(new_n797), .B1(new_n763), .B2(G283), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n799), .A2(KEYINPUT102), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(KEYINPUT102), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n270), .B1(new_n759), .B2(new_n219), .ZN(new_n802));
  INV_X1    g0602(.A(new_n757), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G87), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n776), .B2(new_n750), .ZN(new_n805));
  NOR4_X1   g0605(.A1(new_n800), .A2(new_n801), .A3(new_n802), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n754), .A2(new_n473), .ZN(new_n807));
  INV_X1    g0607(.A(new_n746), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n589), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n807), .B(new_n809), .C1(G294), .C2(new_n747), .ZN(new_n810));
  AOI22_X1  g0610(.A1(G150), .A2(new_n763), .B1(new_n797), .B2(G159), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n747), .A2(G143), .ZN(new_n812));
  INV_X1    g0612(.A(G137), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n811), .B(new_n812), .C1(new_n813), .C2(new_n808), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT34), .ZN(new_n815));
  INV_X1    g0615(.A(G132), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n757), .A2(new_n211), .B1(new_n750), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n512), .B1(new_n248), .B2(new_n754), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n817), .B(new_n818), .C1(G50), .C2(new_n760), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n806), .A2(new_n810), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n796), .B1(new_n780), .B2(new_n820), .C1(new_n791), .C2(new_n728), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n794), .A2(new_n821), .ZN(G384));
  NOR2_X1   g0622(.A1(new_n717), .A2(new_n206), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT103), .ZN(new_n824));
  INV_X1    g0624(.A(new_n695), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n688), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n691), .ZN(new_n827));
  OAI211_X1 g0627(.A(KEYINPUT103), .B(new_n695), .C1(new_n827), .C2(new_n680), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n669), .A2(new_n689), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n350), .A2(new_n351), .ZN(new_n830));
  INV_X1    g0630(.A(new_n341), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n351), .A2(new_n648), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n351), .B(new_n648), .C1(new_n350), .C2(new_n341), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n790), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n410), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n398), .A2(new_n400), .ZN(new_n837));
  AOI21_X1  g0637(.A(KEYINPUT16), .B1(new_n837), .B2(new_n396), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n401), .A2(new_n292), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n646), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n434), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n391), .A2(new_n413), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n418), .A2(new_n841), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT37), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n845), .A2(new_n429), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n840), .A2(new_n424), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n845), .A2(new_n849), .A3(new_n842), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n848), .B1(new_n850), .B2(new_n847), .ZN(new_n851));
  AND3_X1   g0651(.A1(new_n844), .A2(KEYINPUT38), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT38), .B1(new_n844), .B2(new_n851), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n829), .B(new_n835), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT40), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT104), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n854), .A2(KEYINPUT104), .A3(new_n855), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n835), .A2(new_n829), .A3(KEYINPUT40), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n845), .A2(new_n429), .A3(new_n846), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(new_n847), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n846), .B1(new_n634), .B2(new_n421), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n844), .A2(KEYINPUT38), .A3(new_n851), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n861), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n860), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n435), .A2(new_n829), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n870), .A2(new_n871), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n872), .A2(new_n655), .A3(new_n873), .ZN(new_n874));
  OR3_X1    g0674(.A1(new_n711), .A2(new_n434), .A3(new_n369), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n640), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT39), .B1(new_n866), .B2(new_n867), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n853), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(KEYINPUT39), .A3(new_n867), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n350), .A2(new_n351), .A3(new_n649), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n878), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n649), .B(new_n791), .C1(new_n626), .C2(new_n631), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n789), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n833), .A2(new_n834), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n885), .B(new_n886), .C1(new_n852), .C2(new_n853), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n633), .A2(new_n646), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n883), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n876), .B(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n823), .B1(new_n874), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n890), .B2(new_n874), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n476), .A2(new_n478), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n893), .A2(KEYINPUT35), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(KEYINPUT35), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n894), .A2(G116), .A3(new_n231), .A4(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT36), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n233), .B(G77), .C1(new_n248), .C2(new_n211), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(G50), .B2(new_n211), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(G1), .A3(new_n716), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n892), .A2(new_n897), .A3(new_n900), .ZN(G367));
  INV_X1    g0701(.A(new_n482), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n704), .B1(new_n902), .B2(new_n649), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n614), .A2(new_n648), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(new_n642), .A3(new_n660), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n906), .A2(KEYINPUT42), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n488), .A2(new_n568), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n648), .B1(new_n908), .B2(new_n491), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(new_n906), .B2(KEYINPUT42), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n533), .A2(new_n648), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n619), .A2(new_n620), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n620), .B2(new_n911), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n907), .A2(new_n910), .B1(KEYINPUT43), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n913), .A2(KEYINPUT43), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n914), .B(new_n915), .Z(new_n916));
  INV_X1    g0716(.A(new_n905), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n658), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n916), .B(new_n918), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n664), .B(KEYINPUT41), .Z(new_n920));
  INV_X1    g0720(.A(new_n661), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT44), .B1(new_n921), .B2(new_n917), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT44), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n661), .A2(new_n905), .A3(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g0725(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n921), .B2(new_n917), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n661), .A2(new_n905), .A3(new_n926), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n925), .A2(new_n930), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n931), .A2(new_n658), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n658), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n660), .A2(new_n642), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n651), .B2(new_n660), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(new_n656), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n712), .A2(new_n937), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n938), .A2(KEYINPUT106), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(KEYINPUT106), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n934), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n920), .B1(new_n941), .B2(new_n713), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n919), .B1(new_n942), .B2(new_n721), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n731), .B1(new_n227), .B2(new_n363), .C1(new_n245), .C2(new_n733), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT107), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n723), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n945), .B2(new_n944), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n754), .A2(new_n211), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n270), .B(new_n948), .C1(G159), .C2(new_n763), .ZN(new_n949));
  AOI22_X1  g0749(.A1(G50), .A2(new_n797), .B1(new_n751), .B2(G137), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n760), .A2(G58), .B1(new_n803), .B2(G77), .ZN(new_n951));
  AOI22_X1  g0751(.A1(G143), .A2(new_n746), .B1(new_n747), .B2(G150), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n949), .A2(new_n950), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n768), .A2(new_n589), .B1(new_n219), .B2(new_n754), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n759), .A2(new_n496), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n954), .B1(KEYINPUT46), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n757), .A2(new_n473), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n741), .A2(new_n773), .B1(new_n750), .B2(new_n764), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n957), .B(new_n958), .C1(G283), .C2(new_n797), .ZN(new_n959));
  XOR2_X1   g0759(.A(KEYINPUT108), .B(G311), .Z(new_n960));
  AOI21_X1  g0760(.A(new_n512), .B1(new_n746), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n956), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n759), .B2(new_n496), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT110), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n953), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT47), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n947), .B1(new_n967), .B2(new_n730), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n913), .B2(new_n783), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n943), .A2(new_n969), .ZN(G387));
  NAND2_X1  g0770(.A1(new_n939), .A2(new_n940), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n715), .B1(new_n712), .B2(new_n937), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n385), .B(new_n957), .C1(G150), .C2(new_n751), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n754), .A2(new_n363), .ZN(new_n975));
  AOI22_X1  g0775(.A1(G50), .A2(new_n747), .B1(new_n746), .B2(G159), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n217), .A2(new_n759), .B1(new_n743), .B2(new_n211), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n361), .B2(new_n763), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n974), .A2(new_n975), .A3(new_n976), .A4(new_n978), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n803), .A2(G116), .B1(new_n751), .B2(G326), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G303), .A2(new_n797), .B1(new_n763), .B2(new_n960), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n768), .B2(new_n764), .C1(new_n769), .C2(new_n808), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT48), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n983), .ZN(new_n985));
  INV_X1    g0785(.A(new_n754), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n986), .A2(G283), .B1(new_n760), .B2(G294), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n984), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT49), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n385), .B(new_n980), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n988), .A2(new_n989), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n979), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n730), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n735), .A2(new_n665), .B1(new_n219), .B2(new_n663), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n241), .A2(new_n278), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n296), .A2(G50), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT50), .ZN(new_n997));
  AOI211_X1 g0797(.A(G45), .B(new_n665), .C1(G68), .C2(G77), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n733), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT111), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n994), .B1(new_n995), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n723), .B1(new_n1001), .B2(new_n731), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n993), .B(new_n1002), .C1(new_n651), .C2(new_n783), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n973), .B(new_n1003), .C1(new_n718), .C2(new_n937), .ZN(G393));
  OAI221_X1 g0804(.A(new_n731), .B1(new_n473), .B2(new_n227), .C1(new_n254), .C2(new_n733), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n724), .A2(new_n1005), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n202), .A2(new_n741), .B1(new_n743), .B2(new_n296), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n754), .A2(new_n217), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1009), .A2(KEYINPUT112), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n804), .B1(new_n211), .B2(new_n759), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G143), .B2(new_n751), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1009), .A2(KEYINPUT112), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1010), .A2(new_n1012), .A3(new_n512), .A4(new_n1013), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G150), .A2(new_n746), .B1(new_n747), .B2(G159), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT51), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G311), .A2(new_n747), .B1(new_n746), .B2(G317), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT52), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n259), .B(new_n758), .C1(G116), .C2(new_n986), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G294), .A2(new_n797), .B1(new_n763), .B2(G303), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n760), .A2(G283), .B1(new_n751), .B2(G322), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n1014), .A2(new_n1016), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1006), .B1(new_n1023), .B2(new_n730), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n905), .B2(new_n783), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n932), .A2(new_n933), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1025), .B1(new_n1026), .B2(new_n718), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT113), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n941), .A2(new_n664), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n934), .B1(new_n939), .B2(new_n940), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n1029), .A2(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(G390));
  INV_X1    g0833(.A(new_n886), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n884), .B2(new_n789), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT39), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n852), .A2(new_n853), .A3(new_n1036), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n1035), .A2(new_n882), .B1(new_n1037), .B2(new_n877), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n707), .A2(new_n649), .A3(new_n788), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n789), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n886), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n882), .B1(new_n866), .B2(new_n867), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n835), .B1(new_n698), .B2(new_n699), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1038), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1038), .A2(new_n1043), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n829), .A2(G330), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n835), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1045), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n721), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n728), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n1037), .B2(new_n877), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n723), .B1(new_n296), .B2(new_n795), .ZN(new_n1054));
  INV_X1    g0854(.A(G159), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n768), .A2(new_n816), .B1(new_n1055), .B2(new_n754), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n760), .A2(G150), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT53), .ZN(new_n1058));
  INV_X1    g0858(.A(G128), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n259), .B1(new_n757), .B2(new_n202), .C1(new_n808), .C2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(KEYINPUT54), .B(G143), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G137), .A2(new_n763), .B1(new_n797), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(G125), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1063), .B1(new_n1064), .B2(new_n750), .ZN(new_n1065));
  OR4_X1    g0865(.A1(new_n1056), .A2(new_n1058), .A3(new_n1060), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1008), .B1(G116), .B2(new_n747), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n772), .B2(new_n808), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n473), .A2(new_n743), .B1(new_n741), .B2(new_n219), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT118), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n259), .B1(new_n760), .B2(G87), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n803), .A2(G68), .B1(new_n751), .B2(G294), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1066), .B1(new_n1068), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1076), .A2(KEYINPUT119), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(KEYINPUT119), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n730), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1053), .B(new_n1054), .C1(new_n1077), .C2(new_n1079), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1051), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n829), .A2(G330), .A3(new_n791), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n1034), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(KEYINPUT114), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1040), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT114), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1082), .A2(new_n1086), .A3(new_n1034), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1084), .A2(new_n1044), .A3(new_n1085), .A4(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(KEYINPUT115), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n697), .A2(new_n655), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT96), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n697), .A2(KEYINPUT96), .A3(new_n655), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1040), .B1(new_n1094), .B2(new_n835), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT115), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1095), .A2(new_n1096), .A3(new_n1087), .A4(new_n1084), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1089), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n885), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n791), .B1(new_n698), .B2(new_n699), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n1034), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1099), .B1(new_n1101), .B2(new_n1048), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1098), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n435), .A2(new_n1047), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n875), .A2(new_n640), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT116), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1045), .B(new_n1109), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n1038), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1048), .B1(new_n1038), .B2(new_n1043), .ZN(new_n1112));
  OAI21_X1  g0912(.A(KEYINPUT116), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n715), .B1(new_n1108), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1106), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n1050), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT117), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1102), .B1(new_n1089), .B2(new_n1097), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1113), .B(new_n1110), .C1(new_n1119), .C2(new_n1106), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1117), .A2(new_n1120), .A3(KEYINPUT117), .A4(new_n664), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1081), .B1(new_n1118), .B2(new_n1122), .ZN(G378));
  INV_X1    g0923(.A(KEYINPUT57), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n854), .A2(KEYINPUT104), .A3(new_n855), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT104), .B1(new_n854), .B2(new_n855), .ZN(new_n1126));
  OAI211_X1 g0926(.A(G330), .B(new_n869), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n889), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n860), .A2(new_n889), .A3(G330), .A4(new_n869), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n304), .A2(new_n841), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT55), .Z(new_n1132));
  XNOR2_X1  g0932(.A(new_n317), .B(new_n1132), .ZN(new_n1133));
  XOR2_X1   g0933(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1134));
  XOR2_X1   g0934(.A(new_n1133), .B(new_n1134), .Z(new_n1135));
  AND3_X1   g0935(.A1(new_n1129), .A2(new_n1130), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1135), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1106), .B1(new_n1104), .B2(new_n1050), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1124), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1107), .B1(new_n1119), .B2(new_n1049), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1141), .B(KEYINPUT57), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1140), .A2(new_n664), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1135), .A2(new_n1052), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n757), .A2(new_n248), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G97), .B2(new_n763), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n512), .A2(G41), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1146), .B(new_n1147), .C1(new_n363), .C2(new_n743), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n768), .A2(new_n219), .B1(new_n808), .B2(new_n496), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n759), .A2(new_n217), .B1(new_n750), .B2(new_n772), .ZN(new_n1150));
  NOR4_X1   g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n948), .A4(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1147), .ZN(new_n1152));
  AOI21_X1  g0952(.A(G50), .B1(new_n268), .B2(new_n277), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1151), .A2(KEYINPUT58), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n816), .A2(new_n741), .B1(new_n743), .B2(new_n813), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT120), .Z(new_n1156));
  OAI22_X1  g0956(.A1(new_n768), .A2(new_n1059), .B1(new_n759), .B2(new_n1061), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n808), .A2(new_n1064), .B1(new_n298), .B2(new_n754), .ZN(new_n1158));
  NOR3_X1   g0958(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1160), .A2(KEYINPUT59), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n268), .B(new_n277), .C1(new_n757), .C2(new_n1055), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G124), .B2(new_n751), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT59), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1163), .B1(new_n1159), .B2(new_n1164), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1154), .B1(KEYINPUT58), .B2(new_n1151), .C1(new_n1161), .C2(new_n1165), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1166), .A2(new_n730), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n723), .B(new_n1167), .C1(new_n202), .C2(new_n795), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1144), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n1138), .B2(new_n718), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1143), .A2(new_n1171), .ZN(G375));
  OR3_X1    g0972(.A1(new_n1119), .A2(KEYINPUT122), .A3(new_n718), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n723), .B1(new_n211), .B2(new_n795), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n975), .B1(new_n768), .B2(new_n772), .C1(new_n773), .C2(new_n808), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n259), .B1(new_n803), .B2(G77), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1176), .B1(new_n219), .B2(new_n743), .C1(new_n496), .C2(new_n741), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n759), .A2(new_n473), .B1(new_n750), .B2(new_n589), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT123), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1175), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT124), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n768), .A2(new_n813), .B1(new_n202), .B2(new_n754), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G132), .B2(new_n746), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n759), .A2(new_n1055), .B1(new_n750), .B2(new_n1059), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n763), .B2(new_n1062), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n385), .B(new_n1145), .C1(G150), .C2(new_n797), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1183), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1181), .A2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1188), .A2(KEYINPUT125), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(KEYINPUT125), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n730), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n727), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1174), .B1(new_n1189), .B2(new_n1191), .C1(new_n886), .C2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(KEYINPUT122), .B1(new_n1119), .B2(new_n718), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1173), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n920), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1119), .A2(new_n1106), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1108), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1195), .A2(new_n1198), .ZN(G381));
  OR3_X1    g0999(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1200));
  NOR4_X1   g1000(.A1(G381), .A2(new_n1200), .A3(G387), .A4(G390), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1141), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n715), .B1(new_n1202), .B2(new_n1124), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1170), .B1(new_n1203), .B2(new_n1142), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n664), .B1(new_n1116), .B2(new_n1205), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1119), .A2(new_n1049), .A3(new_n1106), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1081), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1201), .A2(new_n1204), .A3(new_n1209), .ZN(G407));
  NAND2_X1  g1010(.A1(new_n647), .A2(G213), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1204), .A2(new_n1209), .A3(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(G407), .A2(G213), .A3(new_n1213), .ZN(G409));
  NAND3_X1  g1014(.A1(new_n1117), .A2(new_n1120), .A3(new_n664), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1141), .B(new_n1196), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1081), .B(new_n1215), .C1(new_n1217), .C2(new_n1170), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1081), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT117), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1215), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1219), .B1(new_n1221), .B2(new_n1121), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1218), .B1(G375), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT60), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1197), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1119), .A2(KEYINPUT60), .A3(new_n1106), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1225), .A2(new_n664), .A3(new_n1108), .A4(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(G384), .A2(KEYINPUT126), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  AND3_X1   g1029(.A1(new_n1195), .A2(new_n1227), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(G384), .A2(KEYINPUT126), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1195), .A2(new_n1227), .B1(new_n1231), .B2(new_n1229), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1223), .A2(new_n1211), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(KEYINPUT62), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT61), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G2897), .B(new_n1212), .C1(new_n1230), .C2(new_n1232), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1195), .A2(new_n1227), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1195), .A2(new_n1227), .A3(new_n1229), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1212), .A2(G2897), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1208), .B1(new_n1171), .B2(new_n1216), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G378), .B2(new_n1204), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1237), .B(new_n1243), .C1(new_n1245), .C2(new_n1212), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT62), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1223), .A2(new_n1247), .A3(new_n1233), .A4(new_n1211), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1235), .A2(new_n1236), .A3(new_n1246), .A4(new_n1248), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(G393), .B(G396), .ZN(new_n1250));
  INV_X1    g1050(.A(G390), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(G387), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n943), .A2(G390), .A3(new_n969), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1250), .B1(new_n1254), .B2(KEYINPUT127), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n943), .A2(G390), .A3(new_n969), .ZN(new_n1256));
  AOI21_X1  g1056(.A(G390), .B1(new_n943), .B2(new_n969), .ZN(new_n1257));
  OAI211_X1 g1057(.A(KEYINPUT127), .B(new_n1250), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1255), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1249), .A2(new_n1261), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1242), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1223), .A2(new_n1211), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT61), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1223), .A2(KEYINPUT63), .A3(new_n1211), .A4(new_n1233), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT63), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1234), .A2(new_n1269), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1267), .A2(new_n1268), .A3(new_n1270), .A4(new_n1260), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1262), .A2(new_n1271), .ZN(G405));
  OAI21_X1  g1072(.A(new_n1233), .B1(new_n1255), .B2(new_n1259), .ZN(new_n1273));
  OAI21_X1  g1073(.A(KEYINPUT127), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1250), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1276), .B(new_n1258), .C1(new_n1232), .C2(new_n1230), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1273), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G378), .A2(new_n1204), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G375), .A2(new_n1209), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1278), .A2(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1273), .A2(new_n1277), .A3(new_n1279), .A4(new_n1280), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(G402));
endmodule


