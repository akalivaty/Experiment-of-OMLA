//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1214, new_n1215, new_n1216, new_n1217, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289, new_n1290;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(KEYINPUT65), .ZN(new_n210));
  XNOR2_X1  g0010(.A(KEYINPUT64), .B(G244), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G77), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G68), .A2(G238), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  NAND4_X1  g0014(.A1(new_n210), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n209), .A2(KEYINPUT65), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n206), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n206), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(G250), .B1(G257), .B2(G264), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n201), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  OAI22_X1  g0029(.A1(new_n223), .A2(KEYINPUT0), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT0), .B2(new_n223), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n218), .A2(new_n219), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT66), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT76), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G13), .A3(G20), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n256), .A2(new_n224), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G1), .B2(new_n225), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n255), .B1(new_n251), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT73), .ZN(new_n261));
  OR2_X1    g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(new_n225), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT7), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(KEYINPUT7), .B1(new_n269), .B2(new_n225), .ZN(new_n270));
  OAI21_X1  g0070(.A(G68), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT16), .ZN(new_n272));
  INV_X1    g0072(.A(G58), .ZN(new_n273));
  INV_X1    g0073(.A(G68), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(G20), .B1(new_n275), .B2(new_n201), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G159), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n276), .A2(KEYINPUT72), .A3(new_n278), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n271), .A2(new_n272), .A3(new_n280), .A4(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n272), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n264), .A2(new_n265), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n269), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n274), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n283), .B1(new_n286), .B2(new_n279), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n256), .A2(new_n224), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n261), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI211_X1 g0090(.A(KEYINPUT73), .B(new_n257), .C1(new_n282), .C2(new_n287), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n260), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G190), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G41), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n294), .A2(G1), .A3(G13), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(G232), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G41), .ZN(new_n298));
  INV_X1    g0098(.A(G45), .ZN(new_n299));
  AOI21_X1  g0099(.A(G1), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G274), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n295), .ZN(new_n303));
  INV_X1    g0103(.A(G1698), .ZN(new_n304));
  OAI211_X1 g0104(.A(G223), .B(new_n304), .C1(new_n267), .C2(new_n268), .ZN(new_n305));
  OAI211_X1 g0105(.A(G226), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G33), .A2(G87), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AOI211_X1 g0108(.A(new_n293), .B(new_n302), .C1(new_n303), .C2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G200), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n303), .ZN(new_n311));
  INV_X1    g0111(.A(new_n302), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT74), .B1(new_n309), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n302), .B1(new_n308), .B2(new_n303), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G190), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT74), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n316), .B(new_n317), .C1(new_n310), .C2(new_n315), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT17), .B1(new_n292), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT75), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI211_X1 g0122(.A(KEYINPUT75), .B(KEYINPUT17), .C1(new_n292), .C2(new_n319), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT17), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n314), .A2(new_n318), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n325), .B(new_n260), .C1(new_n291), .C2(new_n290), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n322), .A2(new_n323), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n315), .A2(G169), .ZN(new_n329));
  INV_X1    g0129(.A(G179), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n329), .B1(new_n330), .B2(new_n315), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n292), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT18), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT18), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n292), .A2(new_n334), .A3(new_n331), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n249), .B1(new_n328), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n327), .A2(new_n324), .ZN(new_n338));
  INV_X1    g0138(.A(new_n323), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT75), .B1(new_n326), .B2(KEYINPUT17), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n336), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(KEYINPUT76), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n262), .A2(new_n263), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(G223), .A3(G1698), .ZN(new_n345));
  INV_X1    g0145(.A(G77), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n304), .ZN(new_n347));
  INV_X1    g0147(.A(G222), .ZN(new_n348));
  OAI221_X1 g0148(.A(new_n345), .B1(new_n346), .B2(new_n344), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n303), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n303), .A2(new_n300), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G226), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n350), .A2(new_n301), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G200), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT68), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n353), .A2(KEYINPUT68), .A3(G200), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n258), .A2(G50), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(G50), .B2(new_n254), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n277), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n225), .A2(G33), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n361), .B1(new_n250), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n289), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT9), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n350), .A2(G190), .A3(new_n301), .A4(new_n352), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n358), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT69), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n366), .A2(new_n370), .A3(new_n367), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT10), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n372), .B(new_n371), .C1(new_n358), .C2(new_n368), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n353), .A2(G169), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(new_n330), .B2(new_n353), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n365), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT15), .B(G87), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(new_n362), .ZN(new_n380));
  INV_X1    g0180(.A(new_n277), .ZN(new_n381));
  OAI22_X1  g0181(.A1(new_n250), .A2(new_n381), .B1(new_n225), .B2(new_n346), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n380), .B1(new_n382), .B2(KEYINPUT67), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(KEYINPUT67), .B2(new_n382), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n289), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n258), .A2(G77), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(G77), .B2(new_n254), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n344), .A2(G238), .A3(G1698), .ZN(new_n388));
  INV_X1    g0188(.A(G107), .ZN(new_n389));
  INV_X1    g0189(.A(G232), .ZN(new_n390));
  OAI221_X1 g0190(.A(new_n388), .B1(new_n389), .B2(new_n344), .C1(new_n347), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n303), .ZN(new_n392));
  INV_X1    g0192(.A(new_n301), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n351), .B2(new_n211), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n395), .A2(G190), .ZN(new_n396));
  AOI21_X1  g0196(.A(G200), .B1(new_n392), .B2(new_n394), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n385), .B(new_n387), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n385), .A2(new_n387), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n395), .A2(new_n330), .ZN(new_n400));
  INV_X1    g0200(.A(G169), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n401), .B1(new_n392), .B2(new_n394), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n399), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n374), .A2(new_n375), .A3(new_n378), .A4(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT12), .ZN(new_n406));
  INV_X1    g0206(.A(G13), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n407), .A2(G1), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n274), .A2(G20), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n406), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n408), .A2(KEYINPUT12), .A3(G20), .A4(new_n274), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n411), .B(new_n412), .C1(new_n258), .C2(new_n274), .ZN(new_n413));
  XOR2_X1   g0213(.A(new_n413), .B(KEYINPUT70), .Z(new_n414));
  OAI221_X1 g0214(.A(new_n410), .B1(new_n362), .B2(new_n346), .C1(new_n381), .C2(new_n202), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n289), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT11), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n344), .A2(G232), .A3(G1698), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G97), .ZN(new_n421));
  INV_X1    g0221(.A(G226), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n420), .B(new_n421), .C1(new_n347), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n303), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT13), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n393), .B1(new_n351), .B2(G238), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n425), .B1(new_n424), .B2(new_n426), .ZN(new_n428));
  OAI21_X1  g0228(.A(G169), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(KEYINPUT71), .A2(KEYINPUT14), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n427), .A2(new_n428), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n429), .A2(new_n431), .B1(new_n432), .B2(G179), .ZN(new_n433));
  OR2_X1    g0233(.A1(new_n429), .A2(new_n431), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n419), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n432), .A2(new_n293), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n310), .B1(new_n427), .B2(new_n428), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n418), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n405), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n337), .A2(new_n343), .A3(new_n439), .ZN(new_n440));
  OAI211_X1 g0240(.A(G250), .B(new_n304), .C1(new_n267), .C2(new_n268), .ZN(new_n441));
  OAI211_X1 g0241(.A(G257), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G294), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n303), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n299), .A2(G1), .ZN(new_n446));
  NOR2_X1   g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  AND2_X1   g0247(.A1(KEYINPUT5), .A2(G41), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n446), .B(G274), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT77), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g0251(.A(KEYINPUT5), .B(G41), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n452), .A2(KEYINPUT77), .A3(G274), .A4(new_n446), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n224), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n452), .A2(new_n446), .B1(new_n455), .B2(new_n294), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G264), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n445), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n310), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n444), .A2(new_n303), .B1(new_n456), .B2(G264), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(new_n293), .A3(new_n454), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT22), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(KEYINPUT83), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(KEYINPUT83), .ZN(new_n466));
  AOI21_X1  g0266(.A(G20), .B1(new_n262), .B2(new_n263), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n466), .B1(new_n467), .B2(G87), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n225), .B(G87), .C1(new_n267), .C2(new_n268), .ZN(new_n469));
  INV_X1    g0269(.A(new_n466), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n465), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  OR3_X1    g0272(.A1(new_n225), .A2(KEYINPUT23), .A3(G107), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n225), .A2(G33), .A3(G116), .ZN(new_n474));
  OAI21_X1  g0274(.A(KEYINPUT23), .B1(new_n225), .B2(G107), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n472), .A2(KEYINPUT24), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT24), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n469), .A2(new_n470), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n344), .A2(new_n225), .A3(G87), .A4(new_n466), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n464), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n479), .B1(new_n482), .B2(new_n476), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n478), .A2(new_n483), .A3(new_n289), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n408), .A2(G20), .A3(new_n389), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n485), .B(KEYINPUT25), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n252), .A2(G33), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n257), .A2(new_n253), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n486), .B1(G107), .B2(new_n489), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n462), .A2(new_n484), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n460), .A2(G179), .A3(new_n454), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n458), .A2(G169), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n484), .A2(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT84), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n484), .A2(new_n490), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(new_n492), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT84), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n462), .A2(new_n484), .A3(new_n490), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT21), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT20), .ZN(new_n504));
  INV_X1    g0304(.A(G116), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n225), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G283), .ZN(new_n507));
  INV_X1    g0307(.A(G97), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(G33), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n506), .B1(new_n509), .B2(new_n225), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n504), .B1(new_n510), .B2(new_n257), .ZN(new_n511));
  INV_X1    g0311(.A(G33), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G97), .ZN(new_n513));
  AOI21_X1  g0313(.A(G20), .B1(new_n513), .B2(new_n507), .ZN(new_n514));
  OAI211_X1 g0314(.A(KEYINPUT20), .B(new_n289), .C1(new_n514), .C2(new_n506), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n488), .A2(G116), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n253), .A2(new_n505), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(G264), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n521));
  OAI211_X1 g0321(.A(G257), .B(new_n304), .C1(new_n267), .C2(new_n268), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n262), .A2(G303), .A3(new_n263), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n303), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n456), .A2(G270), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(new_n454), .A3(new_n526), .ZN(new_n527));
  AND4_X1   g0327(.A1(KEYINPUT82), .A2(new_n520), .A3(G169), .A4(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n401), .B1(new_n516), .B2(new_n519), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT82), .B1(new_n529), .B2(new_n527), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n503), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n520), .A2(KEYINPUT21), .A3(new_n527), .A4(G169), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT81), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT81), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n529), .A2(new_n534), .A3(KEYINPUT21), .A4(new_n527), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  OR2_X1    g0336(.A1(new_n527), .A2(new_n330), .ZN(new_n537));
  INV_X1    g0337(.A(new_n520), .ZN(new_n538));
  OR2_X1    g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n527), .A2(new_n310), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n527), .A2(G190), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AND4_X1   g0342(.A1(new_n531), .A2(new_n536), .A3(new_n539), .A4(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n225), .ZN(new_n545));
  NOR2_X1   g0345(.A1(G87), .A2(G97), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n389), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n547), .A3(KEYINPUT79), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n225), .B(G68), .C1(new_n267), .C2(new_n268), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT19), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(new_n421), .B2(G20), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT79), .B1(new_n545), .B2(new_n547), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n289), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n379), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(new_n253), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n489), .A2(new_n555), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n554), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(G250), .B1(new_n299), .B2(G1), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n252), .A2(G45), .A3(G274), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n560), .A2(new_n561), .B1(new_n455), .B2(new_n294), .ZN(new_n562));
  OAI211_X1 g0362(.A(G238), .B(new_n304), .C1(new_n267), .C2(new_n268), .ZN(new_n563));
  OAI211_X1 g0363(.A(G244), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G33), .A2(G116), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n562), .B1(new_n566), .B2(new_n303), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n567), .A2(KEYINPUT78), .A3(new_n330), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n559), .A2(new_n568), .ZN(new_n569));
  AOI211_X1 g0369(.A(G179), .B(new_n562), .C1(new_n566), .C2(new_n303), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT78), .B1(new_n567), .B2(G169), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n567), .A2(new_n293), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(G200), .B2(new_n567), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n489), .A2(G87), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n554), .A2(new_n557), .A3(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n569), .A2(new_n573), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n254), .A2(G97), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n488), .B2(G97), .ZN(new_n580));
  XNOR2_X1  g0380(.A(G97), .B(G107), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT6), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n582), .A2(new_n508), .A3(G107), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n586), .A2(G20), .B1(G77), .B2(new_n277), .ZN(new_n587));
  OAI21_X1  g0387(.A(G107), .B1(new_n266), .B2(new_n270), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n580), .B1(new_n589), .B2(new_n289), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT4), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n591), .A2(G1698), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n592), .B(G244), .C1(new_n268), .C2(new_n267), .ZN(new_n593));
  INV_X1    g0393(.A(G244), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n262), .B2(new_n263), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n593), .B(new_n507), .C1(new_n595), .C2(KEYINPUT4), .ZN(new_n596));
  OAI21_X1  g0396(.A(G250), .B1(new_n267), .B2(new_n268), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n304), .B1(new_n597), .B2(KEYINPUT4), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n303), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n451), .A2(new_n453), .B1(new_n456), .B2(G257), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n599), .A2(new_n293), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(G200), .B1(new_n599), .B2(new_n600), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n590), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n584), .B1(new_n582), .B2(new_n581), .ZN(new_n604));
  OAI22_X1  g0404(.A1(new_n604), .A2(new_n225), .B1(new_n346), .B2(new_n381), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n389), .B1(new_n284), .B2(new_n285), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n289), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n580), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n599), .A2(G179), .A3(new_n600), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n401), .B1(new_n599), .B2(new_n600), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n578), .A2(KEYINPUT80), .A3(new_n603), .A4(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT80), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n603), .A2(new_n612), .ZN(new_n615));
  INV_X1    g0415(.A(new_n553), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n616), .A2(new_n548), .A3(new_n549), .A4(new_n551), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n556), .B1(new_n617), .B2(new_n289), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n567), .A2(new_n293), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n567), .A2(G200), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n618), .B(new_n576), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n566), .A2(new_n303), .ZN(new_n622));
  INV_X1    g0422(.A(new_n562), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n401), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n570), .B1(new_n625), .B2(KEYINPUT78), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n559), .A2(new_n568), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n621), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n614), .B1(new_n615), .B2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n502), .A2(new_n543), .A3(new_n613), .A4(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n440), .A2(new_n630), .ZN(G372));
  INV_X1    g0431(.A(new_n440), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  INV_X1    g0433(.A(new_n612), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n633), .B1(new_n578), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n571), .A2(new_n559), .A3(new_n625), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n621), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n634), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n635), .B1(new_n639), .B2(new_n633), .ZN(new_n640));
  INV_X1    g0440(.A(new_n636), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n531), .A2(new_n498), .A3(new_n536), .A4(new_n539), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n500), .A2(new_n603), .A3(new_n612), .A4(new_n621), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n632), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n374), .A2(new_n375), .ZN(new_n647));
  INV_X1    g0447(.A(new_n438), .ZN(new_n648));
  INV_X1    g0448(.A(new_n403), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n648), .B1(new_n435), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n328), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT85), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n292), .A2(new_n334), .A3(new_n331), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n334), .B1(new_n292), .B2(new_n331), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n333), .A2(KEYINPUT85), .A3(new_n335), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n647), .B1(new_n651), .B2(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n658), .A2(new_n378), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n646), .A2(new_n659), .ZN(G369));
  NAND3_X1  g0460(.A1(new_n531), .A2(new_n536), .A3(new_n539), .ZN(new_n661));
  OR3_X1    g0461(.A1(new_n409), .A2(KEYINPUT27), .A3(G20), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT27), .B1(new_n409), .B2(G20), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n520), .A2(new_n666), .ZN(new_n667));
  MUX2_X1   g0467(.A(new_n661), .B(new_n543), .S(new_n667), .Z(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(G330), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n496), .A2(new_n666), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n502), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n494), .A2(new_n666), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n666), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n661), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT86), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n494), .A2(new_n677), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n676), .A2(new_n680), .A3(new_n681), .ZN(G399));
  NOR2_X1   g0482(.A1(new_n221), .A2(G41), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n546), .A2(new_n389), .A3(new_n505), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n684), .A2(G1), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n229), .B2(new_n684), .ZN(new_n688));
  XOR2_X1   g0488(.A(new_n688), .B(KEYINPUT28), .Z(new_n689));
  NAND2_X1  g0489(.A1(new_n645), .A2(new_n677), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT29), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n633), .B1(new_n628), .B2(new_n612), .ZN(new_n693));
  OAI22_X1  g0493(.A1(new_n693), .A2(KEYINPUT88), .B1(new_n638), .B2(new_n633), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n693), .A2(KEYINPUT88), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n644), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n696), .A2(KEYINPUT29), .A3(new_n677), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(G330), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT31), .B1(new_n630), .B2(new_n666), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n599), .A2(new_n600), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(new_n454), .B2(new_n460), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n527), .A2(new_n330), .A3(new_n624), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n460), .A2(new_n567), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n537), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n701), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n704), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT87), .ZN(new_n710));
  AOI211_X1 g0510(.A(new_n710), .B(KEYINPUT30), .C1(new_n706), .C2(new_n701), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n707), .A2(new_n708), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n710), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n677), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n700), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  INV_X1    g0518(.A(new_n709), .ZN(new_n719));
  AOI211_X1 g0519(.A(new_n718), .B(new_n677), .C1(new_n719), .C2(new_n713), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n699), .B1(new_n717), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n698), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n689), .B1(new_n724), .B2(new_n252), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT89), .ZN(G364));
  AOI21_X1  g0526(.A(new_n224), .B1(G20), .B2(new_n401), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n330), .A2(new_n310), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n225), .A2(new_n293), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n225), .A2(G190), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n730), .A2(new_n202), .B1(new_n732), .B2(new_n274), .ZN(new_n733));
  INV_X1    g0533(.A(new_n731), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n734), .A2(new_n330), .A3(G200), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n344), .B1(new_n736), .B2(new_n346), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G179), .A2(G200), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n225), .B1(new_n738), .B2(G190), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI211_X1 g0540(.A(new_n733), .B(new_n737), .C1(G97), .C2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n731), .A2(new_n738), .ZN(new_n742));
  INV_X1    g0542(.A(G159), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT32), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n310), .A2(G179), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n731), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G107), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n729), .A2(G179), .A3(new_n310), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n729), .A2(new_n746), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n751), .A2(G58), .B1(new_n753), .B2(G87), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n741), .A2(new_n745), .A3(new_n749), .A4(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(KEYINPUT92), .ZN(new_n757));
  INV_X1    g0557(.A(new_n732), .ZN(new_n758));
  XNOR2_X1  g0558(.A(KEYINPUT33), .B(G317), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n751), .A2(G322), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT93), .ZN(new_n761));
  AOI22_X1  g0561(.A1(G303), .A2(new_n753), .B1(new_n748), .B2(G283), .ZN(new_n762));
  INV_X1    g0562(.A(new_n742), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n735), .A2(G311), .B1(G329), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G326), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n269), .B1(new_n730), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(G294), .B2(new_n740), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n761), .A2(new_n762), .A3(new_n764), .A4(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT92), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n768), .B1(new_n755), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n727), .B1(new_n757), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n407), .A2(G20), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G45), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n684), .A2(G1), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n221), .A2(new_n269), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n775), .A2(G355), .B1(new_n505), .B2(new_n221), .ZN(new_n776));
  AOI21_X1  g0576(.A(G45), .B1(new_n228), .B2(G50), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(new_n244), .B2(G45), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n221), .A2(new_n344), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n776), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G13), .A2(G33), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n225), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT91), .Z(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n727), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n774), .B1(new_n781), .B2(new_n786), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n771), .B(new_n787), .C1(new_n668), .C2(new_n784), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT94), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n668), .A2(G330), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(KEYINPUT90), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n669), .A2(KEYINPUT90), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n774), .B(new_n791), .C1(new_n792), .C2(new_n790), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n789), .A2(new_n793), .ZN(G396));
  INV_X1    g0594(.A(new_n774), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n727), .A2(new_n782), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n795), .B1(G77), .B2(new_n797), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n736), .A2(new_n505), .B1(new_n389), .B2(new_n752), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n344), .B(new_n799), .C1(G311), .C2(new_n763), .ZN(new_n800));
  INV_X1    g0600(.A(G294), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n750), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G303), .ZN(new_n803));
  INV_X1    g0603(.A(G283), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n730), .A2(new_n803), .B1(new_n732), .B2(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n802), .B(new_n805), .C1(G87), .C2(new_n748), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n800), .B(new_n806), .C1(new_n508), .C2(new_n739), .ZN(new_n807));
  INV_X1    g0607(.A(G137), .ZN(new_n808));
  INV_X1    g0608(.A(G150), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n730), .A2(new_n808), .B1(new_n732), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT95), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n735), .A2(G159), .B1(new_n751), .B2(G143), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT34), .Z(new_n814));
  AOI21_X1  g0614(.A(new_n269), .B1(new_n753), .B2(G50), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n763), .A2(G132), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n748), .A2(G68), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n740), .A2(G58), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n815), .A2(new_n816), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n807), .B1(new_n814), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n798), .B1(new_n820), .B2(new_n727), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n399), .A2(new_n666), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n398), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n403), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n403), .A2(new_n666), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n782), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n821), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT96), .Z(new_n831));
  NAND2_X1  g0631(.A1(new_n690), .A2(new_n827), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n645), .A2(new_n677), .A3(new_n828), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(new_n722), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n795), .B1(new_n834), .B2(new_n722), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n831), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G384));
  NOR2_X1   g0639(.A1(new_n772), .A2(new_n252), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n286), .A2(new_n279), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT16), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n260), .B1(new_n842), .B2(new_n257), .ZN(new_n843));
  INV_X1    g0643(.A(new_n664), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n331), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n326), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(KEYINPUT37), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n664), .B(KEYINPUT97), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n292), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n332), .A2(new_n849), .A3(new_n850), .A4(new_n326), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n322), .A2(new_n323), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n336), .B1(new_n853), .B2(new_n338), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n843), .A2(new_n844), .ZN(new_n855));
  OAI211_X1 g0655(.A(KEYINPUT38), .B(new_n852), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(KEYINPUT98), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n844), .B(new_n843), .C1(new_n328), .C2(new_n336), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT98), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n858), .A2(new_n859), .A3(KEYINPUT38), .A4(new_n852), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n855), .B1(new_n341), .B2(new_n342), .ZN(new_n862));
  INV_X1    g0662(.A(new_n852), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n857), .A2(new_n860), .A3(new_n864), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n718), .B(new_n677), .C1(new_n712), .C2(new_n714), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n827), .B1(new_n717), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n435), .A2(new_n438), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n418), .A2(new_n666), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n869), .B(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT40), .B1(new_n865), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n849), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n657), .B2(new_n328), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n332), .A2(new_n849), .A3(new_n326), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT37), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n851), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT38), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n862), .A2(new_n861), .A3(new_n863), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT40), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n882), .A2(new_n872), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n874), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n717), .A2(new_n867), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n632), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n884), .B(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(G330), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n888), .B(KEYINPUT100), .Z(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n848), .B1(new_n655), .B2(new_n656), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n833), .A2(new_n826), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n871), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n891), .B1(new_n865), .B2(new_n894), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n857), .A2(KEYINPUT39), .A3(new_n860), .A4(new_n864), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n435), .A2(new_n677), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT99), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT39), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n880), .B2(new_n881), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n896), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n692), .A2(new_n697), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n378), .B(new_n658), .C1(new_n440), .C2(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n903), .B(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n840), .B1(new_n890), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n890), .B2(new_n906), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n229), .A2(new_n346), .A3(new_n275), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n274), .A2(G50), .ZN(new_n910));
  OAI211_X1 g0710(.A(G1), .B(new_n407), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(G116), .B(new_n226), .C1(new_n586), .C2(KEYINPUT35), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(KEYINPUT35), .B2(new_n586), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n913), .B(KEYINPUT36), .Z(new_n914));
  NAND3_X1  g0714(.A1(new_n908), .A2(new_n911), .A3(new_n914), .ZN(G367));
  AOI21_X1  g0715(.A(new_n615), .B1(new_n609), .B2(new_n666), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n916), .B(KEYINPUT102), .Z(new_n917));
  NAND2_X1  g0717(.A1(new_n634), .A2(new_n666), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  OR3_X1    g0720(.A1(new_n680), .A2(new_n920), .A3(KEYINPUT42), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT42), .B1(new_n680), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n612), .B1(new_n917), .B2(new_n498), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n677), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n921), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT43), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n577), .A2(new_n677), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n637), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n927), .A2(new_n636), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n925), .B1(new_n926), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n675), .A2(new_n919), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n926), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT101), .Z(new_n935));
  XNOR2_X1  g0735(.A(new_n933), .B(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n932), .B(new_n936), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n683), .B(KEYINPUT41), .Z(new_n938));
  NAND2_X1  g0738(.A1(new_n680), .A2(new_n681), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(new_n920), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT45), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n920), .ZN(new_n942));
  XNOR2_X1  g0742(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n941), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n675), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n941), .A2(new_n676), .A3(new_n944), .A4(new_n945), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n674), .B(new_n679), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT104), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n669), .A2(new_n950), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n949), .B(new_n951), .Z(new_n952));
  NOR2_X1   g0752(.A1(new_n952), .A2(new_n724), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n947), .A2(new_n948), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n938), .B1(new_n954), .B2(new_n723), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n773), .A2(G1), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n937), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n240), .A2(new_n780), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n786), .B1(new_n220), .B2(new_n379), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n736), .A2(new_n202), .B1(new_n747), .B2(new_n346), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n269), .B(new_n960), .C1(G137), .C2(new_n763), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n751), .A2(G150), .B1(new_n758), .B2(G159), .ZN(new_n962));
  INV_X1    g0762(.A(new_n730), .ZN(new_n963));
  AOI22_X1  g0763(.A1(G143), .A2(new_n963), .B1(new_n753), .B2(G58), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n739), .A2(new_n274), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n961), .A2(new_n962), .A3(new_n964), .A4(new_n966), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n736), .A2(new_n804), .B1(new_n801), .B2(new_n732), .ZN(new_n968));
  XOR2_X1   g0768(.A(KEYINPUT105), .B(G311), .Z(new_n969));
  OAI22_X1  g0769(.A1(new_n730), .A2(new_n969), .B1(new_n750), .B2(new_n803), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(KEYINPUT106), .B1(new_n752), .B2(new_n505), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT46), .Z(new_n973));
  OAI211_X1 g0773(.A(new_n971), .B(new_n973), .C1(new_n389), .C2(new_n739), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n747), .A2(new_n508), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n344), .B(new_n975), .C1(G317), .C2(new_n763), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT107), .Z(new_n977));
  OAI21_X1  g0777(.A(new_n967), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT47), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n727), .B1(new_n978), .B2(new_n979), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n795), .B1(new_n958), .B2(new_n959), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT108), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n784), .B2(new_n930), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n957), .A2(new_n984), .ZN(G387));
  NOR2_X1   g0785(.A1(new_n953), .A2(new_n684), .ZN(new_n986));
  INV_X1    g0786(.A(new_n952), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n986), .B1(new_n723), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n251), .A2(new_n202), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT50), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n686), .B(new_n299), .C1(new_n274), .C2(new_n346), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n779), .B1(new_n990), .B2(new_n991), .C1(new_n237), .C2(new_n299), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n775), .A2(new_n685), .B1(new_n389), .B2(new_n221), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n774), .B1(new_n994), .B2(new_n786), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n344), .B1(new_n748), .B2(G116), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n752), .A2(new_n801), .B1(new_n739), .B2(new_n804), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n969), .A2(new_n732), .ZN(new_n998));
  INV_X1    g0798(.A(G322), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n736), .A2(new_n803), .B1(new_n999), .B2(new_n730), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n998), .B(new_n1000), .C1(G317), .C2(new_n751), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n997), .B1(new_n1001), .B2(KEYINPUT48), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(KEYINPUT48), .B2(new_n1001), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT49), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n996), .B1(new_n765), .B2(new_n742), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n1004), .B2(new_n1003), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n735), .A2(G68), .B1(new_n758), .B2(new_n251), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT109), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G77), .A2(new_n753), .B1(new_n763), .B2(G150), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n202), .B2(new_n750), .C1(new_n743), .C2(new_n730), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n739), .A2(new_n379), .ZN(new_n1011));
  NOR4_X1   g0811(.A1(new_n1010), .A2(new_n269), .A3(new_n975), .A4(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1006), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n727), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n995), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n674), .B2(new_n785), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(new_n987), .B2(new_n956), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n988), .A2(new_n1017), .ZN(G393));
  AND2_X1   g0818(.A1(new_n954), .A2(new_n683), .ZN(new_n1019));
  AND2_X1   g0819(.A1(new_n947), .A2(new_n948), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1019), .B1(new_n1020), .B2(new_n953), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n956), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n786), .B1(new_n508), .B2(new_n220), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n247), .A2(new_n780), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n795), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n750), .A2(new_n743), .B1(new_n730), .B2(new_n809), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT51), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G50), .A2(new_n758), .B1(new_n763), .B2(G143), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n735), .A2(new_n251), .B1(new_n753), .B2(G68), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n739), .A2(new_n346), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n269), .B(new_n1030), .C1(G87), .C2(new_n748), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n752), .A2(new_n804), .B1(new_n742), .B2(new_n999), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT110), .Z(new_n1034));
  AOI22_X1  g0834(.A1(new_n735), .A2(G294), .B1(new_n758), .B2(G303), .ZN(new_n1035));
  AND3_X1   g0835(.A1(new_n1035), .A2(new_n269), .A3(new_n749), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1034), .B(new_n1036), .C1(new_n505), .C2(new_n739), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n751), .A2(G311), .B1(new_n963), .B2(G317), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT52), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1032), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1025), .B1(new_n1040), .B2(new_n727), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n919), .B2(new_n784), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1021), .A2(new_n1022), .A3(new_n1042), .ZN(G390));
  XNOR2_X1  g0843(.A(KEYINPUT54), .B(G143), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n735), .A2(new_n1045), .B1(new_n758), .B2(G137), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT117), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n269), .B1(new_n963), .B2(G128), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n743), .B2(new_n739), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n751), .A2(G132), .B1(new_n748), .B2(G50), .ZN(new_n1050));
  INV_X1    g0850(.A(G125), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1050), .B1(new_n1051), .B2(new_n742), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT53), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n752), .B2(new_n809), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n753), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1049), .B(new_n1052), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n730), .A2(new_n804), .B1(new_n742), .B2(new_n801), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n344), .B1(new_n753), .B2(G87), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1058), .B(new_n817), .C1(new_n736), .C2(new_n508), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1057), .B(new_n1059), .C1(G107), .C2(new_n758), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1030), .B1(G116), .B2(new_n751), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT118), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1047), .A2(new_n1056), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n795), .B1(new_n251), .B2(new_n797), .C1(new_n1063), .C2(new_n1014), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n896), .A2(new_n901), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1064), .B1(new_n1065), .B2(new_n782), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n896), .A2(new_n901), .B1(new_n898), .B2(new_n893), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT113), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n629), .A2(new_n613), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1069), .A2(new_n543), .A3(new_n502), .A4(new_n677), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n715), .B1(new_n1070), .B2(KEYINPUT31), .ZN(new_n1071));
  OAI211_X1 g0871(.A(G330), .B(new_n828), .C1(new_n1071), .C2(new_n720), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n871), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1068), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n722), .A2(KEYINPUT113), .A3(new_n828), .A4(new_n871), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  AND3_X1   g0877(.A1(new_n696), .A2(new_n677), .A3(new_n824), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n871), .B1(new_n1078), .B2(new_n825), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n898), .B(new_n1079), .C1(new_n880), .C2(new_n881), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n1067), .A2(new_n1077), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT112), .ZN(new_n1083));
  OAI211_X1 g0883(.A(G330), .B(new_n828), .C1(new_n1071), .C2(new_n866), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1083), .B1(new_n1084), .B2(new_n1073), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n868), .A2(KEYINPUT112), .A3(G330), .A4(new_n871), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n893), .A2(new_n898), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1081), .B1(new_n1065), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1088), .B1(new_n1090), .B2(KEYINPUT111), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT111), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n1067), .B2(new_n1081), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1082), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1066), .B1(new_n1094), .B2(new_n956), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT115), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1085), .A2(new_n1086), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n892), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n825), .B(new_n1078), .C1(new_n1084), .C2(new_n1073), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1076), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n866), .B1(new_n700), .B2(new_n716), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n440), .A2(new_n1103), .A3(new_n699), .ZN(new_n1104));
  OAI21_X1  g0904(.A(KEYINPUT114), .B1(new_n905), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n632), .A2(new_n698), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n647), .A2(new_n869), .A3(new_n378), .A4(new_n404), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n341), .A2(new_n342), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1107), .B1(new_n249), .B2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1109), .A2(new_n885), .A3(G330), .A4(new_n343), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT114), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1106), .A2(new_n1110), .A3(new_n659), .A4(new_n1111), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n1105), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1096), .B1(new_n1102), .B2(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1098), .A2(new_n892), .B1(new_n1076), .B2(new_n1100), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1105), .A2(new_n1112), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n1115), .A2(KEYINPUT115), .A3(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(KEYINPUT116), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(KEYINPUT115), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1102), .A2(new_n1096), .A3(new_n1113), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT116), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1094), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1065), .A2(new_n1089), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1125), .A2(KEYINPUT111), .A3(new_n1080), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1126), .A2(new_n1093), .A3(new_n1087), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1082), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n683), .B1(new_n1124), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1095), .B1(new_n1123), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(KEYINPUT119), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT119), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1133), .B(new_n1095), .C1(new_n1123), .C2(new_n1130), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1132), .A2(new_n1134), .ZN(G378));
  INV_X1    g0935(.A(G132), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n730), .A2(new_n1051), .B1(new_n732), .B2(new_n1136), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n751), .A2(G128), .B1(new_n753), .B2(new_n1045), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n808), .B2(new_n736), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1137), .B(new_n1139), .C1(G150), .C2(new_n740), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1141), .A2(KEYINPUT59), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(KEYINPUT59), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n512), .B(new_n298), .C1(new_n747), .C2(new_n743), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(G124), .B2(new_n763), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1142), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n736), .A2(new_n379), .B1(new_n508), .B2(new_n732), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n298), .B(new_n269), .C1(new_n752), .C2(new_n346), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n1147), .A2(new_n965), .A3(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n747), .A2(new_n273), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT120), .Z(new_n1151));
  NAND2_X1  g0951(.A1(new_n963), .A2(G116), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n751), .A2(G107), .B1(new_n763), .B2(G283), .ZN(new_n1153));
  AND4_X1   g0953(.A1(new_n1149), .A2(new_n1151), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(KEYINPUT58), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1154), .A2(KEYINPUT58), .ZN(new_n1156));
  AOI21_X1  g0956(.A(G50), .B1(new_n512), .B2(new_n298), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n344), .B2(G41), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1146), .A2(new_n1155), .A3(new_n1156), .A4(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n727), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n774), .B1(new_n202), .B2(new_n796), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n647), .A2(new_n378), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n365), .A2(new_n844), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1162), .B(new_n1163), .ZN(new_n1164));
  XOR2_X1   g0964(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1165));
  XNOR2_X1  g0965(.A(new_n1164), .B(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1160), .B(new_n1161), .C1(new_n1167), .C2(new_n829), .ZN(new_n1168));
  OR3_X1    g0968(.A1(new_n874), .A2(new_n883), .A3(new_n699), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n903), .A2(new_n1167), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n895), .A2(new_n902), .A3(new_n1166), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n874), .A2(new_n883), .A3(new_n699), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n895), .A2(new_n902), .A3(new_n1166), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1166), .B1(new_n895), .B2(new_n902), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1172), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n956), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1168), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1113), .B1(new_n1124), .B2(new_n1129), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1177), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT57), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1116), .B1(new_n1094), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(KEYINPUT57), .B1(new_n1185), .B2(new_n1177), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1179), .B1(new_n1187), .B2(new_n683), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(G375));
  OAI21_X1  g0989(.A(new_n795), .B1(G68), .B2(new_n797), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT121), .Z(new_n1191));
  AOI22_X1  g0991(.A1(G97), .A2(new_n753), .B1(new_n763), .B2(G303), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n801), .B2(new_n730), .C1(new_n389), .C2(new_n736), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n269), .B1(new_n747), .B2(new_n346), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT122), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n750), .A2(new_n804), .B1(new_n732), .B2(new_n505), .ZN(new_n1196));
  NOR4_X1   g0996(.A1(new_n1193), .A2(new_n1195), .A3(new_n1011), .A4(new_n1196), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT123), .Z(new_n1198));
  OAI21_X1  g0998(.A(new_n344), .B1(new_n750), .B2(new_n808), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n736), .A2(new_n809), .B1(new_n1136), .B2(new_n730), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(G50), .C2(new_n740), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n763), .A2(G128), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G159), .A2(new_n753), .B1(new_n758), .B2(new_n1045), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1201), .A2(new_n1151), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1198), .A2(new_n1204), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1191), .B1(new_n1014), .B2(new_n1205), .C1(new_n871), .C2(new_n829), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n1115), .B2(new_n1178), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n938), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1208), .B1(new_n1209), .B2(new_n1212), .ZN(G381));
  OR2_X1    g1013(.A1(G393), .A2(G396), .ZN(new_n1214));
  OR4_X1    g1014(.A1(G384), .A2(G390), .A3(G387), .A4(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1131), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1188), .A2(new_n1216), .ZN(new_n1217));
  OR3_X1    g1017(.A1(new_n1215), .A2(G381), .A3(new_n1217), .ZN(G407));
  OAI211_X1 g1018(.A(G407), .B(G213), .C1(G343), .C2(new_n1217), .ZN(G409));
  XOR2_X1   g1019(.A(G393), .B(G396), .Z(new_n1220));
  NAND2_X1  g1020(.A1(G387), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(KEYINPUT126), .B1(new_n957), .B2(new_n984), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1221), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(G390), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1221), .B(G390), .C1(new_n1220), .C2(new_n1222), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1182), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1185), .A2(KEYINPUT57), .A3(new_n1177), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n683), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1179), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1231), .A2(new_n1132), .A3(new_n1134), .A4(new_n1232), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1185), .A2(new_n1177), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1179), .B1(new_n1234), .B2(new_n1211), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1235), .A2(new_n1131), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1233), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(G213), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1239), .A2(G343), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT60), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n683), .B1(new_n1210), .B2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1119), .A2(new_n1120), .A3(KEYINPUT60), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1243), .B1(new_n1244), .B2(new_n1210), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n838), .B1(new_n1245), .B2(new_n1207), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1245), .A2(new_n838), .A3(new_n1207), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1238), .A2(new_n1241), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT62), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT127), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT61), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1240), .B1(new_n1233), .B2(new_n1237), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1244), .A2(new_n1210), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1243), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(G384), .A3(new_n1208), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT125), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n1259), .A3(new_n1246), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1240), .A2(G2897), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(KEYINPUT125), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1259), .B(new_n1261), .C1(new_n1258), .C2(new_n1246), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1252), .B(new_n1253), .C1(new_n1254), .C2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT62), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1254), .A2(new_n1270), .A3(new_n1249), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1251), .A2(new_n1269), .A3(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1266), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1236), .B1(G378), .B2(new_n1188), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1273), .B1(new_n1274), .B2(new_n1240), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1252), .B1(new_n1275), .B2(new_n1253), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1228), .B1(new_n1272), .B2(new_n1276), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1227), .B(new_n1253), .C1(new_n1254), .C2(new_n1268), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT63), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1250), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT124), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1254), .A2(KEYINPUT63), .A3(new_n1249), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT124), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1250), .A2(new_n1284), .A3(new_n1280), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1279), .A2(new_n1282), .A3(new_n1283), .A4(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1277), .A2(new_n1286), .ZN(G405));
  INV_X1    g1087(.A(new_n1249), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1227), .B(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1233), .B1(new_n1131), .B2(new_n1188), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1289), .B(new_n1290), .ZN(G402));
endmodule


