//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n564, new_n565,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(KEYINPUT3), .A3(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n470), .A2(new_n473), .A3(G137), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n465), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(KEYINPUT70), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT70), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n465), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n473), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n475), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G125), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT67), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G113), .ZN(new_n487));
  OR3_X1    g062(.A1(new_n487), .A2(new_n467), .A3(KEYINPUT68), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT68), .B1(new_n487), .B2(new_n467), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n486), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NOR3_X1   g065(.A1(new_n484), .A2(KEYINPUT67), .A3(new_n485), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n482), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n481), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G160));
  OAI221_X1 g069(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n473), .C2(G112), .ZN(new_n495));
  XOR2_X1   g070(.A(new_n495), .B(KEYINPUT71), .Z(new_n496));
  INV_X1    g071(.A(G124), .ZN(new_n497));
  INV_X1    g072(.A(new_n475), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(new_n482), .ZN(new_n500));
  INV_X1    g075(.A(G136), .ZN(new_n501));
  INV_X1    g076(.A(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  OAI221_X1 g078(.A(new_n496), .B1(new_n497), .B2(new_n500), .C1(new_n501), .C2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G162));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(G114), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(G2105), .ZN(new_n508));
  AND2_X1   g083(.A1(G126), .A2(G2105), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n470), .A2(new_n475), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT72), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n470), .A2(new_n512), .A3(new_n475), .A4(new_n509), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n508), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n473), .A2(G138), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(new_n499), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n517), .A2(KEYINPUT4), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n515), .A2(new_n519), .ZN(G164));
  XNOR2_X1  g095(.A(KEYINPUT5), .B(G543), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT6), .B(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G50), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G651), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n527), .A2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  INV_X1    g109(.A(G89), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n523), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n536), .B(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n539));
  INV_X1    g114(.A(G51), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n525), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n541), .B(new_n542), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n538), .A2(new_n543), .ZN(G168));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  INV_X1    g120(.A(G52), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n523), .A2(new_n545), .B1(new_n525), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n529), .ZN(new_n549));
  OR3_X1    g124(.A1(new_n547), .A2(new_n549), .A3(KEYINPUT75), .ZN(new_n550));
  OAI21_X1  g125(.A(KEYINPUT75), .B1(new_n547), .B2(new_n549), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(G171));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  INV_X1    g128(.A(G43), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n523), .A2(new_n553), .B1(new_n525), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT76), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n529), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT77), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XNOR2_X1  g138(.A(KEYINPUT78), .B(KEYINPUT8), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT79), .ZN(new_n565));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  NAND2_X1  g143(.A1(new_n523), .A2(KEYINPUT80), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT80), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n521), .A2(new_n522), .A3(new_n570), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G91), .ZN(new_n573));
  INV_X1    g148(.A(G543), .ZN(new_n574));
  OR2_X1    g149(.A1(KEYINPUT6), .A2(G651), .ZN(new_n575));
  NAND2_X1  g150(.A1(KEYINPUT6), .A2(G651), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G53), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT9), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n521), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(new_n529), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n573), .A2(new_n579), .A3(new_n581), .ZN(G299));
  INV_X1    g157(.A(G171), .ZN(G301));
  NAND2_X1  g158(.A1(new_n538), .A2(new_n543), .ZN(G286));
  NAND3_X1  g159(.A1(new_n569), .A2(G87), .A3(new_n571), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n521), .A2(G74), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(new_n577), .B2(G49), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT81), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n588), .B1(new_n585), .B2(new_n587), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n589), .A2(new_n590), .ZN(G288));
  NAND2_X1  g166(.A1(new_n572), .A2(G86), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  XOR2_X1   g168(.A(KEYINPUT5), .B(G543), .Z(new_n594));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(new_n577), .B2(G48), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n592), .A2(new_n597), .ZN(G305));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  XNOR2_X1  g174(.A(KEYINPUT82), .B(G47), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n523), .A2(new_n599), .B1(new_n525), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(new_n529), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NOR2_X1   g181(.A1(G301), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n572), .A2(G92), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n572), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(G79), .A2(G543), .ZN(new_n613));
  INV_X1    g188(.A(G66), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n594), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n615), .A2(G651), .B1(new_n577), .B2(G54), .ZN(new_n616));
  AND3_X1   g191(.A1(new_n612), .A2(KEYINPUT83), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g192(.A(KEYINPUT83), .B1(new_n612), .B2(new_n616), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n607), .B1(new_n619), .B2(new_n606), .ZN(G284));
  AOI21_X1  g195(.A(new_n607), .B1(new_n619), .B2(new_n606), .ZN(G321));
  NAND2_X1  g196(.A1(G299), .A2(new_n606), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G168), .B2(new_n606), .ZN(G297));
  OAI21_X1  g198(.A(new_n622), .B1(G168), .B2(new_n606), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n619), .B1(new_n625), .B2(G860), .ZN(G148));
  OAI21_X1  g201(.A(KEYINPUT84), .B1(new_n560), .B2(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n619), .A2(new_n625), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  MUX2_X1   g204(.A(KEYINPUT84), .B(new_n627), .S(new_n629), .Z(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g206(.A(new_n500), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G123), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT85), .ZN(new_n634));
  OAI221_X1 g209(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n473), .C2(G111), .ZN(new_n635));
  INV_X1    g210(.A(G135), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n503), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2096), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n464), .A2(new_n475), .A3(new_n483), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2100), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n639), .A2(new_n643), .ZN(G156));
  XOR2_X1   g219(.A(KEYINPUT15), .B(G2435), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2438), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2430), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT86), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n646), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(KEYINPUT14), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n651), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(G14), .A3(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2072), .B(G2078), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT18), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n664), .A2(new_n665), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n669), .A2(new_n663), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT87), .B(KEYINPUT17), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n664), .B(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n665), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n670), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n672), .A2(new_n673), .A3(new_n663), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n668), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(G2096), .Z(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT88), .B(G2100), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n682), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT89), .ZN(new_n690));
  OR3_X1    g265(.A1(new_n682), .A2(new_n685), .A3(new_n688), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n687), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n692), .B(new_n693), .Z(new_n694));
  XOR2_X1   g269(.A(G1991), .B(G1996), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n694), .A2(new_n695), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n694), .A2(new_n695), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n700), .A2(new_n697), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G229));
  XOR2_X1   g279(.A(KEYINPUT91), .B(G16), .Z(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(G22), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n706), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1971), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n585), .A2(new_n587), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n711), .B2(G23), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT33), .B(G1976), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n709), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  MUX2_X1   g290(.A(G6), .B(G305), .S(G16), .Z(new_n716));
  XOR2_X1   g291(.A(KEYINPUT32), .B(G1981), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n715), .B(new_n718), .C1(new_n713), .C2(new_n714), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(KEYINPUT34), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT92), .ZN(new_n721));
  OAI221_X1 g296(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n473), .C2(G107), .ZN(new_n722));
  INV_X1    g297(.A(G131), .ZN(new_n723));
  INV_X1    g298(.A(G119), .ZN(new_n724));
  OAI221_X1 g299(.A(new_n722), .B1(new_n503), .B2(new_n723), .C1(new_n724), .C2(new_n500), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G29), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G25), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT90), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT35), .B(G1991), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n706), .A2(G24), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n604), .B2(new_n706), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G1986), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n721), .B(new_n736), .C1(KEYINPUT34), .C2(new_n719), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT36), .ZN(new_n738));
  NOR2_X1   g313(.A1(G5), .A2(G16), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G171), .B2(G16), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1961), .ZN(new_n741));
  INV_X1    g316(.A(G2084), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n727), .B1(KEYINPUT24), .B2(G34), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(KEYINPUT24), .B2(G34), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n493), .B2(G29), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n741), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n705), .A2(G19), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT94), .Z(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n560), .B2(new_n705), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(G1341), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n705), .A2(G20), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT23), .ZN(new_n752));
  INV_X1    g327(.A(G299), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(new_n711), .ZN(new_n754));
  INV_X1    g329(.A(G1956), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n746), .A2(new_n750), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n711), .A2(G21), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G168), .B2(new_n711), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G1966), .ZN(new_n760));
  NOR2_X1   g335(.A1(G29), .A2(G35), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G162), .B2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT29), .B(G2090), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT25), .ZN(new_n765));
  NAND2_X1  g340(.A1(G103), .A2(G2104), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n765), .B1(new_n482), .B2(new_n766), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n473), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n768));
  NAND2_X1  g343(.A1(G115), .A2(G2104), .ZN(new_n769));
  INV_X1    g344(.A(G127), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n484), .B2(new_n770), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n767), .A2(new_n768), .B1(new_n771), .B2(new_n482), .ZN(new_n772));
  INV_X1    g347(.A(G139), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n503), .ZN(new_n774));
  MUX2_X1   g349(.A(G33), .B(new_n774), .S(G29), .Z(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(G2072), .Z(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT31), .B(G11), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT30), .B(G28), .Z(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(G29), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n638), .B2(G29), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n776), .B(new_n780), .C1(new_n742), .C2(new_n745), .ZN(new_n781));
  NOR4_X1   g356(.A1(new_n757), .A2(new_n760), .A3(new_n764), .A4(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G4), .A2(G16), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n619), .B2(G16), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT93), .B(G1348), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT97), .B(KEYINPUT28), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n727), .A2(G26), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  OAI221_X1 g365(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n473), .C2(G116), .ZN(new_n791));
  INV_X1    g366(.A(G140), .ZN(new_n792));
  INV_X1    g367(.A(G128), .ZN(new_n793));
  OAI221_X1 g368(.A(new_n791), .B1(new_n503), .B2(new_n792), .C1(new_n793), .C2(new_n500), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT95), .ZN(new_n795));
  AND3_X1   g370(.A1(new_n795), .A2(KEYINPUT96), .A3(G29), .ZN(new_n796));
  AOI21_X1  g371(.A(KEYINPUT96), .B1(new_n795), .B2(G29), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n790), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2067), .ZN(new_n799));
  NAND3_X1  g374(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT26), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n464), .A2(G105), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G141), .ZN(new_n805));
  INV_X1    g380(.A(G129), .ZN(new_n806));
  OAI221_X1 g381(.A(new_n804), .B1(new_n503), .B2(new_n805), .C1(new_n806), .C2(new_n500), .ZN(new_n807));
  MUX2_X1   g382(.A(G32), .B(new_n807), .S(G29), .Z(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT27), .Z(new_n809));
  NOR2_X1   g384(.A1(new_n809), .A2(G1996), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(G1996), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n727), .A2(G27), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G164), .B2(new_n727), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT98), .B(G2078), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  NOR4_X1   g391(.A1(new_n787), .A2(new_n799), .A3(new_n810), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n738), .A2(new_n817), .ZN(G150));
  INV_X1    g393(.A(G150), .ZN(G311));
  NAND2_X1  g394(.A1(new_n619), .A2(G559), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(G93), .ZN(new_n823));
  INV_X1    g398(.A(G55), .ZN(new_n824));
  OAI22_X1  g399(.A1(new_n523), .A2(new_n823), .B1(new_n525), .B2(new_n824), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n826), .A2(new_n529), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n559), .B(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n822), .B(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT39), .ZN(new_n832));
  AOI21_X1  g407(.A(G860), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n832), .B2(new_n831), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n829), .A2(G860), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT100), .B(KEYINPUT37), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n834), .A2(new_n837), .ZN(G145));
  INV_X1    g413(.A(new_n519), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT101), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n511), .A2(new_n513), .ZN(new_n841));
  INV_X1    g416(.A(new_n508), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI211_X1 g418(.A(KEYINPUT101), .B(new_n508), .C1(new_n511), .C2(new_n513), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n839), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n795), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n725), .ZN(new_n847));
  OAI221_X1 g422(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n473), .C2(G118), .ZN(new_n848));
  INV_X1    g423(.A(G142), .ZN(new_n849));
  INV_X1    g424(.A(G130), .ZN(new_n850));
  OAI221_X1 g425(.A(new_n848), .B1(new_n503), .B2(new_n849), .C1(new_n850), .C2(new_n500), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT102), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n641), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n807), .B(new_n774), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n847), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n847), .A2(new_n855), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n504), .B(new_n493), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n638), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(G37), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n856), .A2(new_n860), .A3(new_n857), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g441(.A(new_n830), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n628), .B(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n612), .A2(new_n616), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(G299), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT41), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n753), .A2(new_n612), .A3(new_n616), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT103), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n875));
  INV_X1    g450(.A(new_n873), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n871), .B1(new_n870), .B2(new_n872), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n868), .A2(new_n874), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n870), .A2(new_n872), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n879), .B1(new_n881), .B2(new_n868), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n882), .A2(KEYINPUT42), .ZN(new_n883));
  XNOR2_X1  g458(.A(G305), .B(G290), .ZN(new_n884));
  XNOR2_X1  g459(.A(G166), .B(new_n710), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n882), .A2(KEYINPUT42), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n883), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n887), .B1(new_n883), .B2(new_n888), .ZN(new_n890));
  OAI21_X1  g465(.A(G868), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n829), .A2(new_n606), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(G295));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n892), .ZN(G331));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n880), .A2(KEYINPUT41), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT103), .B1(new_n896), .B2(new_n873), .ZN(new_n897));
  INV_X1    g472(.A(new_n874), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT106), .B1(G301), .B2(G168), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT106), .ZN(new_n900));
  NAND3_X1  g475(.A1(G171), .A2(G286), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n903));
  NAND3_X1  g478(.A1(G301), .A2(G168), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT105), .B1(G171), .B2(G286), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n902), .A2(new_n830), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n830), .B1(new_n902), .B2(new_n906), .ZN(new_n909));
  OAI22_X1  g484(.A1(new_n897), .A2(new_n898), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n902), .A2(new_n906), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n867), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n912), .A2(new_n881), .A3(new_n907), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n910), .A2(new_n886), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  AOI22_X1  g490(.A1(new_n878), .A2(new_n874), .B1(new_n912), .B2(new_n907), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n908), .A2(new_n880), .A3(new_n909), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n887), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n863), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n915), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n918), .A2(KEYINPUT107), .A3(new_n863), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI22_X1  g499(.A1(new_n912), .A2(new_n907), .B1(new_n873), .B2(new_n896), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n887), .B1(new_n917), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n914), .A2(new_n926), .A3(new_n863), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT43), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n895), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n922), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n886), .B1(new_n910), .B2(new_n913), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n920), .B1(new_n932), .B2(G37), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(new_n923), .A3(new_n914), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n931), .B1(new_n934), .B2(new_n930), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n929), .B1(new_n895), .B2(new_n935), .ZN(G397));
  INV_X1    g511(.A(KEYINPUT54), .ZN(new_n937));
  INV_X1    g512(.A(G2078), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n492), .A2(new_n478), .A3(G40), .A4(new_n480), .ZN(new_n939));
  INV_X1    g514(.A(G1384), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(new_n515), .B2(new_n519), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n942), .A2(G1384), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n845), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n944), .B1(new_n845), .B2(new_n945), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n938), .B(new_n943), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT53), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT50), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n845), .A2(new_n951), .A3(new_n940), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n939), .B1(new_n941), .B2(KEYINPUT50), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G1961), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT45), .B1(new_n845), .B2(new_n940), .ZN(new_n957));
  AND4_X1   g532(.A1(G40), .A2(new_n492), .A3(new_n478), .A4(new_n480), .ZN(new_n958));
  INV_X1    g533(.A(new_n945), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n958), .B1(G164), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n961), .A2(KEYINPUT53), .A3(new_n938), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n950), .A2(new_n956), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n937), .B1(new_n964), .B2(G301), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT122), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT118), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n481), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n481), .A2(new_n967), .ZN(new_n969));
  XOR2_X1   g544(.A(KEYINPUT119), .B(G2078), .Z(new_n970));
  NAND4_X1  g545(.A1(new_n492), .A2(KEYINPUT53), .A3(G40), .A4(new_n970), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n957), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n972), .B(new_n973), .C1(new_n947), .C2(new_n946), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n950), .A2(new_n956), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT121), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT121), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n950), .A2(new_n977), .A3(new_n956), .A4(new_n974), .ZN(new_n978));
  AND4_X1   g553(.A1(new_n966), .A2(new_n976), .A3(G171), .A4(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(G301), .B1(new_n975), .B2(KEYINPUT121), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n966), .B1(new_n980), .B2(new_n978), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n965), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT123), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(KEYINPUT123), .B(new_n965), .C1(new_n979), .C2(new_n981), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT61), .ZN(new_n986));
  XNOR2_X1  g561(.A(KEYINPUT56), .B(G2072), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n943), .B(new_n987), .C1(new_n946), .C2(new_n947), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n989));
  AOI21_X1  g564(.A(G1384), .B1(new_n839), .B2(new_n514), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n939), .B1(new_n990), .B2(new_n951), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n845), .A2(new_n940), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n991), .B1(new_n992), .B2(new_n951), .ZN(new_n993));
  AOI22_X1  g568(.A1(new_n988), .A2(new_n989), .B1(new_n993), .B2(new_n755), .ZN(new_n994));
  XNOR2_X1  g569(.A(G299), .B(KEYINPUT57), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n958), .B1(new_n990), .B2(KEYINPUT45), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n845), .A2(new_n945), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT110), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n845), .A2(new_n944), .A3(new_n945), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n997), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1001), .A2(KEYINPUT114), .A3(new_n987), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n994), .A2(new_n996), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n996), .B1(new_n994), .B2(new_n1002), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n986), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n619), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n845), .A2(new_n958), .A3(new_n940), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(G2067), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G1348), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n954), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT115), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(G1348), .B1(new_n952), .B2(new_n953), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1014), .A2(new_n1009), .A3(new_n1015), .ZN(new_n1016));
  OAI211_X1 g591(.A(KEYINPUT60), .B(new_n1007), .C1(new_n1013), .C2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT59), .ZN(new_n1018));
  INV_X1    g593(.A(G1996), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT58), .B(G1341), .Z(new_n1020));
  AOI22_X1  g595(.A1(new_n1001), .A2(new_n1019), .B1(new_n1008), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1018), .B1(new_n1021), .B2(new_n559), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1008), .A2(new_n1020), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1023), .B1(new_n1024), .B2(G1996), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1025), .A2(KEYINPUT59), .A3(new_n560), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1017), .A2(new_n1022), .A3(new_n1026), .ZN(new_n1027));
  OR3_X1    g602(.A1(new_n1013), .A2(new_n1016), .A3(KEYINPUT60), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT60), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(new_n1029), .A3(new_n619), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n988), .A2(new_n989), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n993), .A2(new_n755), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1002), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n995), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1034), .A2(KEYINPUT61), .A3(new_n1003), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1006), .A2(new_n1027), .A3(new_n1030), .A4(new_n1035), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1013), .A2(new_n1016), .A3(new_n1007), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1003), .B1(new_n1005), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1966), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n957), .B2(new_n960), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n952), .A2(new_n953), .A3(new_n742), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G286), .A2(G8), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1047), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g624(.A(G8), .B(new_n1049), .C1(new_n1043), .C2(G286), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  AOI211_X1 g626(.A(new_n1045), .B(new_n1049), .C1(new_n1043), .C2(G8), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1046), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G8), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1055), .B(new_n991), .C1(new_n992), .C2(new_n951), .ZN(new_n1056));
  INV_X1    g631(.A(G2090), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n951), .B1(new_n845), .B2(new_n940), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n958), .B1(new_n941), .B2(KEYINPUT50), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT113), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1056), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1971), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1024), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1054), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(G303), .A2(G8), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1065), .B(KEYINPUT55), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1008), .A2(G8), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1981), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n592), .A2(new_n1071), .A3(new_n597), .ZN(new_n1072));
  XOR2_X1   g647(.A(KEYINPUT112), .B(G86), .Z(new_n1073));
  OAI21_X1  g648(.A(new_n597), .B1(new_n523), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G1981), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1072), .A2(KEYINPUT49), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT49), .B1(new_n1075), .B2(new_n1072), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n710), .A2(G1976), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1008), .A2(G8), .A3(new_n1079), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1070), .A2(new_n1078), .B1(new_n1080), .B2(KEYINPUT52), .ZN(new_n1081));
  INV_X1    g656(.A(G1976), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT52), .B1(G288), .B2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1083), .A2(new_n1008), .A3(G8), .A4(new_n1079), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1084), .A2(KEYINPUT111), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(KEYINPUT111), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1081), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n954), .A2(G2090), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1054), .B1(new_n1063), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1087), .B1(new_n1067), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1053), .A2(new_n1068), .A3(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT117), .B1(new_n964), .B2(G301), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n950), .A2(new_n956), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1094), .A2(new_n1095), .A3(G301), .A4(new_n974), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n963), .A2(new_n1097), .A3(G171), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT120), .B1(new_n975), .B2(G171), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1093), .A2(new_n1096), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1092), .B1(new_n1100), .B2(new_n937), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n984), .A2(new_n985), .A3(new_n1039), .A4(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT63), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1080), .A2(KEYINPUT52), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1078), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1104), .B1(new_n1105), .B2(new_n1069), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1084), .A2(KEYINPUT111), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1086), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1063), .A2(new_n1089), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1110), .A2(G8), .A3(new_n1067), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1109), .B(new_n1111), .C1(new_n1067), .C2(new_n1064), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1043), .A2(G8), .A3(G168), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1103), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n1103), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1091), .B(new_n1115), .C1(new_n1067), .C2(new_n1090), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1112), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1093), .A2(new_n1098), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1043), .A2(G8), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1049), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(new_n1044), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n1050), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1123), .A2(KEYINPUT62), .A3(new_n1046), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT62), .B1(new_n1123), .B2(new_n1046), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1118), .B(new_n1119), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  OR3_X1    g701(.A1(new_n1078), .A2(G1976), .A3(G288), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1069), .B1(new_n1127), .B2(new_n1072), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1111), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1128), .B1(new_n1129), .B2(new_n1109), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1117), .A2(new_n1126), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1102), .A2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n973), .A2(new_n939), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1133), .A2(G1996), .A3(new_n807), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1134), .A2(KEYINPUT109), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(KEYINPUT109), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n795), .B(G2067), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n807), .A2(G1996), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1135), .A2(new_n1136), .B1(new_n1133), .B2(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n725), .A2(new_n731), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n725), .A2(new_n731), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1133), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT108), .B1(G290), .B2(G1986), .ZN(new_n1145));
  NAND2_X1  g720(.A1(G290), .A2(G1986), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1145), .B(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1144), .B1(new_n1133), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1132), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1133), .B1(new_n1137), .B2(new_n807), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n1150), .B(KEYINPUT124), .Z(new_n1151));
  NAND2_X1  g726(.A1(new_n1133), .A2(new_n1019), .ZN(new_n1152));
  XOR2_X1   g727(.A(new_n1152), .B(KEYINPUT46), .Z(new_n1153));
  NOR2_X1   g728(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1154), .B(KEYINPUT47), .Z(new_n1155));
  AND2_X1   g730(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n795), .A2(G2067), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1133), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NOR4_X1   g733(.A1(new_n973), .A2(G1986), .A3(G290), .A4(new_n939), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT48), .Z(new_n1160));
  NAND3_X1  g735(.A1(new_n1140), .A2(new_n1143), .A3(new_n1160), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1155), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1149), .A2(new_n1162), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g738(.A1(G227), .A2(KEYINPUT125), .A3(new_n459), .ZN(new_n1165));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n1166));
  AOI21_X1  g740(.A(new_n1166), .B1(new_n679), .B2(G319), .ZN(new_n1167));
  OAI21_X1  g741(.A(new_n661), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n1169));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g744(.A(KEYINPUT126), .B(new_n661), .C1(new_n1165), .C2(new_n1167), .ZN(new_n1171));
  NAND3_X1  g745(.A1(new_n1170), .A2(new_n703), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g746(.A(G37), .B1(new_n858), .B2(new_n861), .ZN(new_n1173));
  AOI21_X1  g747(.A(new_n1172), .B1(new_n1173), .B2(new_n864), .ZN(new_n1174));
  AOI21_X1  g748(.A(new_n922), .B1(new_n921), .B2(new_n923), .ZN(new_n1175));
  OAI211_X1 g749(.A(new_n1174), .B(KEYINPUT127), .C1(new_n1175), .C2(new_n931), .ZN(new_n1176));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n1177));
  AND3_X1   g751(.A1(new_n1170), .A2(new_n703), .A3(new_n1171), .ZN(new_n1178));
  NAND2_X1  g752(.A1(new_n865), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g753(.A(new_n1177), .B1(new_n935), .B2(new_n1179), .ZN(new_n1180));
  AND2_X1   g754(.A1(new_n1176), .A2(new_n1180), .ZN(G308));
  NAND2_X1  g755(.A1(new_n1176), .A2(new_n1180), .ZN(G225));
endmodule


