//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT24), .B(G110), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT73), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G128), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n195), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G110), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT23), .B1(new_n193), .B2(G119), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(new_n194), .ZN(new_n201));
  OR2_X1    g015(.A1(KEYINPUT66), .A2(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT66), .A2(G128), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n202), .A2(KEYINPUT23), .A3(G119), .A4(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n199), .B1(new_n201), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT74), .ZN(new_n206));
  OAI22_X1  g020(.A1(new_n192), .A2(new_n198), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n206), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G125), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(KEYINPUT75), .A3(G140), .ZN(new_n212));
  INV_X1    g026(.A(G140), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G125), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(G140), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g030(.A(KEYINPUT16), .B(new_n212), .C1(new_n216), .C2(KEYINPUT75), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT16), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G146), .ZN(new_n221));
  INV_X1    g035(.A(G146), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n217), .A2(new_n222), .A3(new_n219), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT76), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n201), .A2(new_n204), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(G110), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n191), .A2(KEYINPUT73), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n199), .A2(KEYINPUT24), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n199), .A2(KEYINPUT24), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT73), .ZN(new_n231));
  NOR3_X1   g045(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n198), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n201), .A2(new_n204), .A3(KEYINPUT76), .A4(new_n199), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n227), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n216), .A2(G146), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n236), .B1(new_n220), .B2(G146), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n210), .A2(new_n224), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT77), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n190), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n235), .A2(new_n237), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n226), .A2(G110), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT74), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n243), .B(new_n208), .C1(new_n198), .C2(new_n192), .ZN(new_n244));
  INV_X1    g058(.A(new_n223), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n222), .B1(new_n217), .B2(new_n219), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n241), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT77), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n241), .B(new_n239), .C1(new_n244), .C2(new_n247), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n240), .B1(new_n251), .B2(new_n190), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G217), .ZN(new_n254));
  INV_X1    g068(.A(G902), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n254), .B1(G234), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(G902), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n250), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n228), .A2(new_n232), .ZN(new_n261));
  INV_X1    g075(.A(new_n198), .ZN(new_n262));
  AOI22_X1  g076(.A1(KEYINPUT74), .A2(new_n242), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n224), .A2(new_n263), .A3(new_n208), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n239), .B1(new_n264), .B2(new_n241), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n190), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n190), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n250), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n255), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT25), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n266), .A2(KEYINPUT25), .A3(new_n255), .A4(new_n268), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n259), .B1(new_n273), .B2(new_n256), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT32), .ZN(new_n275));
  INV_X1    g089(.A(G237), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(new_n188), .A3(G210), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n277), .B(KEYINPUT27), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT26), .B(G101), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT11), .ZN(new_n282));
  INV_X1    g096(.A(G134), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n282), .B1(new_n283), .B2(G137), .ZN(new_n284));
  INV_X1    g098(.A(G137), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(KEYINPUT11), .A3(G134), .ZN(new_n286));
  INV_X1    g100(.A(G131), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n283), .A2(G137), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n284), .A2(new_n286), .A3(new_n287), .A4(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n288), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n283), .A2(G137), .ZN(new_n291));
  OAI21_X1  g105(.A(G131), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G143), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT1), .B1(new_n293), .B2(G146), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n222), .A2(G143), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(G146), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n196), .A2(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT1), .ZN(new_n298));
  AND4_X1   g112(.A1(new_n298), .A2(new_n295), .A3(new_n296), .A4(G128), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n289), .B(new_n292), .C1(new_n297), .C2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n284), .A2(new_n288), .A3(new_n286), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G131), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n302), .A2(new_n289), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT64), .ZN(new_n304));
  XNOR2_X1  g118(.A(G143), .B(G146), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT0), .B(G128), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AND2_X1   g121(.A1(KEYINPUT0), .A2(G128), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n295), .A2(new_n296), .ZN(new_n310));
  NOR2_X1   g124(.A1(KEYINPUT0), .A2(G128), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n310), .A2(new_n312), .A3(KEYINPUT64), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n307), .A2(new_n309), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n300), .B1(new_n303), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n197), .A2(G116), .ZN(new_n316));
  INV_X1    g130(.A(G116), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G119), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT2), .B(G113), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n319), .B1(new_n321), .B2(KEYINPUT68), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT68), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n321), .A2(new_n319), .A3(KEYINPUT69), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT69), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n316), .A2(new_n318), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n327), .B1(new_n328), .B2(new_n320), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT28), .B1(new_n315), .B2(new_n331), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n307), .A2(new_n309), .A3(new_n313), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n302), .A2(new_n289), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT28), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n322), .A2(new_n324), .B1(new_n326), .B2(new_n329), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n335), .A2(new_n336), .A3(new_n300), .A4(new_n337), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT67), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n300), .B(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT65), .B1(new_n303), .B2(new_n314), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n313), .A2(new_n309), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT65), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n343), .A2(new_n344), .A3(new_n334), .A4(new_n307), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n337), .B1(new_n341), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n281), .B1(new_n339), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n335), .A2(new_n300), .A3(new_n337), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n280), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT31), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT30), .B1(new_n341), .B2(new_n346), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n335), .A2(KEYINPUT30), .A3(new_n300), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n331), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n351), .B(new_n352), .C1(new_n353), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n348), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT30), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n342), .A2(new_n345), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n300), .B(KEYINPUT67), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n355), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n350), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT70), .B1(new_n363), .B2(new_n352), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n351), .B1(new_n353), .B2(new_n355), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT70), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n366), .A3(KEYINPUT31), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n357), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(G472), .A2(G902), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n275), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n275), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT71), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n353), .A2(new_n355), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n349), .A2(new_n281), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT29), .ZN(new_n378));
  AOI21_X1  g192(.A(G902), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OR3_X1    g193(.A1(new_n339), .A2(new_n347), .A3(KEYINPUT29), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n332), .A2(new_n338), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n315), .A2(new_n331), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT29), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n380), .A2(new_n384), .A3(new_n280), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n379), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G472), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n348), .A2(new_n356), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n365), .A2(new_n366), .A3(KEYINPUT31), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n366), .B1(new_n365), .B2(KEYINPUT31), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT71), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(new_n372), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n371), .A2(new_n374), .A3(new_n387), .A4(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT72), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n368), .A2(KEYINPUT71), .A3(new_n373), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n392), .B1(new_n391), .B2(new_n372), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n391), .A2(new_n369), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n400), .A2(new_n275), .B1(G472), .B2(new_n386), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT72), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n274), .B1(new_n396), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n314), .A2(G125), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n297), .A2(new_n299), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n211), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n188), .A2(G224), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n404), .A2(new_n406), .B1(KEYINPUT7), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT87), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n408), .B(new_n409), .ZN(new_n410));
  XOR2_X1   g224(.A(KEYINPUT85), .B(KEYINPUT8), .Z(new_n411));
  XNOR2_X1  g225(.A(G110), .B(G122), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n411), .B(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G107), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(G104), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT3), .ZN(new_n416));
  INV_X1    g230(.A(G104), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(G107), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n415), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G101), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT80), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n414), .A2(G104), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n421), .B1(new_n422), .B2(KEYINPUT3), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n421), .B(KEYINPUT3), .C1(new_n417), .C2(G107), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n419), .B(new_n420), .C1(new_n423), .C2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(G101), .B1(new_n418), .B2(new_n415), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n319), .A2(KEYINPUT5), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n316), .A2(KEYINPUT5), .ZN(new_n430));
  INV_X1    g244(.A(G113), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n326), .A2(new_n329), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n428), .A2(KEYINPUT86), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n433), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n426), .A2(new_n427), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT86), .B1(new_n428), .B2(new_n433), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n413), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT89), .ZN(new_n441));
  NOR3_X1   g255(.A1(new_n297), .A2(new_n299), .A3(G125), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n442), .B1(G125), .B2(new_n314), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT88), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT7), .A4(new_n407), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n404), .A2(new_n406), .A3(KEYINPUT7), .A4(new_n407), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT88), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n410), .A2(new_n440), .A3(new_n441), .A4(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n435), .A2(new_n436), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT82), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n426), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n417), .A2(G107), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n422), .B2(KEYINPUT3), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT80), .B1(new_n418), .B2(new_n416), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n454), .B1(new_n455), .B2(new_n424), .ZN(new_n456));
  OAI21_X1  g270(.A(G101), .B1(new_n456), .B2(KEYINPUT81), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n419), .B(KEYINPUT81), .C1(new_n423), .C2(new_n425), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n452), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n419), .B1(new_n423), .B2(new_n425), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT81), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n463), .A2(new_n451), .A3(G101), .A4(new_n458), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n460), .A2(KEYINPUT4), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT4), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n463), .A2(new_n466), .A3(G101), .A4(new_n458), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n467), .A2(new_n331), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n450), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n412), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n449), .A2(new_n470), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n408), .A2(new_n409), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n408), .A2(new_n409), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n472), .A2(new_n473), .B1(new_n445), .B2(new_n447), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n441), .B1(new_n474), .B2(new_n440), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n255), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  XOR2_X1   g290(.A(new_n443), .B(new_n407), .Z(new_n477));
  INV_X1    g291(.A(new_n412), .ZN(new_n478));
  AOI211_X1 g292(.A(new_n450), .B(new_n478), .C1(new_n465), .C2(new_n468), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT6), .ZN(new_n480));
  XOR2_X1   g294(.A(new_n412), .B(KEYINPUT84), .Z(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI22_X1  g296(.A1(new_n479), .A2(new_n480), .B1(new_n469), .B2(new_n482), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n465), .A2(new_n468), .ZN(new_n484));
  OAI211_X1 g298(.A(KEYINPUT6), .B(new_n481), .C1(new_n484), .C2(new_n450), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n477), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT90), .B1(new_n476), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n480), .B1(new_n469), .B2(new_n412), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n469), .A2(new_n482), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n477), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT90), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n410), .A2(new_n440), .A3(new_n448), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT89), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n470), .A3(new_n449), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n492), .A2(new_n493), .A3(new_n255), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n487), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(G210), .B1(G237), .B2(G902), .ZN(new_n499));
  XOR2_X1   g313(.A(new_n499), .B(KEYINPUT91), .Z(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n492), .A2(new_n255), .A3(new_n496), .A4(new_n499), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(G214), .B1(G237), .B2(G902), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT9), .B(G234), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(KEYINPUT78), .ZN(new_n506));
  OAI21_X1  g320(.A(G221), .B1(new_n506), .B2(G902), .ZN(new_n507));
  XOR2_X1   g321(.A(new_n507), .B(KEYINPUT79), .Z(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT83), .B(G469), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n298), .B1(G143), .B2(new_n222), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n310), .B1(new_n512), .B2(new_n193), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n305), .A2(new_n298), .A3(G128), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n426), .A2(new_n515), .A3(new_n427), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT10), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n297), .A2(new_n299), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n519), .A2(KEYINPUT10), .A3(new_n426), .A4(new_n427), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n467), .A2(new_n333), .ZN(new_n522));
  AOI211_X1 g336(.A(new_n334), .B(new_n521), .C1(new_n465), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n436), .A2(new_n405), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n303), .B1(new_n524), .B2(new_n516), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT12), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(G110), .B(G140), .ZN(new_n528));
  INV_X1    g342(.A(G227), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(G953), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n528), .B(new_n530), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n523), .A2(new_n527), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n531), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n467), .A2(new_n333), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n463), .A2(G101), .A3(new_n458), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n466), .B1(new_n535), .B2(new_n452), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(new_n536), .B2(new_n464), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n334), .B1(new_n537), .B2(new_n521), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n521), .B1(new_n465), .B2(new_n522), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n303), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n533), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n255), .B(new_n511), .C1(new_n532), .C2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(G469), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n531), .B1(new_n523), .B2(new_n527), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n538), .A2(new_n540), .A3(new_n533), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n544), .B1(new_n547), .B2(new_n255), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n509), .B1(new_n543), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(G475), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT92), .B(G143), .ZN(new_n551));
  INV_X1    g365(.A(G214), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n552), .A2(G237), .A3(G953), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n293), .A2(KEYINPUT92), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(G131), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT92), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n553), .B1(new_n559), .B2(G143), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n560), .B(new_n287), .C1(new_n553), .C2(new_n551), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n557), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT94), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n557), .A2(new_n558), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n557), .A2(new_n561), .A3(KEYINPUT94), .A4(new_n558), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n564), .A2(new_n247), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT18), .ZN(new_n568));
  OAI221_X1 g382(.A(new_n560), .B1(new_n568), .B2(new_n287), .C1(new_n553), .C2(new_n551), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n212), .B1(new_n216), .B2(KEYINPUT75), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(new_n222), .ZN(new_n571));
  OAI221_X1 g385(.A(new_n569), .B1(new_n571), .B2(new_n236), .C1(new_n568), .C2(new_n557), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(G113), .B(G122), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(new_n417), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n567), .A2(new_n575), .A3(new_n572), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n550), .B1(new_n579), .B2(new_n255), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n567), .A2(new_n575), .A3(new_n572), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT93), .ZN(new_n582));
  AOI21_X1  g396(.A(KEYINPUT19), .B1(new_n214), .B2(new_n215), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n570), .B2(KEYINPUT19), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(G146), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n582), .B1(new_n585), .B2(new_n246), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n221), .B(KEYINPUT93), .C1(G146), .C2(new_n584), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n557), .A2(new_n561), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n575), .B1(new_n589), .B2(new_n572), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n581), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(G475), .A2(G902), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT20), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT20), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n595), .B(new_n592), .C1(new_n581), .C2(new_n590), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n580), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(G952), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(G953), .ZN(new_n599));
  NAND2_X1  g413(.A1(G234), .A2(G237), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT21), .B(G898), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(G902), .A3(G953), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n317), .A2(G122), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n414), .B1(new_n606), .B2(KEYINPUT14), .ZN(new_n607));
  XNOR2_X1  g421(.A(G116), .B(G122), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OR2_X1    g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n607), .A2(new_n609), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n202), .A2(G143), .A3(new_n203), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n293), .A2(G128), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n283), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n283), .B1(new_n612), .B2(new_n613), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n610), .B(new_n611), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT13), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n613), .B(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n612), .ZN(new_n620));
  OAI21_X1  g434(.A(G134), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n608), .B(new_n414), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n614), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n506), .A2(new_n254), .A3(G953), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n617), .A2(new_n623), .A3(new_n625), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n255), .ZN(new_n630));
  INV_X1    g444(.A(G478), .ZN(new_n631));
  OAI22_X1  g445(.A1(new_n630), .A2(KEYINPUT96), .B1(KEYINPUT15), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT95), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n629), .B2(new_n255), .ZN(new_n634));
  AOI211_X1 g448(.A(KEYINPUT95), .B(G902), .C1(new_n627), .C2(new_n628), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n631), .A2(KEYINPUT15), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT96), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n637), .B1(new_n630), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n632), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n597), .A2(new_n605), .A3(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n549), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n503), .A2(new_n504), .A3(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n403), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(new_n420), .ZN(G3));
  INV_X1    g459(.A(new_n504), .ZN(new_n646));
  INV_X1    g460(.A(new_n499), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n647), .B1(new_n476), .B2(new_n486), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n646), .B1(new_n648), .B2(new_n502), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT33), .ZN(new_n650));
  AOI21_X1  g464(.A(KEYINPUT97), .B1(new_n617), .B2(new_n623), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n629), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n650), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n628), .A3(new_n627), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n631), .A2(G902), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(new_n636), .B2(new_n631), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n597), .A2(new_n659), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n649), .A2(new_n605), .A3(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(G472), .B1(new_n368), .B2(G902), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n274), .A2(new_n400), .A3(new_n663), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n664), .A2(new_n549), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n417), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G6));
  NOR2_X1   g483(.A1(new_n596), .A2(KEYINPUT99), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n580), .ZN(new_n671));
  INV_X1    g485(.A(new_n640), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n594), .A2(KEYINPUT99), .A3(new_n596), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n649), .A2(new_n605), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n665), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT35), .B(G107), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G9));
  AOI21_X1  g493(.A(new_n646), .B1(new_n501), .B2(new_n502), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT25), .B1(new_n252), .B2(new_n255), .ZN(new_n681));
  INV_X1    g495(.A(new_n272), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n256), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n267), .A2(KEYINPUT36), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n248), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n257), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n663), .A2(new_n400), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n680), .A2(new_n642), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT37), .B(G110), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G12));
  NAND2_X1  g507(.A1(new_n394), .A2(new_n395), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n401), .A2(KEYINPUT72), .A3(new_n374), .A4(new_n393), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n601), .B(KEYINPUT101), .Z(new_n697));
  INV_X1    g511(.A(G900), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n600), .A2(new_n698), .A3(G902), .A4(G953), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT100), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n671), .A2(new_n673), .A3(new_n672), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT102), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n688), .A2(new_n549), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n696), .A2(new_n649), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G128), .ZN(G30));
  XOR2_X1   g520(.A(new_n503), .B(KEYINPUT38), .Z(new_n707));
  NOR2_X1   g521(.A1(new_n315), .A2(new_n331), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n280), .B1(new_n375), .B2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n376), .ZN(new_n710));
  AOI21_X1  g524(.A(G902), .B1(new_n710), .B2(new_n382), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(G472), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n399), .A2(new_n371), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n597), .A2(new_n640), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n714), .A2(new_n504), .A3(new_n688), .A4(new_n715), .ZN(new_n716));
  OR3_X1    g530(.A1(new_n707), .A2(KEYINPUT103), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g531(.A(KEYINPUT103), .B1(new_n707), .B2(new_n716), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n701), .B(KEYINPUT39), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n549), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT40), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n717), .A2(new_n718), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G143), .ZN(G45));
  INV_X1    g538(.A(KEYINPUT104), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(new_n660), .B2(new_n701), .ZN(new_n726));
  INV_X1    g540(.A(new_n701), .ZN(new_n727));
  NOR4_X1   g541(.A1(new_n597), .A2(new_n659), .A3(KEYINPUT104), .A4(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n696), .A2(new_n649), .A3(new_n704), .A4(new_n729), .ZN(new_n730));
  XOR2_X1   g544(.A(KEYINPUT105), .B(G146), .Z(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G48));
  NOR2_X1   g546(.A1(new_n539), .A2(new_n303), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n531), .B1(new_n733), .B2(new_n523), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n525), .B(KEYINPUT12), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n540), .A2(new_n735), .A3(new_n533), .ZN(new_n736));
  AOI21_X1  g550(.A(G902), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n542), .B(new_n507), .C1(new_n544), .C2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n734), .A2(new_n736), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n255), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(G469), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(KEYINPUT106), .A3(new_n542), .A4(new_n507), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n696), .A2(new_n274), .A3(new_n661), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT41), .B(G113), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G15));
  NAND4_X1  g562(.A1(new_n696), .A2(new_n274), .A3(new_n675), .A4(new_n745), .ZN(new_n749));
  XNOR2_X1  g563(.A(KEYINPUT107), .B(G116), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G18));
  AND3_X1   g565(.A1(new_n740), .A2(new_n649), .A3(new_n744), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n687), .A2(new_n597), .A3(new_n605), .A4(new_n640), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n696), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G119), .ZN(G21));
  NAND2_X1  g570(.A1(new_n740), .A2(new_n744), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n648), .A2(new_n502), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n504), .A3(new_n715), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n363), .A2(new_n352), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n383), .A2(new_n281), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n356), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n369), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n274), .A2(new_n663), .A3(new_n605), .A4(new_n763), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n757), .A2(new_n759), .A3(new_n764), .ZN(new_n765));
  XOR2_X1   g579(.A(new_n765), .B(G122), .Z(G24));
  INV_X1    g580(.A(KEYINPUT108), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n663), .A2(new_n763), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n767), .B1(new_n688), .B2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n687), .A2(KEYINPUT108), .A3(new_n663), .A4(new_n763), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n729), .A3(new_n752), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G125), .ZN(G27));
  INV_X1    g587(.A(new_n500), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n774), .B1(new_n487), .B2(new_n497), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n507), .B1(new_n543), .B2(new_n548), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n502), .A2(new_n504), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n274), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n391), .A2(new_n372), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n779), .B1(new_n401), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n729), .A2(new_n778), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT42), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n726), .A2(new_n728), .A3(KEYINPUT42), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(new_n696), .A3(new_n274), .A4(new_n778), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(new_n287), .ZN(G33));
  NAND4_X1  g601(.A1(new_n696), .A2(new_n274), .A3(new_n703), .A4(new_n778), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G134), .ZN(G36));
  INV_X1    g603(.A(new_n547), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(KEYINPUT45), .ZN(new_n791));
  OAI21_X1  g605(.A(G469), .B1(new_n790), .B2(KEYINPUT45), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n544), .A2(new_n255), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n795), .A2(KEYINPUT46), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(KEYINPUT46), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n542), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n507), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n720), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT109), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n775), .A2(new_n777), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n659), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n597), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT43), .Z(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n689), .A3(new_n687), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n803), .B1(new_n808), .B2(KEYINPUT44), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n809), .B1(KEYINPUT44), .B2(new_n808), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n801), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(new_n285), .ZN(G39));
  XNOR2_X1  g626(.A(new_n799), .B(KEYINPUT47), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n729), .A2(new_n779), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n813), .A2(new_n696), .A3(new_n803), .A4(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(KEYINPUT110), .B(G140), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n815), .B(new_n816), .ZN(G42));
  INV_X1    g631(.A(new_n765), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n746), .A2(new_n749), .A3(new_n755), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT112), .ZN(new_n820));
  INV_X1    g634(.A(new_n605), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n664), .A2(new_n549), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n660), .A2(KEYINPUT113), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(new_n597), .B2(new_n659), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n597), .A2(new_n672), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n823), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n680), .A2(new_n822), .A3(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n691), .B(new_n828), .C1(new_n403), .C2(new_n643), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n640), .A2(new_n671), .A3(new_n673), .A4(new_n701), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n696), .A2(new_n704), .A3(new_n802), .A4(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n771), .A2(new_n729), .A3(new_n778), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n783), .A2(new_n785), .A3(new_n788), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n753), .B1(new_n694), .B2(new_n695), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n765), .B1(new_n752), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT112), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n838), .A3(new_n746), .A4(new_n749), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n820), .A2(new_n834), .A3(new_n835), .A4(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OR3_X1    g656(.A1(new_n687), .A2(KEYINPUT116), .A3(new_n727), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT116), .B1(new_n687), .B2(new_n727), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n759), .ZN(new_n846));
  INV_X1    g660(.A(new_n776), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n845), .A2(new_n714), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n705), .A2(new_n848), .A3(new_n730), .A4(new_n772), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(KEYINPUT52), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n705), .A2(new_n772), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n705), .A2(new_n772), .A3(KEYINPUT115), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n853), .A2(new_n730), .A3(new_n848), .A4(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n850), .B1(new_n855), .B2(KEYINPUT52), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n783), .A2(new_n785), .A3(new_n788), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n857), .A2(new_n829), .A3(new_n833), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n858), .A2(KEYINPUT114), .A3(new_n820), .A4(new_n839), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n842), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n849), .A2(KEYINPUT52), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(new_n850), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n842), .A2(KEYINPUT53), .A3(new_n859), .A4(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n860), .A2(KEYINPUT117), .A3(new_n861), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n864), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g683(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n842), .A2(new_n859), .A3(new_n866), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n819), .A2(new_n861), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n858), .A2(new_n872), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n871), .A2(new_n861), .B1(new_n856), .B2(new_n873), .ZN(new_n874));
  AOI22_X1  g688(.A1(new_n869), .A2(KEYINPUT54), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n745), .A2(new_n802), .ZN(new_n876));
  NOR4_X1   g690(.A1(new_n876), .A2(new_n714), .A3(new_n779), .A4(new_n601), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n660), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n274), .A2(new_n663), .A3(new_n763), .ZN(new_n879));
  INV_X1    g693(.A(new_n697), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n806), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n752), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n878), .A2(new_n883), .A3(new_n599), .ZN(new_n884));
  INV_X1    g698(.A(new_n876), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(new_n880), .A3(new_n806), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT119), .Z(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n781), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(KEYINPUT48), .Z(new_n889));
  INV_X1    g703(.A(KEYINPUT51), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n743), .A2(new_n542), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n813), .B1(new_n509), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(new_n802), .A3(new_n882), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n887), .A2(new_n771), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n707), .A2(new_n882), .A3(new_n646), .A4(new_n745), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT50), .Z(new_n896));
  NAND3_X1  g710(.A1(new_n877), .A2(new_n597), .A3(new_n659), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n893), .A2(new_n894), .A3(new_n896), .A4(new_n897), .ZN(new_n898));
  AOI211_X1 g712(.A(new_n884), .B(new_n889), .C1(new_n890), .C2(new_n898), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n875), .B(new_n899), .C1(new_n890), .C2(new_n898), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n598), .A2(new_n188), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n804), .A2(new_n504), .A3(new_n509), .A4(new_n597), .ZN(new_n903));
  AOI211_X1 g717(.A(new_n779), .B(new_n903), .C1(KEYINPUT49), .C2(new_n891), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT111), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT49), .ZN(new_n906));
  INV_X1    g720(.A(new_n891), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n714), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n905), .A2(new_n707), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n902), .A2(new_n909), .ZN(G75));
  NOR2_X1   g724(.A1(new_n188), .A2(G952), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n490), .B(KEYINPUT120), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT55), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n477), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n874), .A2(new_n255), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(G210), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT56), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n915), .A2(new_n500), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n914), .A2(new_n917), .ZN(new_n920));
  AOI211_X1 g734(.A(new_n911), .B(new_n918), .C1(new_n919), .C2(new_n920), .ZN(G51));
  XNOR2_X1  g735(.A(new_n874), .B(new_n870), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n794), .B(KEYINPUT57), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n741), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n915), .A2(new_n793), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n911), .B1(new_n925), .B2(new_n926), .ZN(G54));
  NAND2_X1  g741(.A1(KEYINPUT58), .A2(G475), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT121), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n915), .A2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n591), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n932), .A2(new_n933), .A3(new_n911), .ZN(G60));
  NAND2_X1  g748(.A1(G478), .A2(G902), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT59), .Z(new_n936));
  NAND2_X1  g750(.A1(new_n868), .A2(new_n867), .ZN(new_n937));
  AOI21_X1  g751(.A(KEYINPUT117), .B1(new_n860), .B2(new_n861), .ZN(new_n938));
  OAI21_X1  g752(.A(KEYINPUT54), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n874), .A2(new_n870), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n936), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n655), .B(KEYINPUT122), .ZN(new_n942));
  OAI21_X1  g756(.A(KEYINPUT123), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT123), .ZN(new_n944));
  INV_X1    g758(.A(new_n942), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n944), .B(new_n945), .C1(new_n875), .C2(new_n936), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n945), .A2(new_n936), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n911), .B1(new_n922), .B2(new_n947), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n943), .A2(new_n946), .A3(new_n948), .ZN(G63));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n950), .A2(KEYINPUT125), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n871), .A2(new_n861), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n856), .A2(new_n873), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(G217), .A2(G902), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT60), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n954), .A2(KEYINPUT124), .A3(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT124), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n874), .B2(new_n956), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n958), .A2(new_n960), .A3(new_n253), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n911), .B1(KEYINPUT125), .B2(new_n950), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n685), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n958), .B2(new_n960), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n951), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n958), .A2(new_n960), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n685), .ZN(new_n968));
  INV_X1    g782(.A(new_n951), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n968), .A2(new_n969), .A3(new_n961), .A4(new_n962), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n966), .A2(new_n970), .ZN(G66));
  AOI21_X1  g785(.A(new_n188), .B1(new_n603), .B2(G224), .ZN(new_n972));
  INV_X1    g786(.A(new_n829), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n820), .A2(new_n973), .A3(new_n839), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n972), .B1(new_n974), .B2(new_n188), .ZN(new_n975));
  INV_X1    g789(.A(G898), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n912), .B1(new_n976), .B2(G953), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n975), .B(new_n977), .ZN(G69));
  AND2_X1   g792(.A1(new_n361), .A2(new_n354), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(new_n584), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n811), .A2(new_n815), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n853), .A2(new_n730), .A3(new_n854), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n846), .A2(new_n781), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n801), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n981), .A2(new_n835), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n188), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n698), .A2(G953), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n980), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(G953), .B1(new_n529), .B2(new_n698), .ZN(new_n989));
  INV_X1    g803(.A(new_n980), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n989), .B1(new_n990), .B2(KEYINPUT126), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n723), .A2(new_n982), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n992), .A2(KEYINPUT62), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(KEYINPUT62), .ZN(new_n994));
  INV_X1    g808(.A(new_n403), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n995), .A2(new_n721), .A3(new_n802), .A4(new_n827), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n981), .A2(new_n993), .A3(new_n994), .A4(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n990), .B1(new_n997), .B2(new_n188), .ZN(new_n998));
  OR3_X1    g812(.A1(new_n988), .A2(new_n991), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n991), .B1(new_n988), .B2(new_n998), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(G72));
  NAND2_X1  g815(.A1(G472), .A2(G902), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT63), .Z(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT127), .Z(new_n1004));
  OAI21_X1  g818(.A(new_n1004), .B1(new_n985), .B2(new_n974), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n911), .B1(new_n1005), .B2(new_n377), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1004), .B1(new_n997), .B2(new_n974), .ZN(new_n1007));
  INV_X1    g821(.A(new_n709), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1003), .ZN(new_n1011));
  NOR3_X1   g825(.A1(new_n1008), .A2(new_n377), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1010), .B1(new_n869), .B2(new_n1012), .ZN(G57));
endmodule


