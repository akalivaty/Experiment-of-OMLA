//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939;
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G128), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n188), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G128), .ZN(new_n193));
  AOI22_X1  g007(.A1(new_n188), .A2(new_n190), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n188), .A2(G143), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n189), .A2(G146), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n194), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G137), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT11), .A3(G134), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(G137), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n203), .A2(new_n205), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n207), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n202), .A2(G137), .ZN(new_n210));
  OAI21_X1  g024(.A(G131), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n200), .A2(new_n208), .A3(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n203), .A2(new_n207), .A3(new_n205), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G131), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n208), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT0), .A2(G128), .ZN(new_n216));
  XNOR2_X1  g030(.A(G143), .B(G146), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n197), .A2(new_n198), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT0), .B(G128), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT64), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n215), .A2(KEYINPUT65), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT65), .B1(new_n215), .B2(new_n223), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n187), .B(new_n212), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n212), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n215), .A2(new_n223), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT68), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n215), .A2(new_n223), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n227), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n226), .B1(new_n232), .B2(new_n187), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT2), .B(G113), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G119), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(G116), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G116), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT66), .B(G119), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n235), .B(new_n238), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n236), .A2(KEYINPUT66), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G119), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n239), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n234), .B1(new_n245), .B2(new_n237), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n241), .A2(new_n246), .A3(KEYINPUT67), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n238), .B1(new_n240), .B2(new_n239), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n249), .A3(new_n234), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n250), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n247), .A2(KEYINPUT69), .A3(new_n250), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n233), .A2(new_n251), .B1(new_n256), .B2(new_n232), .ZN(new_n257));
  XOR2_X1   g071(.A(KEYINPUT26), .B(G101), .Z(new_n258));
  NOR2_X1   g072(.A1(G237), .A2(G953), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G210), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n258), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT31), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n257), .A2(KEYINPUT31), .A3(new_n264), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n256), .A2(new_n232), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n212), .B1(new_n224), .B2(new_n225), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(new_n251), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n272), .B1(new_n271), .B2(new_n251), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT28), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n256), .A2(new_n228), .A3(new_n212), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n263), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n269), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(G472), .A2(G902), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n283), .B(KEYINPUT72), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT32), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT32), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n282), .A2(new_n287), .A3(new_n284), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n256), .B(new_n232), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n289), .A2(KEYINPUT28), .B1(new_n279), .B2(KEYINPUT74), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(KEYINPUT74), .A3(KEYINPUT28), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n291), .A2(KEYINPUT29), .A3(new_n264), .A4(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n280), .A2(new_n263), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n257), .A2(new_n264), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT29), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT73), .B1(new_n257), .B2(new_n264), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n293), .B(new_n294), .C1(new_n295), .C2(new_n301), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n286), .A2(new_n288), .B1(new_n302), .B2(G472), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n242), .A2(new_n244), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G128), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n305), .B1(new_n236), .B2(G128), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT24), .B(G110), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT77), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT77), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n306), .A2(new_n310), .A3(new_n307), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT75), .B(KEYINPUT23), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n312), .B1(new_n304), .B2(G128), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n195), .A2(KEYINPUT23), .A3(G119), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n305), .A3(new_n314), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n309), .B(new_n311), .C1(G110), .C2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(G125), .B(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n188), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT16), .ZN(new_n319));
  INV_X1    g133(.A(G140), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(G125), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n320), .A2(KEYINPUT76), .A3(G125), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n322), .B1(new_n317), .B2(KEYINPUT76), .ZN(new_n323));
  OAI211_X1 g137(.A(G146), .B(new_n321), .C1(new_n323), .C2(new_n319), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n316), .A2(new_n318), .A3(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n321), .B1(new_n323), .B2(new_n319), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n188), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n327), .A2(new_n324), .B1(G110), .B2(new_n315), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n328), .B1(new_n306), .B2(new_n307), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G953), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(G221), .A3(G234), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(KEYINPUT22), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(G137), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n325), .A2(new_n329), .A3(new_n334), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT25), .B1(new_n338), .B2(G902), .ZN(new_n339));
  INV_X1    g153(.A(G217), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n340), .B1(G234), .B2(new_n294), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT25), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n336), .A2(new_n342), .A3(new_n294), .A4(new_n337), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n339), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n338), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n341), .A2(G902), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n303), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G104), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT3), .B1(new_n350), .B2(G107), .ZN(new_n351));
  INV_X1    g165(.A(G107), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT78), .B1(new_n352), .B2(G104), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(new_n352), .A3(G104), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(new_n350), .A3(G107), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n351), .A2(new_n353), .A3(new_n355), .A4(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT4), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(G101), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n360), .B(new_n361), .ZN(new_n362));
  AND4_X1   g176(.A1(new_n351), .A2(new_n353), .A3(new_n355), .A4(new_n357), .ZN(new_n363));
  INV_X1    g177(.A(G101), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n358), .A2(G101), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(KEYINPUT4), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n251), .A2(new_n362), .A3(new_n367), .ZN(new_n368));
  OR2_X1    g182(.A1(new_n368), .A2(KEYINPUT84), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT5), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n245), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n371), .B(G113), .C1(new_n248), .C2(new_n370), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n352), .A2(G104), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n350), .A2(G107), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n364), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n375), .B1(new_n363), .B2(new_n364), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n372), .A2(new_n376), .A3(new_n241), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n368), .A2(KEYINPUT84), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n369), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  XOR2_X1   g193(.A(G110), .B(G122), .Z(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n380), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n369), .A2(new_n382), .A3(new_n377), .A4(new_n378), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(KEYINPUT6), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n200), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(G125), .ZN(new_n386));
  INV_X1    g200(.A(G125), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n387), .B1(new_n219), .B2(new_n222), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G224), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(G953), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n389), .B(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n379), .A2(new_n393), .A3(new_n380), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n384), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT7), .ZN(new_n396));
  AOI211_X1 g210(.A(new_n396), .B(new_n389), .C1(KEYINPUT88), .C2(new_n391), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n397), .B1(KEYINPUT88), .B2(new_n391), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n372), .A2(new_n241), .ZN(new_n399));
  INV_X1    g213(.A(new_n375), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(new_n358), .B2(G101), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT85), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(new_n377), .ZN(new_n404));
  XOR2_X1   g218(.A(new_n380), .B(KEYINPUT8), .Z(new_n405));
  NAND3_X1  g219(.A1(new_n399), .A2(KEYINPUT85), .A3(new_n401), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT86), .B(KEYINPUT7), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n389), .B1(new_n391), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(KEYINPUT87), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n383), .A2(new_n398), .A3(new_n407), .A4(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n395), .A2(new_n294), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(G210), .B1(G237), .B2(G902), .ZN(new_n413));
  XOR2_X1   g227(.A(new_n413), .B(KEYINPUT89), .Z(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(G214), .B1(G237), .B2(G902), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n395), .A2(new_n294), .A3(new_n411), .A4(new_n414), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(G110), .B(G140), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n331), .A2(G227), .ZN(new_n421));
  XOR2_X1   g235(.A(new_n420), .B(new_n421), .Z(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n215), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT10), .ZN(new_n425));
  NOR3_X1   g239(.A1(new_n385), .A2(new_n401), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT80), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n199), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n217), .A2(KEYINPUT80), .A3(new_n196), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n428), .A2(new_n194), .A3(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(KEYINPUT81), .B1(new_n430), .B2(new_n401), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT81), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n428), .A2(new_n429), .A3(new_n194), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n376), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n426), .B1(new_n435), .B2(new_n425), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n362), .A2(new_n367), .A3(new_n223), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n424), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n430), .A2(KEYINPUT81), .A3(new_n401), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n432), .B1(new_n376), .B2(new_n433), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n425), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n426), .ZN(new_n442));
  AND4_X1   g256(.A1(new_n424), .A2(new_n441), .A3(new_n437), .A4(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n423), .B1(new_n438), .B2(new_n443), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n441), .A2(new_n437), .A3(new_n424), .A4(new_n442), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT82), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT12), .B1(new_n215), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n431), .A2(new_n434), .B1(new_n401), .B2(new_n385), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n448), .B1(new_n449), .B2(new_n424), .ZN(new_n450));
  OAI22_X1  g264(.A1(new_n439), .A2(new_n440), .B1(new_n376), .B2(new_n200), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n215), .A3(new_n447), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n445), .A2(new_n450), .A3(new_n452), .A4(new_n422), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n444), .A2(KEYINPUT83), .A3(new_n453), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n453), .A2(KEYINPUT83), .ZN(new_n455));
  INV_X1    g269(.A(G469), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n454), .A2(new_n455), .A3(new_n456), .A4(new_n294), .ZN(new_n457));
  NAND2_X1  g271(.A1(G469), .A2(G902), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n441), .A2(new_n437), .A3(new_n442), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n215), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n423), .B1(new_n460), .B2(new_n445), .ZN(new_n461));
  AND4_X1   g275(.A1(new_n423), .A2(new_n445), .A3(new_n450), .A4(new_n452), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n457), .B(new_n458), .C1(new_n456), .C2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(KEYINPUT9), .B(G234), .ZN(new_n465));
  OAI21_X1  g279(.A(G221), .B1(new_n465), .B2(G902), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n419), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(G113), .B(G122), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(new_n350), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n317), .A2(KEYINPUT76), .ZN(new_n471));
  INV_X1    g285(.A(new_n322), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(KEYINPUT19), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT19), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n317), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT93), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n320), .A2(G125), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n387), .A2(G140), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n477), .A2(new_n478), .A3(new_n474), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT93), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n473), .A2(new_n476), .A3(new_n188), .A4(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT94), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n323), .A2(KEYINPUT19), .B1(new_n480), .B2(new_n479), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n485), .A2(KEYINPUT94), .A3(new_n188), .A4(new_n476), .ZN(new_n486));
  INV_X1    g300(.A(G237), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n331), .A3(G214), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n189), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n259), .A2(G143), .A3(G214), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n489), .A2(new_n206), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT92), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n489), .A2(new_n490), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(G131), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n489), .A2(KEYINPUT92), .A3(new_n206), .A4(new_n490), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n493), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n484), .A2(new_n486), .A3(new_n324), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(KEYINPUT18), .A2(G131), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n494), .B(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n323), .A2(G146), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n501), .A2(KEYINPUT91), .A3(new_n318), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT91), .B1(new_n501), .B2(new_n318), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n500), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n470), .B1(new_n498), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT17), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n493), .A2(new_n495), .A3(new_n506), .A4(new_n496), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n494), .A2(KEYINPUT17), .A3(G131), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n507), .A2(new_n327), .A3(new_n324), .A4(new_n508), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n504), .A2(new_n509), .A3(new_n470), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT20), .ZN(new_n512));
  INV_X1    g326(.A(G475), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n511), .A2(new_n512), .A3(new_n513), .A4(new_n294), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n513), .B(new_n294), .C1(new_n505), .C2(new_n510), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n504), .A2(new_n509), .ZN(new_n519));
  INV_X1    g333(.A(new_n470), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n504), .A2(new_n509), .A3(new_n470), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n513), .B1(new_n523), .B2(new_n294), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT95), .B1(new_n518), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT95), .ZN(new_n527));
  AOI211_X1 g341(.A(new_n527), .B(new_n524), .C1(new_n514), .C2(new_n517), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n331), .A2(G952), .ZN(new_n531));
  INV_X1    g345(.A(G234), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n531), .B1(new_n532), .B2(new_n487), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  AOI211_X1 g348(.A(new_n294), .B(new_n331), .C1(G234), .C2(G237), .ZN(new_n535));
  XOR2_X1   g349(.A(KEYINPUT21), .B(G898), .Z(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n534), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(G128), .B(G143), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT13), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n195), .A2(KEYINPUT13), .A3(G143), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(new_n202), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n540), .A2(new_n542), .B1(new_n202), .B2(new_n539), .ZN(new_n543));
  INV_X1    g357(.A(G122), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT96), .B1(new_n544), .B2(G116), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT96), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n239), .A3(G122), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n239), .A2(G122), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n551), .A2(G107), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n352), .B1(new_n548), .B2(new_n550), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n543), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n539), .B(new_n202), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n352), .B1(new_n550), .B2(KEYINPUT14), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n548), .B(new_n550), .C1(KEYINPUT14), .C2(new_n352), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n465), .A2(new_n340), .A3(G953), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT97), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n554), .A2(new_n559), .A3(new_n561), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n560), .A2(KEYINPUT97), .A3(new_n562), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n294), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G478), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n569), .A2(KEYINPUT15), .ZN(new_n570));
  XOR2_X1   g384(.A(new_n568), .B(new_n570), .Z(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n530), .A2(new_n538), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n349), .A2(new_n468), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(G101), .ZN(G3));
  INV_X1    g389(.A(new_n419), .ZN(new_n576));
  INV_X1    g390(.A(new_n538), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n563), .A2(KEYINPUT33), .A3(new_n565), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT98), .B(KEYINPUT33), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n566), .A2(new_n567), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT99), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n566), .A2(KEYINPUT99), .A3(new_n567), .A4(new_n580), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n579), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n569), .A2(G902), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT100), .ZN(new_n587));
  INV_X1    g401(.A(new_n568), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n587), .B1(new_n588), .B2(G478), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n568), .A2(KEYINPUT100), .A3(new_n569), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n585), .A2(new_n586), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n530), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n578), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n467), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n267), .A2(new_n268), .B1(new_n280), .B2(new_n263), .ZN(new_n596));
  OAI21_X1  g410(.A(G472), .B1(new_n596), .B2(G902), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n597), .A2(new_n285), .ZN(new_n598));
  INV_X1    g412(.A(new_n348), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n595), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT34), .B(G104), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G6));
  OAI21_X1  g417(.A(KEYINPUT101), .B1(new_n515), .B2(new_n516), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n604), .B(new_n517), .Z(new_n605));
  NOR4_X1   g419(.A1(new_n578), .A2(new_n571), .A3(new_n524), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n600), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT35), .B(G107), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G9));
  NOR2_X1   g423(.A1(new_n335), .A2(KEYINPUT36), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n330), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n346), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n344), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n468), .A2(new_n573), .A3(new_n598), .A4(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(new_n615), .B(KEYINPUT37), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(G110), .ZN(G12));
  NOR4_X1   g431(.A1(new_n303), .A2(new_n419), .A3(new_n467), .A4(new_n613), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT102), .B(G900), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n534), .B1(new_n535), .B2(new_n619), .ZN(new_n620));
  NOR4_X1   g434(.A1(new_n605), .A2(new_n571), .A3(new_n524), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT103), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G128), .ZN(G30));
  XNOR2_X1  g438(.A(new_n620), .B(KEYINPUT39), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n467), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n416), .A2(new_n418), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n629), .B(KEYINPUT38), .Z(new_n630));
  NAND2_X1  g444(.A1(new_n286), .A2(new_n288), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n294), .B1(new_n289), .B2(new_n264), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n257), .A2(new_n263), .ZN(new_n633));
  OAI21_X1  g447(.A(G472), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n529), .A2(new_n571), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n635), .A2(new_n417), .A3(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n628), .A2(new_n630), .A3(new_n613), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT105), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(new_n189), .ZN(G45));
  OR2_X1    g454(.A1(new_n303), .A2(new_n613), .ZN(new_n641));
  INV_X1    g455(.A(new_n620), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n592), .B(new_n642), .C1(new_n526), .C2(new_n528), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT106), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n419), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n643), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n576), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n467), .B1(new_n648), .B2(new_n644), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G146), .ZN(G48));
  INV_X1    g465(.A(KEYINPUT108), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n454), .A2(new_n294), .A3(new_n455), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(G469), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n654), .A2(KEYINPUT107), .A3(new_n457), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT107), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n653), .A2(new_n656), .A3(G469), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n652), .B1(new_n658), .B2(new_n466), .ZN(new_n659));
  INV_X1    g473(.A(new_n466), .ZN(new_n660));
  AOI211_X1 g474(.A(KEYINPUT108), .B(new_n660), .C1(new_n655), .C2(new_n657), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n662), .A2(new_n349), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n594), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT41), .B(G113), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G15));
  NAND2_X1  g480(.A1(new_n663), .A2(new_n606), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G116), .ZN(G18));
  INV_X1    g482(.A(new_n641), .ZN(new_n669));
  AOI21_X1  g483(.A(KEYINPUT109), .B1(new_n662), .B2(new_n576), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT109), .ZN(new_n671));
  NOR4_X1   g485(.A1(new_n659), .A2(new_n661), .A3(new_n671), .A4(new_n419), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n573), .B(new_n669), .C1(new_n670), .C2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G119), .ZN(G21));
  NAND3_X1  g488(.A1(new_n662), .A2(new_n576), .A3(new_n636), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n264), .B1(new_n291), .B2(new_n292), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n267), .A2(new_n268), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n284), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n678), .A2(new_n597), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n679), .A2(new_n599), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n577), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(new_n544), .ZN(G24));
  NAND2_X1  g497(.A1(new_n679), .A2(new_n614), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n643), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n685), .B1(new_n670), .B2(new_n672), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G125), .ZN(G27));
  INV_X1    g501(.A(KEYINPUT110), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n629), .A2(new_n417), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n349), .A2(new_n595), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n689), .B1(new_n691), .B2(new_n643), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n691), .A2(new_n689), .A3(new_n643), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n688), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n694), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(KEYINPUT110), .A3(new_n692), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G131), .ZN(G33));
  INV_X1    g513(.A(new_n690), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n467), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n349), .A3(new_n622), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n702), .B(KEYINPUT111), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G134), .ZN(G36));
  AOI21_X1  g518(.A(new_n613), .B1(new_n597), .B2(new_n285), .ZN(new_n705));
  AOI21_X1  g519(.A(KEYINPUT43), .B1(new_n529), .B2(new_n592), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n707));
  NOR4_X1   g521(.A1(new_n526), .A2(new_n528), .A3(new_n591), .A4(new_n707), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n705), .B(KEYINPUT44), .C1(new_n706), .C2(new_n708), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n709), .A2(KEYINPUT113), .A3(new_n690), .ZN(new_n710));
  AOI21_X1  g524(.A(KEYINPUT113), .B1(new_n709), .B2(new_n690), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n705), .B1(new_n706), .B2(new_n708), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n625), .ZN(new_n716));
  INV_X1    g530(.A(new_n457), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n718));
  OAI21_X1  g532(.A(KEYINPUT112), .B1(new_n463), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n456), .B1(new_n463), .B2(new_n718), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT112), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n721), .B(KEYINPUT45), .C1(new_n461), .C2(new_n462), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n458), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT46), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n717), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n723), .A2(KEYINPUT46), .A3(new_n458), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n660), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n715), .A2(new_n716), .A3(new_n728), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n712), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G137), .ZN(G39));
  INV_X1    g545(.A(KEYINPUT47), .ZN(new_n732));
  AOI211_X1 g546(.A(new_n732), .B(new_n660), .C1(new_n726), .C2(new_n727), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n724), .A2(new_n725), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n457), .A3(new_n727), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT47), .B1(new_n735), .B2(new_n466), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n647), .B(new_n690), .C1(new_n733), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n303), .A2(new_n348), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G140), .ZN(G42));
  INV_X1    g554(.A(new_n662), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n741), .A2(new_n533), .A3(new_n700), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n631), .A2(new_n599), .A3(new_n634), .ZN(new_n744));
  OR3_X1    g558(.A1(new_n743), .A2(KEYINPUT117), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT117), .B1(new_n743), .B2(new_n744), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n530), .A2(new_n592), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n706), .A2(new_n708), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n742), .A2(new_n614), .A3(new_n679), .A4(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n680), .A3(new_n534), .ZN(new_n751));
  NOR4_X1   g565(.A1(new_n741), .A2(new_n630), .A3(new_n751), .A4(new_n417), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT50), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n748), .A2(new_n750), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  AOI211_X1 g569(.A(new_n736), .B(new_n733), .C1(new_n660), .C2(new_n658), .ZN(new_n756));
  OR3_X1    g570(.A1(new_n756), .A2(new_n700), .A3(new_n751), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n755), .B(new_n757), .C1(KEYINPUT116), .C2(KEYINPUT51), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n748), .A2(new_n750), .A3(new_n753), .A4(new_n757), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n759), .B(new_n760), .C1(new_n754), .C2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n758), .A2(new_n531), .A3(new_n762), .ZN(new_n763));
  AND4_X1   g577(.A1(new_n530), .A2(new_n745), .A3(new_n592), .A4(new_n746), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n742), .A2(new_n349), .A3(new_n749), .ZN(new_n765));
  XOR2_X1   g579(.A(new_n765), .B(KEYINPUT48), .Z(new_n766));
  NOR3_X1   g580(.A1(new_n763), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n751), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n768), .B1(new_n670), .B2(new_n672), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n529), .A2(new_n572), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n593), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n600), .A2(new_n576), .A3(new_n577), .A4(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n615), .A3(new_n574), .ZN(new_n773));
  AOI22_X1  g587(.A1(new_n646), .A2(new_n649), .B1(new_n618), .B2(new_n622), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n686), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n629), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n614), .A2(new_n620), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n637), .A2(new_n776), .A3(new_n595), .A4(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n775), .A2(KEYINPUT52), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n686), .A2(new_n774), .A3(new_n778), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n773), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  NOR4_X1   g597(.A1(new_n605), .A2(new_n572), .A3(new_n524), .A4(new_n620), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT114), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n641), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n701), .B1(new_n786), .B2(new_n685), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n703), .A2(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n673), .A2(new_n667), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n664), .B1(new_n675), .B2(new_n681), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n698), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT53), .B1(new_n789), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n783), .A2(new_n788), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n798), .A2(new_n799), .A3(new_n795), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT54), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n696), .A2(new_n692), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n794), .A2(KEYINPUT115), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n805));
  OAI21_X1  g619(.A(KEYINPUT53), .B1(new_n793), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n789), .A2(new_n802), .A3(new_n804), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n799), .B1(new_n798), .B2(new_n795), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n767), .A2(new_n769), .A3(new_n801), .A4(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n812), .B1(G952), .B2(G953), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT49), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n417), .B1(new_n658), .B2(new_n814), .ZN(new_n815));
  AOI211_X1 g629(.A(new_n744), .B(new_n815), .C1(new_n814), .C2(new_n658), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n466), .ZN(new_n817));
  OR4_X1    g631(.A1(new_n530), .A2(new_n817), .A3(new_n591), .A4(new_n630), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n813), .A2(new_n818), .ZN(G75));
  NAND2_X1  g633(.A1(new_n384), .A2(new_n394), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(new_n392), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(KEYINPUT55), .Z(new_n822));
  INV_X1    g636(.A(new_n802), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n798), .A2(new_n803), .A3(new_n806), .A4(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(G902), .B1(new_n824), .B2(new_n797), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n415), .ZN(new_n826));
  OAI211_X1 g640(.A(KEYINPUT118), .B(new_n822), .C1(new_n826), .C2(KEYINPUT56), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n331), .A2(G952), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n294), .B1(new_n808), .B2(new_n810), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT56), .B1(new_n829), .B2(new_n414), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n822), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n833), .B1(new_n830), .B2(new_n831), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n827), .A2(new_n832), .A3(new_n834), .ZN(G51));
  NAND2_X1  g649(.A1(new_n458), .A2(KEYINPUT57), .ZN(new_n836));
  INV_X1    g650(.A(new_n811), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n809), .B1(new_n808), .B2(new_n810), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n458), .A2(KEYINPUT57), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n454), .B(new_n455), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n825), .A2(new_n723), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n828), .B1(new_n841), .B2(new_n842), .ZN(G54));
  NAND3_X1  g657(.A1(new_n829), .A2(KEYINPUT58), .A3(G475), .ZN(new_n844));
  INV_X1    g658(.A(new_n511), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n846), .A2(new_n847), .A3(new_n828), .ZN(G60));
  OAI21_X1  g662(.A(new_n585), .B1(new_n837), .B2(new_n838), .ZN(new_n849));
  NAND2_X1  g663(.A1(G478), .A2(G902), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n850), .B(KEYINPUT59), .Z(new_n851));
  NOR2_X1   g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n828), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n851), .B1(new_n801), .B2(new_n811), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(new_n854), .B2(new_n585), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n852), .A2(new_n855), .ZN(G63));
  NAND2_X1  g670(.A1(G217), .A2(G902), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT60), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n611), .B(new_n859), .C1(new_n824), .C2(new_n797), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n858), .B1(new_n808), .B2(new_n810), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n860), .B(new_n853), .C1(new_n345), .C2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n862), .A2(new_n863), .A3(KEYINPUT61), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT61), .B1(new_n862), .B2(new_n863), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(G66));
  OAI21_X1  g680(.A(G953), .B1(new_n537), .B2(new_n390), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n793), .A2(new_n773), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n867), .B1(new_n868), .B2(G953), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n869), .B(KEYINPUT120), .Z(new_n870));
  OAI21_X1  g684(.A(new_n820), .B1(G898), .B2(new_n331), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n870), .B(new_n871), .ZN(G69));
  AOI21_X1  g686(.A(new_n331), .B1(G227), .B2(G900), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n686), .A2(new_n638), .A3(new_n774), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT62), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n771), .A2(KEYINPUT121), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n349), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n593), .A2(new_n879), .A3(new_n770), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n690), .A2(new_n880), .A3(new_n626), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n876), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(new_n737), .B2(new_n738), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n690), .A2(new_n880), .A3(new_n626), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n884), .A2(KEYINPUT122), .A3(new_n349), .A4(new_n877), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(new_n712), .B2(new_n729), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n686), .A2(new_n638), .A3(new_n888), .A4(new_n774), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n875), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n331), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n485), .A2(new_n476), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n233), .B(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT123), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n891), .A2(new_n896), .A3(new_n893), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n703), .A2(new_n698), .A3(new_n739), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n728), .A2(new_n716), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n901), .A2(new_n576), .A3(new_n349), .A4(new_n636), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n775), .A2(new_n730), .A3(new_n902), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n899), .A2(G953), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(G900), .A2(G953), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n904), .A2(new_n893), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n873), .B1(new_n898), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n895), .A2(KEYINPUT124), .A3(new_n897), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n896), .B1(new_n891), .B2(new_n893), .ZN(new_n911));
  INV_X1    g725(.A(new_n893), .ZN(new_n912));
  AOI211_X1 g726(.A(KEYINPUT123), .B(new_n912), .C1(new_n890), .C2(new_n331), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n910), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  OR3_X1    g728(.A1(new_n904), .A2(new_n893), .A3(new_n906), .ZN(new_n915));
  INV_X1    g729(.A(new_n873), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n909), .A2(new_n914), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n917), .A2(KEYINPUT125), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n907), .B1(new_n898), .B2(new_n910), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n911), .A2(new_n913), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n873), .B1(new_n921), .B2(KEYINPUT124), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n919), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n908), .B1(new_n918), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI211_X1 g740(.A(KEYINPUT126), .B(new_n908), .C1(new_n918), .C2(new_n923), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(G72));
  NAND2_X1  g742(.A1(G472), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT63), .Z(new_n930));
  INV_X1    g744(.A(new_n868), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n930), .B1(new_n931), .B2(new_n890), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n633), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT127), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n931), .A2(new_n903), .A3(new_n899), .ZN(new_n935));
  INV_X1    g749(.A(new_n930), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n263), .B(new_n257), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n298), .A2(new_n265), .A3(new_n300), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n930), .B(new_n938), .C1(new_n797), .C2(new_n800), .ZN(new_n939));
  AND4_X1   g753(.A1(new_n853), .A2(new_n934), .A3(new_n937), .A4(new_n939), .ZN(G57));
endmodule


