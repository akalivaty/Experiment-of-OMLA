//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951;
  INV_X1    g000(.A(KEYINPUT34), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT25), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT24), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n204), .A2(G183gat), .A3(G190gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(G183gat), .B(G190gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(new_n204), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n203), .B1(new_n207), .B2(KEYINPUT65), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  INV_X1    g008(.A(G176gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(KEYINPUT64), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n214));
  NOR2_X1   g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n214), .B1(new_n215), .B2(KEYINPUT23), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G190gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(G183gat), .ZN(new_n219));
  INV_X1    g018(.A(G183gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(G190gat), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT24), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n224), .B1(KEYINPUT23), .B2(new_n215), .ZN(new_n225));
  AND3_X1   g024(.A1(new_n222), .A2(new_n225), .A3(new_n205), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n208), .A2(new_n217), .A3(new_n226), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n217), .A2(new_n225), .A3(new_n222), .A4(new_n205), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n222), .A2(new_n229), .A3(new_n205), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n203), .A3(new_n230), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n215), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT26), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n211), .A2(new_n234), .A3(new_n223), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(KEYINPUT27), .B(G183gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(new_n218), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT28), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n237), .A2(KEYINPUT28), .A3(new_n218), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n236), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT69), .B1(new_n232), .B2(new_n242), .ZN(new_n243));
  OR2_X1    g042(.A1(KEYINPUT66), .A2(G134gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(KEYINPUT66), .A2(G134gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(G127gat), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G127gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G134gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT67), .ZN(new_n249));
  INV_X1    g048(.A(G134gat), .ZN(new_n250));
  OR3_X1    g049(.A1(new_n250), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n246), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(G113gat), .B(G120gat), .Z(new_n253));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OR2_X1    g054(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n250), .A2(G127gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n258));
  AND4_X1   g057(.A1(new_n248), .A2(new_n256), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n252), .A2(new_n255), .B1(new_n259), .B2(new_n253), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n242), .B1(new_n227), .B2(new_n231), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n243), .A2(new_n263), .ZN(new_n264));
  OAI211_X1 g063(.A(KEYINPUT69), .B(new_n260), .C1(new_n232), .C2(new_n242), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G227gat), .ZN(new_n267));
  INV_X1    g066(.A(G233gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n202), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  AOI211_X1 g070(.A(KEYINPUT34), .B(new_n269), .C1(new_n264), .C2(new_n265), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n264), .A2(new_n269), .A3(new_n265), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT32), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT33), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G15gat), .B(G43gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT70), .ZN(new_n279));
  INV_X1    g078(.A(G71gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G99gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n275), .A2(new_n277), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n283), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n274), .B(KEYINPUT32), .C1(new_n276), .C2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n273), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n273), .A2(new_n284), .A3(KEYINPUT72), .A4(new_n286), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n292));
  XNOR2_X1  g091(.A(G141gat), .B(G148gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G155gat), .ZN(new_n295));
  INV_X1    g094(.A(G162gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(KEYINPUT2), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n294), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n298), .B(new_n297), .C1(new_n293), .C2(KEYINPUT2), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n292), .B1(new_n303), .B2(KEYINPUT3), .ZN(new_n304));
  XNOR2_X1  g103(.A(G197gat), .B(G204gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT22), .ZN(new_n306));
  INV_X1    g105(.A(G211gat), .ZN(new_n307));
  INV_X1    g106(.A(G218gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n305), .A3(new_n309), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(KEYINPUT73), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n314), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n304), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n303), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n313), .A2(KEYINPUT84), .A3(new_n314), .ZN(new_n321));
  OR2_X1    g120(.A1(new_n314), .A2(KEYINPUT84), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(new_n322), .A3(new_n292), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT3), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n320), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G228gat), .ZN(new_n326));
  OAI22_X1  g125(.A1(new_n319), .A2(new_n325), .B1(new_n326), .B2(new_n268), .ZN(new_n327));
  INV_X1    g126(.A(G22gat), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT29), .B1(new_n313), .B2(new_n314), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n303), .B1(new_n329), .B2(KEYINPUT3), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT85), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n304), .A2(new_n315), .A3(new_n318), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n326), .A2(new_n268), .ZN(new_n334));
  OAI211_X1 g133(.A(KEYINPUT85), .B(new_n303), .C1(new_n329), .C2(KEYINPUT3), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n327), .A2(new_n328), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n328), .B1(new_n327), .B2(new_n336), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT83), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G78gat), .B(G106gat), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n340), .B(KEYINPUT82), .Z(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT31), .B(G50gat), .ZN(new_n343));
  INV_X1    g142(.A(new_n341), .ZN(new_n344));
  OAI211_X1 g143(.A(KEYINPUT83), .B(new_n344), .C1(new_n337), .C2(new_n338), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n343), .B1(new_n342), .B2(new_n345), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n284), .A2(new_n286), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n349), .B1(new_n271), .B2(new_n272), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n291), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(G1gat), .B(G29gat), .Z(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G57gat), .B(G85gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G225gat), .A2(G233gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n252), .A2(new_n255), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n259), .A2(new_n253), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(new_n303), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT4), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n320), .A2(new_n324), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n303), .A2(KEYINPUT3), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT77), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n361), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n260), .A2(KEYINPUT77), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n358), .B(new_n363), .C1(new_n366), .C2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT78), .B1(new_n361), .B2(new_n303), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n320), .A2(new_n260), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n375), .A2(KEYINPUT4), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n372), .A2(new_n374), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n368), .A2(new_n303), .A3(new_n369), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n358), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT5), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT79), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n379), .A2(new_n372), .A3(new_n374), .ZN(new_n383));
  INV_X1    g182(.A(new_n358), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT79), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT5), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n377), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n358), .B1(new_n370), .B2(new_n366), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n389), .A2(KEYINPUT5), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT81), .B1(new_n362), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(new_n375), .B2(new_n391), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n372), .A2(new_n374), .A3(KEYINPUT81), .A4(KEYINPUT4), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n390), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n357), .B1(new_n388), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n386), .B1(new_n385), .B2(KEYINPUT5), .ZN(new_n398));
  AOI211_X1 g197(.A(KEYINPUT79), .B(new_n381), .C1(new_n383), .C2(new_n384), .ZN(new_n399));
  OAI22_X1  g198(.A1(new_n398), .A2(new_n399), .B1(new_n376), .B2(new_n371), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(new_n356), .A3(new_n395), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT6), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n397), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(new_n395), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n404), .A2(KEYINPUT6), .A3(new_n357), .ZN(new_n405));
  NAND2_X1  g204(.A1(G226gat), .A2(G233gat), .ZN(new_n406));
  OR2_X1    g205(.A1(new_n261), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n292), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n406), .B1(new_n261), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n318), .A2(new_n315), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n406), .B1(new_n261), .B2(KEYINPUT29), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n407), .A2(new_n415), .A3(KEYINPUT75), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n261), .A2(KEYINPUT75), .A3(new_n406), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n412), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT30), .ZN(new_n421));
  XOR2_X1   g220(.A(G8gat), .B(G36gat), .Z(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(KEYINPUT76), .ZN(new_n423));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n420), .A2(new_n421), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n425), .B1(new_n414), .B2(new_n419), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n261), .A2(new_n406), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT75), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n417), .B1(new_n431), .B2(new_n415), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n413), .B(new_n426), .C1(new_n432), .C2(new_n412), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n428), .A2(KEYINPUT30), .A3(new_n433), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n403), .A2(new_n405), .B1(new_n427), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n351), .A2(new_n436), .A3(KEYINPUT35), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT71), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n273), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT71), .B1(new_n271), .B2(new_n272), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(new_n349), .A3(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n435), .A2(new_n291), .A3(new_n348), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT35), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT86), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT86), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n442), .A2(new_n445), .A3(KEYINPUT35), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n437), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT37), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n448), .B(new_n413), .C1(new_n432), .C2(new_n412), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n449), .A2(new_n425), .ZN(new_n450));
  OR2_X1    g249(.A1(new_n432), .A2(new_n411), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n448), .B1(new_n410), .B2(new_n411), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT38), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n450), .A2(new_n453), .B1(new_n420), .B2(new_n426), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n420), .A2(new_n448), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n449), .A2(new_n425), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT38), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n454), .A2(new_n457), .A3(new_n405), .A4(new_n403), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n393), .B(new_n394), .C1(new_n370), .C2(new_n366), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT39), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n460), .A3(new_n384), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n459), .A2(new_n384), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT39), .B1(new_n383), .B2(new_n384), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n356), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT40), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n464), .A2(new_n465), .B1(new_n404), .B2(new_n357), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n466), .A2(new_n467), .A3(new_n427), .A4(new_n434), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n458), .A2(new_n468), .A3(new_n348), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT36), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n291), .A2(new_n470), .A3(new_n350), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n291), .A2(new_n441), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n469), .B(new_n471), .C1(new_n472), .C2(new_n470), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n435), .A2(new_n348), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n447), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(G15gat), .B(G22gat), .ZN(new_n477));
  OR2_X1    g276(.A1(new_n477), .A2(G1gat), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT16), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n477), .B1(new_n479), .B2(G1gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(G8gat), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT90), .B1(new_n477), .B2(G1gat), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n478), .B(new_n480), .C1(KEYINPUT90), .C2(G8gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G43gat), .B(G50gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT15), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT88), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT14), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(G29gat), .B2(G36gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(G29gat), .A2(G36gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT14), .ZN(new_n493));
  NAND2_X1  g292(.A1(G29gat), .A2(G36gat), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT89), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(KEYINPUT89), .A2(G29gat), .A3(G36gat), .ZN(new_n497));
  AND4_X1   g296(.A1(new_n491), .A2(new_n493), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n487), .A2(KEYINPUT15), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT88), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n487), .A2(new_n500), .A3(KEYINPUT15), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n489), .A2(new_n498), .A3(new_n499), .A4(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n493), .A2(new_n494), .A3(new_n491), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n503), .A2(KEYINPUT15), .A3(new_n487), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT17), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n505), .B1(new_n502), .B2(new_n504), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n486), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G229gat), .A2(G233gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n502), .A2(new_n504), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(new_n485), .A3(new_n484), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT18), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n486), .A2(new_n504), .A3(new_n502), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n511), .ZN(new_n516));
  XOR2_X1   g315(.A(new_n509), .B(KEYINPUT13), .Z(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n508), .A2(KEYINPUT18), .A3(new_n509), .A4(new_n511), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n514), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G113gat), .B(G141gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(G169gat), .B(G197gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT12), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n520), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n514), .A2(new_n518), .A3(new_n519), .A4(new_n526), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n476), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(G57gat), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n533), .A2(G64gat), .ZN(new_n534));
  INV_X1    g333(.A(G64gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n535), .A2(G57gat), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT9), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OR2_X1    g336(.A1(G71gat), .A2(G78gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(G71gat), .A2(G78gat), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT91), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(new_n533), .B2(G64gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n535), .A2(KEYINPUT91), .A3(G57gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n533), .A2(G64gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT9), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n539), .B1(new_n538), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n537), .A2(new_n540), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT92), .B(KEYINPUT21), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(G127gat), .B(G155gat), .Z(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n484), .A2(new_n485), .B1(KEYINPUT21), .B2(new_n548), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n553), .B(new_n554), .Z(new_n555));
  NAND2_X1  g354(.A1(G231gat), .A2(G233gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT93), .ZN(new_n557));
  XOR2_X1   g356(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G183gat), .B(G211gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n555), .B(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT94), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT7), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT7), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT94), .ZN(new_n567));
  AND2_X1   g366(.A1(G85gat), .A2(G92gat), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(G92gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT95), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT95), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(G92gat), .ZN(new_n573));
  INV_X1    g372(.A(G85gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G99gat), .A2(G106gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT8), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n564), .A2(KEYINPUT7), .ZN(new_n578));
  NAND2_X1  g377(.A1(G85gat), .A2(G92gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n569), .A2(new_n575), .A3(new_n577), .A4(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G99gat), .B(G106gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n578), .A2(new_n579), .B1(KEYINPUT8), .B2(new_n576), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n585), .A2(new_n582), .A3(new_n569), .A4(new_n575), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n587), .B1(new_n506), .B2(new_n507), .ZN(new_n588));
  INV_X1    g387(.A(new_n587), .ZN(new_n589));
  AND2_X1   g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n589), .A2(new_n510), .B1(KEYINPUT41), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n595), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n588), .A2(new_n597), .A3(new_n591), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n600));
  XNOR2_X1  g399(.A(G134gat), .B(G162gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n596), .A2(new_n602), .A3(new_n598), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n563), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT98), .ZN(new_n610));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n587), .A2(new_n549), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n584), .A2(new_n548), .A3(new_n586), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(G230gat), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(new_n268), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT10), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n614), .A2(new_n621), .A3(new_n615), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n584), .A2(new_n548), .A3(new_n586), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT10), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n618), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n613), .B1(new_n620), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n548), .B1(new_n584), .B2(new_n586), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n623), .A2(new_n627), .A3(KEYINPUT10), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n615), .A2(new_n621), .ZN(new_n629));
  OAI22_X1  g428(.A1(new_n628), .A2(new_n629), .B1(new_n617), .B2(new_n268), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n630), .A2(new_n619), .A3(new_n612), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n608), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n532), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n403), .A2(new_n405), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT99), .B(G1gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(G1324gat));
  NAND2_X1  g439(.A1(new_n434), .A2(new_n427), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n636), .A2(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n642), .A2(KEYINPUT100), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(KEYINPUT100), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(G8gat), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT16), .B(G8gat), .Z(new_n646));
  NAND3_X1  g445(.A1(new_n642), .A2(KEYINPUT42), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n646), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n648), .B1(new_n643), .B2(new_n644), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n645), .B(new_n647), .C1(new_n649), .C2(KEYINPUT42), .ZN(G1325gat));
  AOI21_X1  g449(.A(new_n470), .B1(new_n291), .B2(new_n441), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n291), .A2(new_n350), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n651), .B1(new_n470), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(G15gat), .B1(new_n636), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n652), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n655), .A2(G15gat), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n654), .B1(new_n636), .B2(new_n656), .ZN(G1326gat));
  NOR2_X1   g456(.A1(new_n636), .A2(new_n348), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT43), .B(G22gat), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1327gat));
  INV_X1    g459(.A(KEYINPUT45), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n562), .A2(new_n632), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n607), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT101), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n532), .A2(new_n664), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n665), .A2(G29gat), .A3(new_n637), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n661), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n670), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n672), .A2(KEYINPUT45), .A3(new_n668), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n606), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n675), .B1(new_n447), .B2(new_n475), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n531), .A2(new_n562), .A3(new_n632), .ZN(new_n677));
  OR3_X1    g476(.A1(new_n351), .A2(new_n436), .A3(KEYINPUT35), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n442), .A2(new_n445), .A3(KEYINPUT35), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n445), .B1(new_n442), .B2(KEYINPUT35), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n474), .A2(KEYINPUT103), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n683), .B1(new_n435), .B2(new_n348), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n653), .A2(new_n469), .A3(new_n682), .A4(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n606), .B1(new_n681), .B2(new_n685), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n676), .B(new_n677), .C1(new_n686), .C2(KEYINPUT44), .ZN(new_n687));
  OAI21_X1  g486(.A(G29gat), .B1(new_n687), .B2(new_n637), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n671), .A2(new_n673), .A3(new_n688), .ZN(G1328gat));
  INV_X1    g488(.A(KEYINPUT46), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n665), .A2(G36gat), .A3(new_n641), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n691), .A2(new_n692), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n690), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n695), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n697), .A2(KEYINPUT46), .A3(new_n693), .ZN(new_n698));
  OAI21_X1  g497(.A(G36gat), .B1(new_n687), .B2(new_n641), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n696), .A2(new_n698), .A3(new_n699), .ZN(G1329gat));
  OR3_X1    g499(.A1(new_n665), .A2(G43gat), .A3(new_n655), .ZN(new_n701));
  OAI21_X1  g500(.A(G43gat), .B1(new_n687), .B2(new_n653), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT105), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n703), .B(new_n705), .ZN(G1330gat));
  OAI21_X1  g505(.A(G50gat), .B1(new_n687), .B2(new_n348), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n348), .A2(G50gat), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n707), .B1(new_n665), .B2(new_n708), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT48), .Z(G1331gat));
  NAND3_X1  g509(.A1(new_n608), .A2(new_n531), .A3(new_n632), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n681), .B2(new_n685), .ZN(new_n712));
  INV_X1    g511(.A(new_n637), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(G57gat), .ZN(G1332gat));
  INV_X1    g514(.A(new_n641), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT49), .B(G64gat), .Z(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n717), .B2(new_n719), .ZN(G1333gat));
  INV_X1    g519(.A(new_n653), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n280), .B1(new_n712), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n655), .A2(G71gat), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n722), .B1(new_n712), .B2(new_n723), .ZN(new_n724));
  XOR2_X1   g523(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1334gat));
  INV_X1    g525(.A(new_n348), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g528(.A1(new_n562), .A2(new_n530), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n682), .A2(new_n684), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n473), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n607), .B(new_n730), .C1(new_n447), .C2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT51), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n686), .A2(KEYINPUT51), .A3(new_n730), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n737), .A2(new_n574), .A3(new_n713), .A4(new_n632), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n530), .A2(new_n562), .A3(new_n633), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n676), .B(new_n739), .C1(new_n686), .C2(KEYINPUT44), .ZN(new_n740));
  OAI21_X1  g539(.A(G85gat), .B1(new_n740), .B2(new_n637), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n741), .ZN(G1336gat));
  NOR2_X1   g541(.A1(new_n740), .A2(new_n641), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n743), .A2(KEYINPUT109), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n571), .A2(new_n573), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(KEYINPUT109), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n737), .A2(new_n570), .A3(new_n716), .A4(new_n632), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n751));
  INV_X1    g550(.A(new_n745), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n743), .B2(new_n752), .ZN(new_n753));
  OAI211_X1 g552(.A(KEYINPUT108), .B(new_n745), .C1(new_n740), .C2(new_n641), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n753), .A2(new_n754), .A3(new_n749), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n750), .B1(new_n748), .B2(new_n755), .ZN(G1337gat));
  OR2_X1    g555(.A1(new_n740), .A2(new_n653), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n282), .B1(new_n757), .B2(KEYINPUT110), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(KEYINPUT110), .B2(new_n757), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n737), .A2(new_n282), .A3(new_n652), .A4(new_n632), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(G1338gat));
  NOR3_X1   g560(.A1(new_n348), .A2(G106gat), .A3(new_n633), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT53), .B1(new_n737), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n740), .A2(new_n348), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n764), .A2(KEYINPUT114), .ZN(new_n765));
  OAI21_X1  g564(.A(G106gat), .B1(new_n764), .B2(KEYINPUT114), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n763), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768));
  OAI21_X1  g567(.A(G106gat), .B1(new_n740), .B2(new_n348), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n762), .B(KEYINPUT111), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n735), .B2(new_n736), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n769), .B1(KEYINPUT112), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n733), .A2(new_n734), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT51), .B1(new_n686), .B2(new_n730), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n770), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n768), .B(KEYINPUT53), .C1(new_n773), .C2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n776), .A2(new_n777), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n772), .A2(KEYINPUT112), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(new_n782), .A3(new_n769), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n768), .B1(new_n783), .B2(KEYINPUT53), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n767), .B1(new_n780), .B2(new_n784), .ZN(G1339gat));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n622), .A2(new_n624), .A3(new_n618), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT115), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n622), .A2(new_n789), .A3(new_n624), .A4(new_n618), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n788), .A2(KEYINPUT54), .A3(new_n630), .A4(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n612), .B1(new_n625), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n791), .A2(KEYINPUT55), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n631), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT55), .B1(new_n791), .B2(new_n793), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n786), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n791), .A2(new_n793), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n800), .A2(KEYINPUT116), .A3(new_n631), .A4(new_n794), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n797), .A2(new_n530), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n517), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n515), .A2(new_n511), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT117), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n515), .A2(new_n511), .A3(new_n806), .A4(new_n803), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n509), .B1(new_n508), .B2(new_n511), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n525), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n810), .A2(new_n529), .A3(new_n632), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n607), .B1(new_n802), .B2(new_n811), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n607), .A2(new_n529), .A3(new_n810), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n813), .A2(new_n797), .A3(new_n801), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n563), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n634), .A2(new_n530), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n815), .A2(KEYINPUT118), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT118), .B1(new_n815), .B2(new_n817), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n637), .A2(new_n716), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n351), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(G113gat), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n825), .A2(new_n826), .A3(new_n531), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n472), .A2(new_n348), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n823), .A2(new_n828), .A3(new_n530), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n827), .B1(new_n826), .B2(new_n829), .ZN(G1340gat));
  OAI21_X1  g629(.A(G120gat), .B1(new_n825), .B2(new_n633), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(KEYINPUT119), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n823), .A2(new_n828), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n633), .A2(G120gat), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(G1341gat));
  OAI21_X1  g634(.A(G127gat), .B1(new_n825), .B2(new_n563), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n562), .A2(new_n247), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n833), .B2(new_n837), .ZN(G1342gat));
  NAND2_X1  g637(.A1(new_n244), .A2(new_n245), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n833), .A2(new_n839), .A3(new_n606), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n841), .A2(KEYINPUT56), .ZN(new_n842));
  OAI21_X1  g641(.A(G134gat), .B1(new_n825), .B2(new_n606), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(KEYINPUT56), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(G1343gat));
  NAND2_X1  g644(.A1(new_n653), .A2(new_n727), .ZN(new_n846));
  NOR4_X1   g645(.A1(new_n822), .A2(G141gat), .A3(new_n531), .A4(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(KEYINPUT58), .ZN(new_n848));
  INV_X1    g647(.A(G141gat), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n727), .A2(KEYINPUT57), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n800), .A2(new_n631), .A3(new_n794), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n851), .A2(new_n531), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT121), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n811), .B(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n607), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n563), .B1(new_n855), .B2(new_n814), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n816), .B1(new_n856), .B2(KEYINPUT122), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n858), .B(new_n563), .C1(new_n855), .C2(new_n814), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n850), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n815), .A2(new_n817), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n815), .A2(new_n817), .A3(KEYINPUT118), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n727), .A3(new_n864), .ZN(new_n865));
  XNOR2_X1  g664(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n860), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n653), .A2(new_n821), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n867), .A2(new_n531), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n848), .B1(new_n849), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n860), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n818), .A2(new_n819), .A3(new_n348), .ZN(new_n872));
  INV_X1    g671(.A(new_n866), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n868), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(KEYINPUT123), .A3(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT123), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n867), .B2(new_n868), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n878), .A3(new_n530), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n847), .B1(new_n879), .B2(G141gat), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT58), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n870), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n870), .B(KEYINPUT124), .C1(new_n880), .C2(new_n881), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1344gat));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n822), .A2(new_n846), .ZN(new_n888));
  AOI211_X1 g687(.A(new_n887), .B(G148gat), .C1(new_n888), .C2(new_n632), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n876), .A2(new_n878), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n887), .B1(new_n890), .B2(new_n633), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n811), .B(KEYINPUT121), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n851), .A2(new_n531), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n606), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n813), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n895), .B2(new_n851), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n896), .A2(KEYINPUT125), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n562), .B1(new_n896), .B2(KEYINPUT125), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n348), .B1(new_n899), .B2(new_n817), .ZN(new_n900));
  OAI22_X1  g699(.A1(new_n900), .A2(KEYINPUT57), .B1(new_n865), .B2(new_n866), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n901), .A2(KEYINPUT59), .A3(new_n632), .A4(new_n875), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n891), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n889), .B1(new_n903), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g703(.A(G155gat), .B1(new_n890), .B2(new_n563), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n888), .A2(new_n295), .A3(new_n562), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1346gat));
  NOR3_X1   g706(.A1(new_n890), .A2(new_n296), .A3(new_n606), .ZN(new_n908));
  AOI21_X1  g707(.A(G162gat), .B1(new_n888), .B2(new_n607), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(G1347gat));
  NOR2_X1   g709(.A1(new_n713), .A2(new_n641), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n820), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n912), .A2(new_n828), .ZN(new_n913));
  AOI21_X1  g712(.A(G169gat), .B1(new_n913), .B2(new_n530), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n824), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n915), .A2(new_n209), .A3(new_n531), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n914), .A2(new_n916), .ZN(G1348gat));
  NAND3_X1  g716(.A1(new_n913), .A2(new_n210), .A3(new_n632), .ZN(new_n918));
  OAI21_X1  g717(.A(G176gat), .B1(new_n915), .B2(new_n633), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1349gat));
  NOR2_X1   g719(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n913), .A2(new_n237), .A3(new_n562), .ZN(new_n922));
  OAI21_X1  g721(.A(G183gat), .B1(new_n915), .B2(new_n563), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n925));
  XOR2_X1   g724(.A(new_n924), .B(new_n925), .Z(G1350gat));
  OAI21_X1  g725(.A(G190gat), .B1(new_n915), .B2(new_n606), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n927), .A2(KEYINPUT127), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(KEYINPUT127), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(KEYINPUT61), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n913), .A2(new_n218), .A3(new_n607), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n930), .B(new_n931), .C1(KEYINPUT61), .C2(new_n929), .ZN(G1351gat));
  AND2_X1   g731(.A1(new_n653), .A2(new_n911), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n901), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(G197gat), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n531), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n872), .A2(new_n530), .A3(new_n933), .ZN(new_n937));
  AOI22_X1  g736(.A1(new_n934), .A2(new_n936), .B1(new_n935), .B2(new_n937), .ZN(G1352gat));
  NAND2_X1  g737(.A1(new_n872), .A2(new_n933), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n939), .A2(G204gat), .A3(new_n633), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT62), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n934), .A2(new_n632), .ZN(new_n942));
  INV_X1    g741(.A(G204gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(G1353gat));
  AOI21_X1  g743(.A(new_n307), .B1(new_n934), .B2(new_n562), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n945), .A2(KEYINPUT63), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n945), .A2(KEYINPUT63), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n562), .A2(new_n307), .ZN(new_n948));
  OAI22_X1  g747(.A1(new_n946), .A2(new_n947), .B1(new_n939), .B2(new_n948), .ZN(G1354gat));
  AND2_X1   g748(.A1(new_n934), .A2(new_n607), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n607), .A2(new_n308), .ZN(new_n951));
  OAI22_X1  g750(.A1(new_n950), .A2(new_n308), .B1(new_n939), .B2(new_n951), .ZN(G1355gat));
endmodule


