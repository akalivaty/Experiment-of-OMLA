

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U553 ( .A1(n736), .A2(n735), .ZN(n737) );
  OR2_X1 U554 ( .A1(n738), .A2(n524), .ZN(n736) );
  AND2_X1 U555 ( .A1(G2105), .A2(G2104), .ZN(n877) );
  NOR2_X2 U556 ( .A1(n535), .A2(n534), .ZN(G160) );
  XNOR2_X1 U557 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n531) );
  NOR2_X1 U558 ( .A1(G2105), .A2(G2104), .ZN(n530) );
  NOR2_X2 U559 ( .A1(G164), .A2(G1384), .ZN(n771) );
  BUF_X1 U560 ( .A(n536), .Z(n520) );
  NAND2_X1 U561 ( .A1(n694), .A2(n693), .ZN(n696) );
  INV_X1 U562 ( .A(KEYINPUT93), .ZN(n695) );
  XNOR2_X1 U563 ( .A(n527), .B(n526), .ZN(n528) );
  INV_X1 U564 ( .A(KEYINPUT13), .ZN(n570) );
  NOR2_X1 U565 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U566 ( .A1(G651), .A2(G543), .ZN(n645) );
  NOR2_X2 U567 ( .A1(G2104), .A2(n525), .ZN(n537) );
  XNOR2_X2 U568 ( .A(n531), .B(n530), .ZN(n617) );
  XOR2_X1 U569 ( .A(G543), .B(KEYINPUT0), .Z(n521) );
  XOR2_X1 U570 ( .A(n758), .B(KEYINPUT97), .Z(n522) );
  AND2_X1 U571 ( .A1(n1011), .A2(n815), .ZN(n523) );
  XOR2_X2 U572 ( .A(KEYINPUT15), .B(n591), .Z(n992) );
  NAND2_X2 U573 ( .A1(n684), .A2(n771), .ZN(n729) );
  NAND2_X1 U574 ( .A1(G286), .A2(G8), .ZN(n524) );
  NOR2_X1 U575 ( .A1(n729), .A2(n969), .ZN(n686) );
  NOR2_X1 U576 ( .A1(n689), .A2(n1009), .ZN(n697) );
  XNOR2_X1 U577 ( .A(KEYINPUT30), .B(KEYINPUT94), .ZN(n720) );
  XNOR2_X1 U578 ( .A(n721), .B(n720), .ZN(n722) );
  INV_X1 U579 ( .A(KEYINPUT95), .ZN(n743) );
  XNOR2_X1 U580 ( .A(n744), .B(n743), .ZN(n745) );
  NAND2_X1 U581 ( .A1(G8), .A2(n729), .ZN(n765) );
  INV_X1 U582 ( .A(G2105), .ZN(n525) );
  AND2_X1 U583 ( .A1(n525), .A2(G2104), .ZN(n536) );
  NOR2_X1 U584 ( .A1(n803), .A2(n523), .ZN(n804) );
  INV_X1 U585 ( .A(KEYINPUT23), .ZN(n526) );
  NAND2_X1 U586 ( .A1(n805), .A2(n804), .ZN(n818) );
  NAND2_X1 U587 ( .A1(n575), .A2(n574), .ZN(n1009) );
  NAND2_X1 U588 ( .A1(n537), .A2(G125), .ZN(n529) );
  NAND2_X1 U589 ( .A1(G101), .A2(n536), .ZN(n527) );
  NAND2_X1 U590 ( .A1(n529), .A2(n528), .ZN(n535) );
  NAND2_X1 U591 ( .A1(G137), .A2(n617), .ZN(n533) );
  NAND2_X1 U592 ( .A1(G113), .A2(n877), .ZN(n532) );
  NAND2_X1 U593 ( .A1(n533), .A2(n532), .ZN(n534) );
  AND2_X1 U594 ( .A1(G138), .A2(n617), .ZN(n543) );
  NAND2_X1 U595 ( .A1(G102), .A2(n520), .ZN(n541) );
  AND2_X1 U596 ( .A1(G126), .A2(n537), .ZN(n539) );
  AND2_X1 U597 ( .A1(G114), .A2(n877), .ZN(n538) );
  NOR2_X1 U598 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U599 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U600 ( .A1(n543), .A2(n542), .ZN(G164) );
  NAND2_X1 U601 ( .A1(G85), .A2(n645), .ZN(n545) );
  INV_X1 U602 ( .A(G651), .ZN(n546) );
  XNOR2_X1 U603 ( .A(KEYINPUT66), .B(n521), .ZN(n635) );
  NOR2_X2 U604 ( .A1(n546), .A2(n635), .ZN(n648) );
  NAND2_X1 U605 ( .A1(G72), .A2(n648), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n552) );
  NOR2_X1 U607 ( .A1(G543), .A2(n546), .ZN(n548) );
  XNOR2_X1 U608 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n547) );
  XNOR2_X2 U609 ( .A(n548), .B(n547), .ZN(n644) );
  NAND2_X1 U610 ( .A1(G60), .A2(n644), .ZN(n550) );
  NOR2_X2 U611 ( .A1(G651), .A2(n635), .ZN(n652) );
  NAND2_X1 U612 ( .A1(G47), .A2(n652), .ZN(n549) );
  NAND2_X1 U613 ( .A1(n550), .A2(n549), .ZN(n551) );
  OR2_X1 U614 ( .A1(n552), .A2(n551), .ZN(G290) );
  AND2_X1 U615 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U616 ( .A(G57), .ZN(G237) );
  INV_X1 U617 ( .A(G132), .ZN(G219) );
  INV_X1 U618 ( .A(G82), .ZN(G220) );
  NAND2_X1 U619 ( .A1(G89), .A2(n645), .ZN(n553) );
  XOR2_X1 U620 ( .A(KEYINPUT4), .B(n553), .Z(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(KEYINPUT73), .ZN(n556) );
  NAND2_X1 U622 ( .A1(G76), .A2(n648), .ZN(n555) );
  NAND2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(KEYINPUT5), .ZN(n562) );
  NAND2_X1 U625 ( .A1(G63), .A2(n644), .ZN(n559) );
  NAND2_X1 U626 ( .A1(G51), .A2(n652), .ZN(n558) );
  NAND2_X1 U627 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U628 ( .A(KEYINPUT6), .B(n560), .Z(n561) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U631 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U632 ( .A1(G7), .A2(G661), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n564), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U634 ( .A(G223), .ZN(n820) );
  NAND2_X1 U635 ( .A1(n820), .A2(G567), .ZN(n565) );
  XOR2_X1 U636 ( .A(KEYINPUT11), .B(n565), .Z(G234) );
  NAND2_X1 U637 ( .A1(G56), .A2(n644), .ZN(n566) );
  XOR2_X1 U638 ( .A(KEYINPUT14), .B(n566), .Z(n573) );
  NAND2_X1 U639 ( .A1(n645), .A2(G81), .ZN(n567) );
  XNOR2_X1 U640 ( .A(n567), .B(KEYINPUT12), .ZN(n569) );
  NAND2_X1 U641 ( .A1(G68), .A2(n648), .ZN(n568) );
  NAND2_X1 U642 ( .A1(n569), .A2(n568), .ZN(n571) );
  XNOR2_X1 U643 ( .A(n571), .B(n570), .ZN(n572) );
  NOR2_X1 U644 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U645 ( .A1(n652), .A2(G43), .ZN(n574) );
  INV_X1 U646 ( .A(G860), .ZN(n606) );
  OR2_X1 U647 ( .A1(n1009), .A2(n606), .ZN(G153) );
  NAND2_X1 U648 ( .A1(G90), .A2(n645), .ZN(n577) );
  NAND2_X1 U649 ( .A1(G77), .A2(n648), .ZN(n576) );
  NAND2_X1 U650 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U651 ( .A(n578), .B(KEYINPUT9), .ZN(n583) );
  NAND2_X1 U652 ( .A1(G64), .A2(n644), .ZN(n580) );
  NAND2_X1 U653 ( .A1(G52), .A2(n652), .ZN(n579) );
  NAND2_X1 U654 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U655 ( .A(KEYINPUT68), .B(n581), .Z(n582) );
  NAND2_X1 U656 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U657 ( .A(n584), .B(KEYINPUT69), .ZN(G171) );
  INV_X1 U658 ( .A(G171), .ZN(G301) );
  NAND2_X1 U659 ( .A1(G868), .A2(G301), .ZN(n593) );
  NAND2_X1 U660 ( .A1(G66), .A2(n644), .ZN(n586) );
  NAND2_X1 U661 ( .A1(G92), .A2(n645), .ZN(n585) );
  NAND2_X1 U662 ( .A1(n586), .A2(n585), .ZN(n590) );
  NAND2_X1 U663 ( .A1(G79), .A2(n648), .ZN(n588) );
  NAND2_X1 U664 ( .A1(G54), .A2(n652), .ZN(n587) );
  NAND2_X1 U665 ( .A1(n588), .A2(n587), .ZN(n589) );
  OR2_X1 U666 ( .A1(n992), .A2(G868), .ZN(n592) );
  NAND2_X1 U667 ( .A1(n593), .A2(n592), .ZN(G284) );
  NAND2_X1 U668 ( .A1(n648), .A2(G78), .ZN(n594) );
  XNOR2_X1 U669 ( .A(n594), .B(KEYINPUT70), .ZN(n596) );
  NAND2_X1 U670 ( .A1(G91), .A2(n645), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U672 ( .A(KEYINPUT71), .B(n597), .ZN(n602) );
  NAND2_X1 U673 ( .A1(G65), .A2(n644), .ZN(n599) );
  NAND2_X1 U674 ( .A1(G53), .A2(n652), .ZN(n598) );
  NAND2_X1 U675 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U676 ( .A(KEYINPUT72), .B(n600), .Z(n601) );
  NAND2_X1 U677 ( .A1(n602), .A2(n601), .ZN(G299) );
  INV_X1 U678 ( .A(G868), .ZN(n665) );
  XNOR2_X1 U679 ( .A(KEYINPUT74), .B(n665), .ZN(n603) );
  NOR2_X1 U680 ( .A1(G286), .A2(n603), .ZN(n605) );
  NOR2_X1 U681 ( .A1(G868), .A2(G299), .ZN(n604) );
  NOR2_X1 U682 ( .A1(n605), .A2(n604), .ZN(G297) );
  NAND2_X1 U683 ( .A1(n606), .A2(G559), .ZN(n607) );
  NAND2_X1 U684 ( .A1(n607), .A2(n992), .ZN(n608) );
  XNOR2_X1 U685 ( .A(n608), .B(KEYINPUT16), .ZN(n609) );
  XOR2_X1 U686 ( .A(KEYINPUT75), .B(n609), .Z(G148) );
  NOR2_X1 U687 ( .A1(G868), .A2(n1009), .ZN(n612) );
  NAND2_X1 U688 ( .A1(G868), .A2(n992), .ZN(n610) );
  NOR2_X1 U689 ( .A1(G559), .A2(n610), .ZN(n611) );
  NOR2_X1 U690 ( .A1(n612), .A2(n611), .ZN(G282) );
  NAND2_X1 U691 ( .A1(G123), .A2(n537), .ZN(n613) );
  XNOR2_X1 U692 ( .A(n613), .B(KEYINPUT76), .ZN(n614) );
  XNOR2_X1 U693 ( .A(n614), .B(KEYINPUT18), .ZN(n616) );
  NAND2_X1 U694 ( .A1(G99), .A2(n520), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n616), .A2(n615), .ZN(n621) );
  NAND2_X1 U696 ( .A1(G135), .A2(n617), .ZN(n619) );
  NAND2_X1 U697 ( .A1(G111), .A2(n877), .ZN(n618) );
  NAND2_X1 U698 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U699 ( .A1(n621), .A2(n620), .ZN(n918) );
  XNOR2_X1 U700 ( .A(n918), .B(G2096), .ZN(n623) );
  INV_X1 U701 ( .A(G2100), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(G156) );
  NAND2_X1 U703 ( .A1(G559), .A2(n992), .ZN(n624) );
  XNOR2_X1 U704 ( .A(n1009), .B(n624), .ZN(n662) );
  NOR2_X1 U705 ( .A1(n662), .A2(G860), .ZN(n631) );
  NAND2_X1 U706 ( .A1(G67), .A2(n644), .ZN(n626) );
  NAND2_X1 U707 ( .A1(G55), .A2(n652), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U709 ( .A1(G93), .A2(n645), .ZN(n628) );
  NAND2_X1 U710 ( .A1(G80), .A2(n648), .ZN(n627) );
  NAND2_X1 U711 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U712 ( .A1(n630), .A2(n629), .ZN(n664) );
  XNOR2_X1 U713 ( .A(n631), .B(n664), .ZN(G145) );
  NAND2_X1 U714 ( .A1(G49), .A2(n652), .ZN(n633) );
  NAND2_X1 U715 ( .A1(G74), .A2(G651), .ZN(n632) );
  NAND2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U717 ( .A1(n644), .A2(n634), .ZN(n637) );
  NAND2_X1 U718 ( .A1(G87), .A2(n635), .ZN(n636) );
  NAND2_X1 U719 ( .A1(n637), .A2(n636), .ZN(G288) );
  NAND2_X1 U720 ( .A1(G88), .A2(n645), .ZN(n639) );
  NAND2_X1 U721 ( .A1(G75), .A2(n648), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n639), .A2(n638), .ZN(n643) );
  NAND2_X1 U723 ( .A1(G62), .A2(n644), .ZN(n641) );
  NAND2_X1 U724 ( .A1(G50), .A2(n652), .ZN(n640) );
  NAND2_X1 U725 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U726 ( .A1(n643), .A2(n642), .ZN(G166) );
  NAND2_X1 U727 ( .A1(G61), .A2(n644), .ZN(n647) );
  NAND2_X1 U728 ( .A1(G86), .A2(n645), .ZN(n646) );
  NAND2_X1 U729 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U730 ( .A1(n648), .A2(G73), .ZN(n649) );
  XOR2_X1 U731 ( .A(KEYINPUT2), .B(n649), .Z(n650) );
  NOR2_X1 U732 ( .A1(n651), .A2(n650), .ZN(n654) );
  NAND2_X1 U733 ( .A1(n652), .A2(G48), .ZN(n653) );
  NAND2_X1 U734 ( .A1(n654), .A2(n653), .ZN(G305) );
  XNOR2_X1 U735 ( .A(KEYINPUT19), .B(KEYINPUT78), .ZN(n656) );
  XNOR2_X1 U736 ( .A(G288), .B(KEYINPUT77), .ZN(n655) );
  XNOR2_X1 U737 ( .A(n656), .B(n655), .ZN(n659) );
  XNOR2_X1 U738 ( .A(G166), .B(G290), .ZN(n657) );
  XNOR2_X1 U739 ( .A(n657), .B(G299), .ZN(n658) );
  XNOR2_X1 U740 ( .A(n659), .B(n658), .ZN(n661) );
  XNOR2_X1 U741 ( .A(G305), .B(n664), .ZN(n660) );
  XNOR2_X1 U742 ( .A(n661), .B(n660), .ZN(n827) );
  XOR2_X1 U743 ( .A(n662), .B(n827), .Z(n663) );
  NAND2_X1 U744 ( .A1(n663), .A2(G868), .ZN(n667) );
  NAND2_X1 U745 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U746 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U747 ( .A(KEYINPUT79), .B(n668), .ZN(G295) );
  NAND2_X1 U748 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(n669), .Z(n670) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n670), .ZN(n671) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n671), .ZN(n672) );
  NAND2_X1 U752 ( .A1(n672), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U753 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U754 ( .A1(G220), .A2(G219), .ZN(n673) );
  XOR2_X1 U755 ( .A(KEYINPUT22), .B(n673), .Z(n674) );
  NOR2_X1 U756 ( .A1(G218), .A2(n674), .ZN(n675) );
  NAND2_X1 U757 ( .A1(G96), .A2(n675), .ZN(n825) );
  NAND2_X1 U758 ( .A1(G2106), .A2(n825), .ZN(n676) );
  XNOR2_X1 U759 ( .A(n676), .B(KEYINPUT80), .ZN(n680) );
  NAND2_X1 U760 ( .A1(G69), .A2(G120), .ZN(n677) );
  NOR2_X1 U761 ( .A1(G237), .A2(n677), .ZN(n678) );
  NAND2_X1 U762 ( .A1(G108), .A2(n678), .ZN(n826) );
  NAND2_X1 U763 ( .A1(G567), .A2(n826), .ZN(n679) );
  NAND2_X1 U764 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U765 ( .A(KEYINPUT81), .B(n681), .ZN(G319) );
  INV_X1 U766 ( .A(G319), .ZN(n905) );
  NAND2_X1 U767 ( .A1(G661), .A2(G483), .ZN(n682) );
  NOR2_X1 U768 ( .A1(n905), .A2(n682), .ZN(n824) );
  NAND2_X1 U769 ( .A1(n824), .A2(G36), .ZN(G176) );
  XOR2_X1 U770 ( .A(KEYINPUT82), .B(G166), .Z(G303) );
  NAND2_X1 U771 ( .A1(G160), .A2(G40), .ZN(n770) );
  INV_X1 U772 ( .A(n770), .ZN(n684) );
  INV_X1 U773 ( .A(G1996), .ZN(n969) );
  XNOR2_X1 U774 ( .A(KEYINPUT26), .B(KEYINPUT91), .ZN(n685) );
  XNOR2_X1 U775 ( .A(n686), .B(n685), .ZN(n688) );
  NAND2_X1 U776 ( .A1(n729), .A2(G1341), .ZN(n687) );
  NAND2_X1 U777 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U778 ( .A1(n697), .A2(n992), .ZN(n694) );
  XNOR2_X2 U779 ( .A(KEYINPUT89), .B(n729), .ZN(n711) );
  NAND2_X1 U780 ( .A1(G2067), .A2(n711), .ZN(n691) );
  NAND2_X1 U781 ( .A1(G1348), .A2(n729), .ZN(n690) );
  NAND2_X1 U782 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U783 ( .A(n692), .B(KEYINPUT92), .ZN(n693) );
  XNOR2_X1 U784 ( .A(n696), .B(n695), .ZN(n699) );
  OR2_X1 U785 ( .A1(n992), .A2(n697), .ZN(n698) );
  NAND2_X1 U786 ( .A1(n699), .A2(n698), .ZN(n704) );
  NAND2_X1 U787 ( .A1(n711), .A2(G2072), .ZN(n700) );
  XNOR2_X1 U788 ( .A(n700), .B(KEYINPUT27), .ZN(n702) );
  INV_X1 U789 ( .A(G1956), .ZN(n941) );
  NOR2_X1 U790 ( .A1(n941), .A2(n711), .ZN(n701) );
  NOR2_X1 U791 ( .A1(n702), .A2(n701), .ZN(n705) );
  INV_X1 U792 ( .A(G299), .ZN(n991) );
  NAND2_X1 U793 ( .A1(n705), .A2(n991), .ZN(n703) );
  NAND2_X1 U794 ( .A1(n704), .A2(n703), .ZN(n709) );
  NOR2_X1 U795 ( .A1(n705), .A2(n991), .ZN(n707) );
  XOR2_X1 U796 ( .A(KEYINPUT28), .B(KEYINPUT90), .Z(n706) );
  XNOR2_X1 U797 ( .A(n707), .B(n706), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U799 ( .A(n710), .B(KEYINPUT29), .ZN(n717) );
  XOR2_X1 U800 ( .A(G2078), .B(KEYINPUT25), .Z(n971) );
  INV_X1 U801 ( .A(n711), .ZN(n712) );
  NOR2_X1 U802 ( .A1(n971), .A2(n712), .ZN(n715) );
  INV_X1 U803 ( .A(n729), .ZN(n713) );
  NOR2_X1 U804 ( .A1(n713), .A2(G1961), .ZN(n714) );
  NOR2_X1 U805 ( .A1(n715), .A2(n714), .ZN(n723) );
  NOR2_X1 U806 ( .A1(G301), .A2(n723), .ZN(n716) );
  NOR2_X1 U807 ( .A1(n717), .A2(n716), .ZN(n728) );
  NOR2_X1 U808 ( .A1(G1966), .A2(n765), .ZN(n739) );
  NOR2_X1 U809 ( .A1(n729), .A2(G2084), .ZN(n718) );
  XNOR2_X1 U810 ( .A(n718), .B(KEYINPUT88), .ZN(n740) );
  NOR2_X1 U811 ( .A1(n739), .A2(n740), .ZN(n719) );
  NAND2_X1 U812 ( .A1(n719), .A2(G8), .ZN(n721) );
  NOR2_X1 U813 ( .A1(G168), .A2(n722), .ZN(n725) );
  AND2_X1 U814 ( .A1(G301), .A2(n723), .ZN(n724) );
  NOR2_X1 U815 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U816 ( .A(n726), .B(KEYINPUT31), .ZN(n727) );
  NOR2_X1 U817 ( .A1(n728), .A2(n727), .ZN(n738) );
  INV_X1 U818 ( .A(G8), .ZN(n734) );
  NOR2_X1 U819 ( .A1(G1971), .A2(n765), .ZN(n731) );
  NOR2_X1 U820 ( .A1(G2090), .A2(n729), .ZN(n730) );
  NOR2_X1 U821 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U822 ( .A1(n732), .A2(G303), .ZN(n733) );
  OR2_X1 U823 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U824 ( .A(n737), .B(KEYINPUT32), .ZN(n746) );
  NOR2_X1 U825 ( .A1(n739), .A2(n738), .ZN(n742) );
  NAND2_X1 U826 ( .A1(G8), .A2(n740), .ZN(n741) );
  NAND2_X1 U827 ( .A1(n742), .A2(n741), .ZN(n744) );
  NAND2_X1 U828 ( .A1(n746), .A2(n745), .ZN(n761) );
  NOR2_X1 U829 ( .A1(G1976), .A2(G288), .ZN(n995) );
  NOR2_X1 U830 ( .A1(G303), .A2(G1971), .ZN(n1015) );
  NOR2_X1 U831 ( .A1(n995), .A2(n1015), .ZN(n747) );
  NAND2_X1 U832 ( .A1(n761), .A2(n747), .ZN(n748) );
  NAND2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n997) );
  NAND2_X1 U834 ( .A1(n748), .A2(n997), .ZN(n749) );
  XNOR2_X1 U835 ( .A(n749), .B(KEYINPUT96), .ZN(n750) );
  NOR2_X2 U836 ( .A1(n750), .A2(n765), .ZN(n751) );
  XNOR2_X1 U837 ( .A(n751), .B(KEYINPUT64), .ZN(n753) );
  INV_X1 U838 ( .A(KEYINPUT33), .ZN(n752) );
  NAND2_X1 U839 ( .A1(n753), .A2(n752), .ZN(n757) );
  INV_X1 U840 ( .A(n765), .ZN(n754) );
  NAND2_X1 U841 ( .A1(n995), .A2(n754), .ZN(n755) );
  NAND2_X1 U842 ( .A1(n755), .A2(KEYINPUT33), .ZN(n756) );
  NAND2_X1 U843 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U844 ( .A(G1981), .B(G305), .Z(n1003) );
  NAND2_X1 U845 ( .A1(n522), .A2(n1003), .ZN(n769) );
  NOR2_X1 U846 ( .A1(G2090), .A2(G303), .ZN(n759) );
  NAND2_X1 U847 ( .A1(G8), .A2(n759), .ZN(n760) );
  NAND2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n762) );
  AND2_X1 U849 ( .A1(n762), .A2(n765), .ZN(n767) );
  NOR2_X1 U850 ( .A1(G1981), .A2(G305), .ZN(n763) );
  XOR2_X1 U851 ( .A(n763), .B(KEYINPUT24), .Z(n764) );
  NOR2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U853 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U854 ( .A1(n769), .A2(n768), .ZN(n805) );
  NOR2_X1 U855 ( .A1(n771), .A2(n770), .ZN(n815) );
  NAND2_X1 U856 ( .A1(G140), .A2(n617), .ZN(n773) );
  NAND2_X1 U857 ( .A1(G104), .A2(n520), .ZN(n772) );
  NAND2_X1 U858 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U859 ( .A(KEYINPUT34), .B(n774), .ZN(n779) );
  NAND2_X1 U860 ( .A1(G128), .A2(n537), .ZN(n776) );
  NAND2_X1 U861 ( .A1(G116), .A2(n877), .ZN(n775) );
  NAND2_X1 U862 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U863 ( .A(n777), .B(KEYINPUT35), .Z(n778) );
  NOR2_X1 U864 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U865 ( .A(KEYINPUT36), .B(n780), .Z(n781) );
  XNOR2_X1 U866 ( .A(KEYINPUT83), .B(n781), .ZN(n888) );
  XNOR2_X1 U867 ( .A(KEYINPUT37), .B(G2067), .ZN(n813) );
  NOR2_X1 U868 ( .A1(n888), .A2(n813), .ZN(n917) );
  NAND2_X1 U869 ( .A1(n815), .A2(n917), .ZN(n811) );
  NAND2_X1 U870 ( .A1(G129), .A2(n537), .ZN(n783) );
  NAND2_X1 U871 ( .A1(G117), .A2(n877), .ZN(n782) );
  NAND2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U873 ( .A(KEYINPUT85), .B(n784), .Z(n787) );
  NAND2_X1 U874 ( .A1(n520), .A2(G105), .ZN(n785) );
  XOR2_X1 U875 ( .A(KEYINPUT38), .B(n785), .Z(n786) );
  NOR2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U877 ( .A(n788), .B(KEYINPUT86), .ZN(n790) );
  NAND2_X1 U878 ( .A1(G141), .A2(n617), .ZN(n789) );
  NAND2_X1 U879 ( .A1(n790), .A2(n789), .ZN(n872) );
  NAND2_X1 U880 ( .A1(G1996), .A2(n872), .ZN(n791) );
  XNOR2_X1 U881 ( .A(n791), .B(KEYINPUT87), .ZN(n800) );
  NAND2_X1 U882 ( .A1(G131), .A2(n617), .ZN(n793) );
  NAND2_X1 U883 ( .A1(G95), .A2(n520), .ZN(n792) );
  NAND2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n796) );
  NAND2_X1 U885 ( .A1(n537), .A2(G119), .ZN(n794) );
  XOR2_X1 U886 ( .A(KEYINPUT84), .B(n794), .Z(n795) );
  NOR2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n798) );
  NAND2_X1 U888 ( .A1(n877), .A2(G107), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n860) );
  AND2_X1 U890 ( .A1(G1991), .A2(n860), .ZN(n799) );
  NOR2_X1 U891 ( .A1(n800), .A2(n799), .ZN(n932) );
  INV_X1 U892 ( .A(n815), .ZN(n801) );
  NOR2_X1 U893 ( .A1(n932), .A2(n801), .ZN(n808) );
  INV_X1 U894 ( .A(n808), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n811), .A2(n802), .ZN(n803) );
  XNOR2_X1 U896 ( .A(G1986), .B(G290), .ZN(n1011) );
  NOR2_X1 U897 ( .A1(G1996), .A2(n872), .ZN(n928) );
  NOR2_X1 U898 ( .A1(G1991), .A2(n860), .ZN(n919) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n806) );
  NOR2_X1 U900 ( .A1(n919), .A2(n806), .ZN(n807) );
  NOR2_X1 U901 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U902 ( .A1(n928), .A2(n809), .ZN(n810) );
  XNOR2_X1 U903 ( .A(n810), .B(KEYINPUT39), .ZN(n812) );
  NAND2_X1 U904 ( .A1(n812), .A2(n811), .ZN(n814) );
  NAND2_X1 U905 ( .A1(n888), .A2(n813), .ZN(n922) );
  NAND2_X1 U906 ( .A1(n814), .A2(n922), .ZN(n816) );
  NAND2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U908 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U909 ( .A(KEYINPUT40), .B(n819), .ZN(G329) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n820), .ZN(G217) );
  NAND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n821) );
  XNOR2_X1 U912 ( .A(KEYINPUT101), .B(n821), .ZN(n822) );
  NAND2_X1 U913 ( .A1(n822), .A2(G661), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U915 ( .A1(n824), .A2(n823), .ZN(G188) );
  INV_X1 U917 ( .A(G120), .ZN(G236) );
  INV_X1 U918 ( .A(G96), .ZN(G221) );
  INV_X1 U919 ( .A(G69), .ZN(G235) );
  NOR2_X1 U920 ( .A1(n826), .A2(n825), .ZN(G325) );
  INV_X1 U921 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U922 ( .A(n1009), .B(n827), .ZN(n829) );
  XNOR2_X1 U923 ( .A(G171), .B(n992), .ZN(n828) );
  XNOR2_X1 U924 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U925 ( .A(G286), .B(n830), .Z(n831) );
  NOR2_X1 U926 ( .A1(G37), .A2(n831), .ZN(G397) );
  XOR2_X1 U927 ( .A(KEYINPUT104), .B(G1976), .Z(n833) );
  XNOR2_X1 U928 ( .A(G1986), .B(G1956), .ZN(n832) );
  XNOR2_X1 U929 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U930 ( .A(n834), .B(KEYINPUT105), .Z(n836) );
  XNOR2_X1 U931 ( .A(G1996), .B(G1991), .ZN(n835) );
  XNOR2_X1 U932 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U933 ( .A(G1981), .B(G1971), .Z(n838) );
  XNOR2_X1 U934 ( .A(G1966), .B(G1961), .ZN(n837) );
  XNOR2_X1 U935 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U936 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U937 ( .A(G2474), .B(KEYINPUT41), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(G229) );
  XOR2_X1 U939 ( .A(G2100), .B(KEYINPUT103), .Z(n844) );
  XNOR2_X1 U940 ( .A(G2678), .B(KEYINPUT43), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U942 ( .A(KEYINPUT42), .B(G2090), .Z(n846) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2072), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U945 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U946 ( .A(KEYINPUT102), .B(G2096), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(n852) );
  XOR2_X1 U948 ( .A(G2078), .B(G2084), .Z(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(G227) );
  NAND2_X1 U950 ( .A1(G124), .A2(n537), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U952 ( .A1(n520), .A2(G100), .ZN(n854) );
  NAND2_X1 U953 ( .A1(n855), .A2(n854), .ZN(n859) );
  NAND2_X1 U954 ( .A1(G136), .A2(n617), .ZN(n857) );
  NAND2_X1 U955 ( .A1(G112), .A2(n877), .ZN(n856) );
  NAND2_X1 U956 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U957 ( .A1(n859), .A2(n858), .ZN(G162) );
  XOR2_X1 U958 ( .A(n918), .B(G162), .Z(n862) );
  XOR2_X1 U959 ( .A(G160), .B(n860), .Z(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U961 ( .A(G164), .B(n863), .ZN(n876) );
  XNOR2_X1 U962 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n874) );
  NAND2_X1 U963 ( .A1(G127), .A2(n537), .ZN(n865) );
  NAND2_X1 U964 ( .A1(G115), .A2(n877), .ZN(n864) );
  NAND2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n866), .B(KEYINPUT47), .ZN(n868) );
  NAND2_X1 U967 ( .A1(G103), .A2(n536), .ZN(n867) );
  NAND2_X1 U968 ( .A1(n868), .A2(n867), .ZN(n871) );
  NAND2_X1 U969 ( .A1(G139), .A2(n617), .ZN(n869) );
  XNOR2_X1 U970 ( .A(KEYINPUT107), .B(n869), .ZN(n870) );
  NOR2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n910) );
  XNOR2_X1 U972 ( .A(n872), .B(n910), .ZN(n873) );
  XNOR2_X1 U973 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n876), .B(n875), .ZN(n887) );
  NAND2_X1 U975 ( .A1(G130), .A2(n537), .ZN(n879) );
  NAND2_X1 U976 ( .A1(G118), .A2(n877), .ZN(n878) );
  NAND2_X1 U977 ( .A1(n879), .A2(n878), .ZN(n885) );
  NAND2_X1 U978 ( .A1(n617), .A2(G142), .ZN(n880) );
  XNOR2_X1 U979 ( .A(n880), .B(KEYINPUT106), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G106), .A2(n536), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U982 ( .A(n883), .B(KEYINPUT45), .Z(n884) );
  NOR2_X1 U983 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U984 ( .A(n887), .B(n886), .Z(n889) );
  XOR2_X1 U985 ( .A(n889), .B(n888), .Z(n890) );
  NOR2_X1 U986 ( .A1(G37), .A2(n890), .ZN(G395) );
  XNOR2_X1 U987 ( .A(G2443), .B(G2446), .ZN(n900) );
  XOR2_X1 U988 ( .A(G2430), .B(KEYINPUT99), .Z(n892) );
  XNOR2_X1 U989 ( .A(G2454), .B(G2435), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n896) );
  XOR2_X1 U991 ( .A(G2438), .B(G2427), .Z(n894) );
  XNOR2_X1 U992 ( .A(G1341), .B(G1348), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U994 ( .A(n896), .B(n895), .Z(n898) );
  XNOR2_X1 U995 ( .A(G2451), .B(KEYINPUT98), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n901) );
  NAND2_X1 U998 ( .A1(n901), .A2(G14), .ZN(n902) );
  XOR2_X1 U999 ( .A(KEYINPUT100), .B(n902), .Z(G401) );
  NOR2_X1 U1000 ( .A1(G229), .A2(G227), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(KEYINPUT49), .B(n903), .ZN(n904) );
  NOR2_X1 U1002 ( .A1(G397), .A2(n904), .ZN(n909) );
  NOR2_X1 U1003 ( .A1(n905), .A2(G401), .ZN(n906) );
  XOR2_X1 U1004 ( .A(KEYINPUT108), .B(n906), .Z(n907) );
  NOR2_X1 U1005 ( .A1(G395), .A2(n907), .ZN(n908) );
  NAND2_X1 U1006 ( .A1(n909), .A2(n908), .ZN(G225) );
  INV_X1 U1007 ( .A(G225), .ZN(G308) );
  INV_X1 U1008 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1009 ( .A(G2072), .B(n910), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(G164), .B(G2078), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(n911), .B(KEYINPUT110), .ZN(n912) );
  NAND2_X1 U1012 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(n914), .B(KEYINPUT111), .ZN(n915) );
  XOR2_X1 U1014 ( .A(KEYINPUT50), .B(n915), .Z(n916) );
  NOR2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(n926) );
  NOR2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1017 ( .A(KEYINPUT109), .B(n920), .Z(n921) );
  NAND2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(n924) );
  XOR2_X1 U1019 ( .A(G160), .B(G2084), .Z(n923) );
  NOR2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n931) );
  XOR2_X1 U1022 ( .A(G2090), .B(G162), .Z(n927) );
  NOR2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1024 ( .A(KEYINPUT51), .B(n929), .ZN(n930) );
  NOR2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n933) );
  NAND2_X1 U1026 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1027 ( .A(n934), .B(KEYINPUT112), .ZN(n935) );
  XNOR2_X1 U1028 ( .A(n935), .B(KEYINPUT52), .ZN(n936) );
  NOR2_X1 U1029 ( .A1(KEYINPUT55), .A2(n936), .ZN(n937) );
  XNOR2_X1 U1030 ( .A(KEYINPUT113), .B(n937), .ZN(n938) );
  NAND2_X1 U1031 ( .A1(n938), .A2(G29), .ZN(n1026) );
  XOR2_X1 U1032 ( .A(G4), .B(KEYINPUT122), .Z(n940) );
  XNOR2_X1 U1033 ( .A(G1348), .B(KEYINPUT59), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(n940), .B(n939), .ZN(n947) );
  XNOR2_X1 U1035 ( .A(G20), .B(n941), .ZN(n945) );
  XNOR2_X1 U1036 ( .A(G1341), .B(G19), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(G1981), .B(G6), .ZN(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1041 ( .A(KEYINPUT123), .B(n948), .Z(n949) );
  XNOR2_X1 U1042 ( .A(KEYINPUT60), .B(n949), .ZN(n963) );
  XNOR2_X1 U1043 ( .A(G1961), .B(G5), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(n950), .B(KEYINPUT121), .ZN(n958) );
  XNOR2_X1 U1045 ( .A(G1971), .B(G22), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G23), .B(G1976), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(G1986), .B(KEYINPUT125), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(n953), .B(G24), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1051 ( .A(KEYINPUT58), .B(n956), .Z(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(G21), .B(G1966), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(KEYINPUT124), .B(n959), .ZN(n960) );
  NOR2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(n964), .B(KEYINPUT61), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(n965), .B(KEYINPUT126), .ZN(n966) );
  NOR2_X1 U1059 ( .A1(G16), .A2(n966), .ZN(n989) );
  XOR2_X1 U1060 ( .A(KEYINPUT55), .B(KEYINPUT115), .Z(n986) );
  XNOR2_X1 U1061 ( .A(G2090), .B(G35), .ZN(n981) );
  XNOR2_X1 U1062 ( .A(G2067), .B(G26), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(G33), .B(G2072), .ZN(n967) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n976) );
  XNOR2_X1 U1065 ( .A(G32), .B(n969), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n970), .A2(G28), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(G27), .B(n971), .ZN(n972) );
  XNOR2_X1 U1068 ( .A(KEYINPUT114), .B(n972), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(G25), .B(G1991), .ZN(n977) );
  NOR2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(KEYINPUT53), .B(n979), .ZN(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n984) );
  XOR2_X1 U1075 ( .A(G2084), .B(G34), .Z(n982) );
  XNOR2_X1 U1076 ( .A(KEYINPUT54), .B(n982), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(n986), .B(n985), .ZN(n987) );
  NOR2_X1 U1079 ( .A1(G29), .A2(n987), .ZN(n988) );
  NOR2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(G11), .A2(n990), .ZN(n1023) );
  XNOR2_X1 U1082 ( .A(G16), .B(KEYINPUT56), .ZN(n1020) );
  XNOR2_X1 U1083 ( .A(n991), .B(G1956), .ZN(n1002) );
  XNOR2_X1 U1084 ( .A(n992), .B(G1348), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(G1971), .A2(G303), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n1000) );
  XOR2_X1 U1087 ( .A(n995), .B(KEYINPUT118), .Z(n996) );
  NAND2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1089 ( .A(KEYINPUT119), .B(n998), .Z(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1008) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G168), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(n1005), .B(KEYINPUT57), .ZN(n1006) );
  XOR2_X1 U1095 ( .A(KEYINPUT116), .B(n1006), .Z(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1018) );
  XNOR2_X1 U1097 ( .A(G1341), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(G1961), .B(KEYINPUT117), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(n1012), .B(G301), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1105 ( .A(KEYINPUT120), .B(n1021), .Z(n1022) );
  NOR2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1107 ( .A(KEYINPUT127), .B(n1024), .Z(n1025) );
  NAND2_X1 U1108 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1027), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

