//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n596,
    new_n597, new_n598, new_n599, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n645, new_n646, new_n649, new_n651, new_n652, new_n653, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160,
    new_n1161, new_n1163, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT65), .B(G2105), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n468), .A2(new_n469), .B1(G101), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n473), .B1(new_n466), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n469), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  OAI221_X1 g054(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n469), .C2(G112), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT67), .Z(new_n481));
  NOR2_X1   g056(.A1(new_n466), .A2(G2105), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(G136), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n466), .A2(new_n469), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT66), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n466), .ZN(new_n492));
  AND2_X1   g067(.A1(G126), .A2(G2105), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n492), .A2(KEYINPUT4), .A3(G138), .A4(new_n469), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  OAI21_X1  g071(.A(G138), .B1(new_n464), .B2(new_n465), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n476), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n494), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n501));
  XOR2_X1   g076(.A(KEYINPUT6), .B(G651), .Z(new_n502));
  AND2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n501), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT68), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G88), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n502), .A2(new_n508), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n505), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(G50), .A2(new_n517), .B1(new_n520), .B2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n516), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n515), .A2(G89), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT69), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n528), .B1(new_n503), .B2(new_n504), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n509), .A2(KEYINPUT69), .A3(new_n510), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT70), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT70), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n529), .A2(new_n530), .A3(new_n534), .A4(new_n531), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT71), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n508), .B1(new_n512), .B2(new_n537), .ZN(new_n538));
  OR2_X1    g113(.A1(KEYINPUT6), .A2(G651), .ZN(new_n539));
  NAND2_X1  g114(.A1(KEYINPUT6), .A2(G651), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n539), .A2(KEYINPUT71), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n538), .A2(G51), .A3(new_n541), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n536), .A2(KEYINPUT72), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(KEYINPUT72), .B1(new_n536), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n527), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(G168));
  NAND3_X1  g121(.A1(new_n529), .A2(new_n530), .A3(G64), .ZN(new_n547));
  NAND2_X1  g122(.A1(G77), .A2(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n538), .A2(G52), .A3(new_n541), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n506), .A2(G90), .A3(new_n513), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(KEYINPUT73), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n550), .A2(new_n555), .A3(new_n551), .A4(new_n552), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(G171));
  INV_X1    g132(.A(G81), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n538), .A2(new_n541), .ZN(new_n559));
  INV_X1    g134(.A(G43), .ZN(new_n560));
  OAI22_X1  g135(.A1(new_n514), .A2(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(G651), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n529), .A2(new_n530), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G56), .ZN(new_n564));
  NAND2_X1  g139(.A1(G68), .A2(G543), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  INV_X1    g147(.A(KEYINPUT74), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT68), .ZN(new_n574));
  AOI21_X1  g149(.A(KEYINPUT68), .B1(new_n511), .B2(new_n512), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n506), .A2(KEYINPUT74), .A3(new_n513), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n576), .A2(new_n577), .A3(G91), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n512), .A2(new_n537), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n579), .A2(G53), .A3(G543), .A4(new_n541), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT9), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT9), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n538), .A2(new_n582), .A3(G53), .A4(new_n541), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(G78), .A2(G543), .ZN(new_n585));
  XOR2_X1   g160(.A(KEYINPUT75), .B(G65), .Z(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n586), .B2(new_n505), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n578), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(KEYINPUT76), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT76), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n578), .A2(new_n584), .A3(new_n591), .A4(new_n588), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G299));
  INV_X1    g169(.A(G171), .ZN(G301));
  NAND2_X1  g170(.A1(new_n545), .A2(KEYINPUT77), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT77), .ZN(new_n597));
  OAI211_X1 g172(.A(new_n597), .B(new_n527), .C1(new_n543), .C2(new_n544), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G286));
  AND2_X1   g175(.A1(new_n576), .A2(new_n577), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G87), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n563), .A2(G74), .ZN(new_n603));
  INV_X1    g178(.A(new_n559), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n603), .A2(G651), .B1(new_n604), .B2(G49), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n602), .A2(new_n605), .ZN(G288));
  INV_X1    g181(.A(G61), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT78), .B1(new_n505), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G73), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n508), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT78), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n511), .A2(new_n611), .A3(G61), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(G651), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT79), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n601), .A2(G86), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n517), .A2(G48), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT80), .Z(new_n619));
  NAND3_X1  g194(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(G305));
  INV_X1    g195(.A(G85), .ZN(new_n621));
  INV_X1    g196(.A(G47), .ZN(new_n622));
  OAI22_X1  g197(.A1(new_n514), .A2(new_n621), .B1(new_n559), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n563), .A2(G60), .ZN(new_n624));
  NAND2_X1  g199(.A1(G72), .A2(G543), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n562), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(G290));
  NAND2_X1  g203(.A1(new_n604), .A2(G54), .ZN(new_n629));
  AND2_X1   g204(.A1(new_n511), .A2(G66), .ZN(new_n630));
  NAND2_X1  g205(.A1(G79), .A2(G543), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT82), .Z(new_n632));
  OAI21_X1  g207(.A(G651), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n576), .A2(new_n577), .A3(G92), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g213(.A1(new_n576), .A2(new_n577), .A3(G92), .A4(new_n636), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n634), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(G868), .ZN(new_n642));
  MUX2_X1   g217(.A(G301), .B(new_n641), .S(new_n642), .Z(G284));
  MUX2_X1   g218(.A(G301), .B(new_n641), .S(new_n642), .Z(G321));
  OAI21_X1  g219(.A(KEYINPUT83), .B1(new_n593), .B2(G868), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n599), .A2(new_n642), .ZN(new_n646));
  MUX2_X1   g221(.A(new_n645), .B(KEYINPUT83), .S(new_n646), .Z(G297));
  MUX2_X1   g222(.A(new_n645), .B(KEYINPUT83), .S(new_n646), .Z(G280));
  INV_X1    g223(.A(G559), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n640), .B1(new_n649), .B2(G860), .ZN(G148));
  INV_X1    g225(.A(new_n567), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(new_n642), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n641), .A2(G559), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n652), .B1(new_n653), .B2(new_n642), .ZN(G323));
  XNOR2_X1  g229(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g230(.A1(new_n492), .A2(new_n471), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT13), .Z(new_n659));
  INV_X1    g234(.A(G2100), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  AOI22_X1  g237(.A1(G123), .A2(new_n484), .B1(new_n482), .B2(G135), .ZN(new_n663));
  OAI221_X1 g238(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n469), .C2(G111), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(G2096), .Z(new_n666));
  NAND3_X1  g241(.A1(new_n661), .A2(new_n662), .A3(new_n666), .ZN(G156));
  XNOR2_X1  g242(.A(KEYINPUT15), .B(G2435), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2438), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2427), .B(G2430), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT85), .B(KEYINPUT14), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT86), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(new_n669), .B2(new_n670), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2443), .B(G2446), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1341), .B(G1348), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2451), .B(G2454), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT16), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n681), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(new_n683), .A3(G14), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(KEYINPUT87), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT87), .ZN(new_n686));
  NAND4_X1  g261(.A1(new_n682), .A2(new_n683), .A3(new_n686), .A4(G14), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT88), .ZN(G401));
  XNOR2_X1  g264(.A(G2067), .B(G2678), .ZN(new_n690));
  NOR2_X1   g265(.A1(G2072), .A2(G2078), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n444), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n690), .B1(new_n693), .B2(KEYINPUT89), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(KEYINPUT89), .B2(new_n693), .ZN(new_n695));
  XOR2_X1   g270(.A(G2084), .B(G2090), .Z(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n692), .B(KEYINPUT17), .ZN(new_n698));
  INV_X1    g273(.A(new_n690), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n695), .B(new_n697), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  NOR3_X1   g275(.A1(new_n697), .A2(new_n692), .A3(new_n699), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT18), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n698), .A2(new_n699), .A3(new_n696), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n700), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(new_n660), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT90), .B(G2096), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(G227));
  XOR2_X1   g282(.A(G1971), .B(G1976), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT19), .ZN(new_n709));
  XOR2_X1   g284(.A(G1956), .B(G2474), .Z(new_n710));
  XOR2_X1   g285(.A(G1961), .B(G1966), .Z(new_n711));
  NAND3_X1  g286(.A1(new_n710), .A2(new_n711), .A3(KEYINPUT91), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT91), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n709), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT20), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n710), .A2(new_n711), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n709), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n718), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(new_n713), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n717), .B(new_n719), .C1(new_n709), .C2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(G1991), .B(G1996), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(G1981), .B(G1986), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(G229));
  INV_X1    g303(.A(G29), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n729), .A2(G33), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT25), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G139), .B2(new_n482), .ZN(new_n733));
  NAND2_X1  g308(.A1(G115), .A2(G2104), .ZN(new_n734));
  INV_X1    g309(.A(G127), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n466), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(new_n476), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(KEYINPUT96), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(KEYINPUT96), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n733), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n730), .B1(new_n740), .B2(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(new_n442), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT97), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n729), .A2(G32), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n482), .A2(G141), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT99), .Z(new_n746));
  NAND2_X1  g321(.A1(new_n484), .A2(G129), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT100), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n484), .A2(KEYINPUT100), .A3(G129), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT26), .Z(new_n753));
  NAND2_X1  g328(.A1(new_n471), .A2(G105), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n746), .A2(new_n751), .A3(new_n753), .A4(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n744), .B1(new_n755), .B2(G29), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT27), .B(G1996), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT24), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(G34), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(G34), .ZN(new_n761));
  AOI21_X1  g336(.A(G29), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n478), .B2(G29), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT98), .Z(new_n764));
  INV_X1    g339(.A(G2084), .ZN(new_n765));
  OAI221_X1 g340(.A(new_n758), .B1(new_n442), .B2(new_n741), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n743), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT101), .Z(new_n768));
  OR2_X1    g343(.A1(new_n756), .A2(new_n757), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n729), .A2(G27), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G164), .B2(new_n729), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(new_n443), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT31), .B(G11), .Z(new_n773));
  NOR2_X1   g348(.A1(new_n665), .A2(new_n729), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT30), .B(G28), .ZN(new_n775));
  AOI211_X1 g350(.A(new_n773), .B(new_n774), .C1(new_n729), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n764), .A2(new_n765), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n769), .A2(new_n772), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G16), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G5), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G171), .B2(new_n779), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n778), .B1(G1961), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n779), .A2(G21), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G168), .B2(new_n779), .ZN(new_n784));
  INV_X1    g359(.A(G1966), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n782), .B(new_n786), .C1(G1961), .C2(new_n781), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n768), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(KEYINPUT102), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n484), .A2(G128), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT93), .Z(new_n791));
  INV_X1    g366(.A(G116), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n470), .B1(new_n476), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G104), .A2(G2105), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT94), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n793), .A2(new_n795), .B1(G140), .B2(new_n482), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(G29), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT95), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n729), .A2(G26), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT28), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2067), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n729), .A2(G35), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G162), .B2(new_n729), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT29), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n803), .B1(G2090), .B2(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n806), .A2(G2090), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n779), .A2(G19), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n567), .B2(new_n779), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(G1341), .Z(new_n811));
  NAND3_X1  g386(.A1(new_n807), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n779), .A2(G20), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT23), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n593), .B2(new_n779), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G1956), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n779), .A2(G4), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n640), .B2(new_n779), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G1348), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n812), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n789), .A2(new_n820), .ZN(new_n821));
  AOI22_X1  g396(.A1(G119), .A2(new_n484), .B1(new_n482), .B2(G131), .ZN(new_n822));
  OAI221_X1 g397(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n469), .C2(G107), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  MUX2_X1   g399(.A(G25), .B(new_n824), .S(G29), .Z(new_n825));
  XOR2_X1   g400(.A(KEYINPUT35), .B(G1991), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(KEYINPUT92), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n779), .A2(G24), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n627), .B2(new_n779), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(G1986), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n831), .A2(G1986), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n829), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  MUX2_X1   g409(.A(G6), .B(G305), .S(G16), .Z(new_n835));
  XOR2_X1   g410(.A(KEYINPUT32), .B(G1981), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n779), .A2(G22), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(G166), .B2(new_n779), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G1971), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n779), .A2(G23), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(G288), .B2(G16), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT33), .B(G1976), .Z(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n842), .A2(new_n844), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n840), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n837), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n834), .B1(new_n848), .B2(KEYINPUT34), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(KEYINPUT34), .B2(new_n848), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n828), .A2(KEYINPUT92), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n850), .B(new_n852), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n788), .A2(KEYINPUT102), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n821), .A2(new_n853), .A3(new_n854), .ZN(G311));
  NAND3_X1  g430(.A1(new_n821), .A2(new_n853), .A3(new_n854), .ZN(G150));
  NAND2_X1  g431(.A1(new_n640), .A2(G559), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT38), .Z(new_n858));
  AOI22_X1  g433(.A1(new_n515), .A2(G93), .B1(new_n604), .B2(G55), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n563), .A2(G67), .ZN(new_n860));
  NAND2_X1  g435(.A1(G80), .A2(G543), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n859), .B1(new_n562), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n651), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n858), .B(new_n864), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n865), .A2(KEYINPUT39), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(KEYINPUT39), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n866), .A2(new_n867), .A3(G860), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n863), .A2(G860), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT37), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n868), .A2(new_n870), .ZN(G145));
  INV_X1    g446(.A(KEYINPUT40), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n755), .B(new_n797), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n499), .B(KEYINPUT103), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n740), .B(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n873), .B(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n658), .B(new_n824), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n484), .A2(G130), .ZN(new_n878));
  OAI221_X1 g453(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n469), .C2(G118), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n482), .A2(G142), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n877), .B(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n876), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n665), .B(new_n478), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n487), .B(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n882), .B(new_n883), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n886), .B(new_n888), .C1(new_n889), .C2(new_n876), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n889), .A2(new_n876), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n893), .A2(KEYINPUT105), .A3(new_n888), .A4(new_n886), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n888), .B1(new_n893), .B2(new_n886), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n896), .A2(G37), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n895), .A2(new_n897), .A3(KEYINPUT106), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT106), .B1(new_n895), .B2(new_n897), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n872), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n895), .A2(new_n897), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n895), .A2(new_n897), .A3(KEYINPUT106), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(KEYINPUT40), .A3(new_n904), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n900), .A2(new_n905), .ZN(G395));
  NAND2_X1  g481(.A1(new_n863), .A2(new_n642), .ZN(new_n907));
  XNOR2_X1  g482(.A(G305), .B(new_n627), .ZN(new_n908));
  XNOR2_X1  g483(.A(G288), .B(G166), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n908), .B(new_n909), .Z(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT42), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n864), .B(new_n653), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n640), .A2(new_n590), .A3(new_n592), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n638), .A2(new_n639), .ZN(new_n914));
  INV_X1    g489(.A(new_n634), .ZN(new_n915));
  AOI22_X1  g490(.A1(new_n590), .A2(new_n592), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n917), .B(KEYINPUT41), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n918), .B1(new_n912), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n911), .B(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n907), .B1(new_n921), .B2(new_n642), .ZN(G295));
  OAI21_X1  g497(.A(new_n907), .B1(new_n921), .B2(new_n642), .ZN(G331));
  AOI21_X1  g498(.A(G301), .B1(new_n596), .B2(new_n598), .ZN(new_n924));
  INV_X1    g499(.A(new_n544), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n536), .A2(KEYINPUT72), .A3(new_n542), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(G171), .B1(new_n927), .B2(new_n527), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n864), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT107), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n928), .B1(new_n599), .B2(G171), .ZN(new_n931));
  INV_X1    g506(.A(new_n864), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n917), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n934), .B(new_n864), .C1(new_n924), .C2(new_n928), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n930), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT108), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n930), .A2(new_n933), .A3(new_n938), .A4(new_n935), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n924), .A2(new_n864), .A3(new_n928), .ZN(new_n941));
  INV_X1    g516(.A(new_n929), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n919), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(G37), .B1(new_n944), .B2(new_n910), .ZN(new_n945));
  INV_X1    g520(.A(new_n910), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n940), .A2(new_n946), .A3(new_n943), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT43), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n947), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  INV_X1    g525(.A(G37), .ZN(new_n951));
  INV_X1    g526(.A(new_n941), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(new_n930), .A3(new_n935), .ZN(new_n953));
  AOI22_X1  g528(.A1(new_n953), .A2(new_n919), .B1(new_n929), .B2(new_n933), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n951), .B1(new_n954), .B2(new_n946), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n949), .A2(new_n950), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT44), .B1(new_n948), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n950), .B1(new_n945), .B2(new_n947), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n949), .A2(KEYINPUT43), .A3(new_n955), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n957), .A2(new_n961), .ZN(G397));
  INV_X1    g537(.A(KEYINPUT61), .ZN(new_n963));
  XNOR2_X1  g538(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n589), .B(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n499), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(KEYINPUT50), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n969), .B1(new_n499), .B2(new_n966), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n472), .A2(G40), .A3(new_n477), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT116), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n968), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT116), .B1(new_n970), .B2(new_n971), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g551(.A(KEYINPUT117), .B(G1956), .Z(new_n977));
  AOI21_X1  g552(.A(KEYINPUT118), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(KEYINPUT118), .A3(new_n977), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT111), .B1(new_n967), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n971), .B1(new_n967), .B2(new_n982), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n499), .A2(new_n985), .A3(KEYINPUT45), .A4(new_n966), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n983), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT56), .B(G2072), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n965), .B1(new_n981), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n980), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n965), .B(new_n990), .C1(new_n992), .C2(new_n978), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n963), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n967), .ZN(new_n996));
  INV_X1    g571(.A(new_n971), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT120), .ZN(new_n999));
  OR3_X1    g574(.A1(new_n967), .A2(KEYINPUT120), .A3(new_n971), .ZN(new_n1000));
  AOI21_X1  g575(.A(G2067), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n968), .A2(new_n971), .A3(new_n970), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1002), .A2(G1348), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT60), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1004), .A2(new_n1005), .A3(new_n640), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n651), .A2(KEYINPUT122), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n987), .A2(G1996), .ZN(new_n1008));
  XOR2_X1   g583(.A(KEYINPUT58), .B(G1341), .Z(new_n1009));
  NAND3_X1  g584(.A1(new_n999), .A2(new_n1000), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1007), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1006), .B1(KEYINPUT59), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1004), .A2(new_n641), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n640), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1005), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1011), .A2(KEYINPUT59), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1012), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n990), .B1(new_n992), .B2(new_n978), .ZN(new_n1018));
  INV_X1    g593(.A(new_n965), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1020), .A2(KEYINPUT61), .A3(new_n993), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n995), .A2(new_n1017), .A3(new_n1021), .ZN(new_n1022));
  XOR2_X1   g597(.A(new_n1014), .B(KEYINPUT121), .Z(new_n1023));
  OAI21_X1  g598(.A(new_n993), .B1(new_n1023), .B2(new_n991), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(G305), .B2(G1981), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n617), .A2(new_n619), .ZN(new_n1028));
  INV_X1    g603(.A(G1981), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1028), .A2(KEYINPUT115), .A3(new_n1029), .A4(new_n616), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G86), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n619), .B1(new_n1032), .B2(new_n514), .ZN(new_n1033));
  INV_X1    g608(.A(new_n614), .ZN(new_n1034));
  OAI21_X1  g609(.A(G1981), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT49), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1031), .A2(KEYINPUT49), .A3(new_n1035), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n998), .A2(G8), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n972), .B1(KEYINPUT50), .B2(new_n967), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(G2084), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n996), .A2(KEYINPUT45), .ZN(new_n1045));
  AOI21_X1  g620(.A(G1966), .B1(new_n1045), .B2(new_n984), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n545), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1046), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1048), .B(G168), .C1(G2084), .C2(new_n1043), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1047), .A2(new_n1049), .A3(G8), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT51), .ZN(new_n1051));
  INV_X1    g626(.A(G8), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1046), .B1(new_n765), .B2(new_n1002), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1052), .B1(new_n1053), .B2(G168), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1051), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1976), .ZN(new_n1058));
  NOR2_X1   g633(.A1(G288), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1040), .B1(new_n1059), .B2(KEYINPUT114), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(KEYINPUT114), .B2(new_n1059), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT52), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT52), .B1(G288), .B2(new_n1058), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1060), .B(new_n1063), .C1(KEYINPUT114), .C2(new_n1059), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(G303), .A2(G8), .ZN(new_n1066));
  XOR2_X1   g641(.A(new_n1066), .B(KEYINPUT55), .Z(new_n1067));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n987), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G1971), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n983), .A2(new_n984), .A3(KEYINPUT112), .A4(new_n986), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(G2090), .B2(new_n976), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1067), .B1(new_n1073), .B2(G8), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1042), .A2(new_n1057), .A3(new_n1065), .A4(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1072), .B1(G2090), .B2(new_n1043), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(G8), .A3(new_n1067), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT113), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n1078), .B(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n1081));
  OR2_X1    g656(.A1(KEYINPUT124), .A2(G2078), .ZN(new_n1082));
  NAND2_X1  g657(.A1(KEYINPUT124), .A2(G2078), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G1961), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n988), .A2(new_n1084), .B1(new_n1085), .B2(new_n1043), .ZN(new_n1086));
  AOI21_X1  g661(.A(G2078), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(new_n1087), .B2(KEYINPUT53), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1088), .A2(G171), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1043), .A2(new_n1085), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1045), .A2(new_n984), .A3(KEYINPUT53), .A4(new_n443), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1091), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1094));
  OAI22_X1  g669(.A1(new_n1093), .A2(new_n1094), .B1(new_n1087), .B2(KEYINPUT53), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(G171), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT54), .B1(new_n1089), .B2(new_n1096), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1076), .A2(new_n1080), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1088), .A2(KEYINPUT125), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT125), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1100), .B(new_n1086), .C1(new_n1087), .C2(KEYINPUT53), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1099), .A2(G171), .A3(new_n1101), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n1102), .A2(KEYINPUT126), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(KEYINPUT126), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1095), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(G301), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1103), .A2(KEYINPUT54), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1025), .A2(new_n1098), .A3(new_n1107), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1042), .A2(new_n1065), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1055), .B1(new_n1054), .B2(new_n1047), .ZN(new_n1110));
  AOI211_X1 g685(.A(KEYINPUT51), .B(new_n1052), .C1(new_n1053), .C2(G168), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT62), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1051), .A2(new_n1113), .A3(new_n1056), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1096), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NOR3_X1   g691(.A1(G286), .A2(new_n1053), .A3(new_n1052), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT63), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1074), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1109), .B1(new_n1120), .B2(new_n1080), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1042), .A2(new_n1058), .A3(new_n602), .A4(new_n605), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n1031), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1077), .A2(G8), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1067), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1042), .A2(new_n1065), .A3(new_n1117), .A4(new_n1126), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1123), .A2(new_n1041), .B1(KEYINPUT63), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1108), .A2(new_n1121), .A3(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n797), .B(G2067), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n996), .A2(KEYINPUT45), .A3(new_n971), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1130), .A2(KEYINPUT109), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT109), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1131), .ZN(new_n1134));
  XOR2_X1   g709(.A(new_n755), .B(G1996), .Z(new_n1135));
  OAI22_X1  g710(.A1(new_n1132), .A2(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT110), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n824), .B(new_n826), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1137), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1139));
  XOR2_X1   g714(.A(new_n627), .B(G1986), .Z(new_n1140));
  AOI21_X1  g715(.A(new_n1139), .B1(new_n1131), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1129), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1137), .A2(new_n826), .A3(new_n823), .A4(new_n822), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n797), .A2(G2067), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1134), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT46), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1134), .A2(new_n1146), .A3(G1996), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1131), .B1(new_n1130), .B2(new_n755), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1147), .B1(new_n1148), .B2(KEYINPUT127), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1146), .B1(new_n1134), .B2(G1996), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1149), .B(new_n1150), .C1(KEYINPUT127), .C2(new_n1148), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT47), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1134), .A2(G1986), .A3(G290), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT48), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1152), .B1(new_n1139), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1145), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1142), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g732(.A1(new_n959), .A2(new_n960), .ZN(new_n1159));
  NOR3_X1   g733(.A1(G229), .A2(new_n462), .A3(G227), .ZN(new_n1160));
  OAI211_X1 g734(.A(new_n688), .B(new_n1160), .C1(new_n898), .C2(new_n899), .ZN(new_n1161));
  NOR2_X1   g735(.A1(new_n1159), .A2(new_n1161), .ZN(G308));
  AND2_X1   g736(.A1(new_n688), .A2(new_n1160), .ZN(new_n1163));
  NAND2_X1  g737(.A1(new_n903), .A2(new_n904), .ZN(new_n1164));
  OAI211_X1 g738(.A(new_n1163), .B(new_n1164), .C1(new_n959), .C2(new_n960), .ZN(G225));
endmodule


