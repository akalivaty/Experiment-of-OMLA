//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G116), .B(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT5), .ZN(new_n192));
  INV_X1    g006(.A(G116), .ZN(new_n193));
  NOR3_X1   g007(.A1(new_n193), .A2(KEYINPUT5), .A3(G119), .ZN(new_n194));
  INV_X1    g008(.A(G113), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT2), .B(G113), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n192), .A2(new_n196), .B1(new_n198), .B2(new_n191), .ZN(new_n199));
  INV_X1    g013(.A(G107), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(KEYINPUT80), .A3(G104), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT80), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G107), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n200), .A2(G104), .ZN(new_n205));
  OAI211_X1 g019(.A(G101), .B(new_n201), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT3), .B1(new_n203), .B2(G107), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(new_n200), .A3(G104), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n203), .A2(G107), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n207), .A2(new_n209), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n206), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n199), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n207), .A2(new_n209), .A3(new_n211), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT4), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(G101), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n198), .A2(KEYINPUT66), .A3(new_n191), .ZN(new_n218));
  XOR2_X1   g032(.A(G116), .B(G119), .Z(new_n219));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n197), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n217), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n215), .A2(G101), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n223), .A2(KEYINPUT4), .A3(new_n212), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n214), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G110), .B(G122), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n226), .B(KEYINPUT85), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT85), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n226), .B(new_n229), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n230), .B(new_n214), .C1(new_n222), .C2(new_n224), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n228), .A2(KEYINPUT6), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G143), .ZN(new_n234));
  INV_X1    g048(.A(G143), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G146), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n234), .A2(new_n236), .A3(KEYINPUT0), .A4(G128), .ZN(new_n237));
  XNOR2_X1  g051(.A(G143), .B(G146), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT0), .B(G128), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G125), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT1), .B1(new_n235), .B2(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G128), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n234), .A2(new_n236), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G125), .ZN(new_n246));
  INV_X1    g060(.A(G128), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(KEYINPUT1), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n238), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n245), .A2(new_n246), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n241), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G224), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(G953), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n253), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(new_n241), .B2(new_n250), .ZN(new_n256));
  OR2_X1    g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n225), .A2(new_n258), .A3(new_n227), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n232), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  OAI22_X1  g074(.A1(new_n254), .A2(new_n256), .B1(KEYINPUT7), .B2(new_n253), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n230), .A2(KEYINPUT8), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT8), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n227), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT87), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n206), .A2(new_n212), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n199), .B(new_n266), .C1(KEYINPUT86), .C2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n192), .A2(new_n196), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n269), .B1(new_n197), .B2(new_n219), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n266), .B2(new_n267), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT86), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT87), .B1(new_n213), .B2(new_n272), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n265), .B(new_n268), .C1(new_n271), .C2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT7), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n251), .A2(new_n275), .A3(new_n255), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n261), .A2(new_n231), .A3(new_n274), .A4(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G902), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n190), .B1(new_n260), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n232), .A2(new_n257), .A3(new_n259), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n281), .A2(new_n278), .A3(new_n189), .A4(new_n277), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n188), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT90), .ZN(new_n284));
  INV_X1    g098(.A(G475), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n278), .ZN(new_n286));
  INV_X1    g100(.A(G140), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G125), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n246), .A2(G140), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT89), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT89), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(KEYINPUT19), .A3(new_n293), .ZN(new_n294));
  OR2_X1    g108(.A1(new_n290), .A2(KEYINPUT19), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n233), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT16), .ZN(new_n297));
  OR3_X1    g111(.A1(new_n246), .A2(KEYINPUT16), .A3(G140), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(G146), .ZN(new_n299));
  OR2_X1    g113(.A1(KEYINPUT68), .A2(G953), .ZN(new_n300));
  INV_X1    g114(.A(G237), .ZN(new_n301));
  NAND2_X1  g115(.A1(KEYINPUT68), .A2(G953), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n300), .A2(G214), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n235), .ZN(new_n304));
  AND2_X1   g118(.A1(KEYINPUT68), .A2(G953), .ZN(new_n305));
  NOR2_X1   g119(.A1(KEYINPUT68), .A2(G953), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n307), .A2(G143), .A3(G214), .A4(new_n301), .ZN(new_n308));
  INV_X1    g122(.A(G131), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n304), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(new_n304), .B2(new_n308), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n296), .B(new_n299), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n304), .A2(new_n308), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(KEYINPUT18), .A3(G131), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n292), .A2(G146), .A3(new_n293), .ZN(new_n315));
  INV_X1    g129(.A(new_n290), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n233), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(KEYINPUT18), .A2(G131), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n304), .A2(new_n308), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n314), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n312), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(G113), .B(G122), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(new_n203), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n299), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT78), .A4(G146), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n297), .A2(new_n298), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n233), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n328), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n311), .A2(KEYINPUT17), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n310), .A2(new_n311), .A3(KEYINPUT17), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n324), .B(new_n321), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n286), .B1(new_n326), .B2(new_n336), .ZN(new_n337));
  XOR2_X1   g151(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n338));
  OAI21_X1  g152(.A(new_n284), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n338), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n324), .B1(new_n312), .B2(new_n321), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT17), .ZN(new_n342));
  AOI211_X1 g156(.A(new_n342), .B(new_n309), .C1(new_n304), .C2(new_n308), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n328), .A2(new_n329), .A3(new_n331), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n311), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n304), .A2(new_n308), .A3(new_n309), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n342), .A3(new_n347), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n318), .A2(new_n320), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n345), .A2(new_n348), .B1(new_n349), .B2(new_n314), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n341), .B1(new_n350), .B2(new_n324), .ZN(new_n351));
  OAI211_X1 g165(.A(KEYINPUT90), .B(new_n340), .C1(new_n351), .C2(new_n286), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT20), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n337), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n339), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n350), .A2(new_n324), .ZN(new_n356));
  INV_X1    g170(.A(new_n336), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n278), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G475), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G952), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(G953), .ZN(new_n362));
  NAND2_X1  g176(.A1(G234), .A2(G237), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XOR2_X1   g178(.A(new_n364), .B(KEYINPUT92), .Z(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT21), .B(G898), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n307), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(G902), .A3(new_n363), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n365), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n193), .A2(KEYINPUT14), .A3(G122), .ZN(new_n371));
  XOR2_X1   g185(.A(G116), .B(G122), .Z(new_n372));
  OAI211_X1 g186(.A(G107), .B(new_n371), .C1(new_n372), .C2(KEYINPUT14), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n235), .A2(G128), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n247), .A2(G143), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G134), .ZN(new_n377));
  INV_X1    g191(.A(G134), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n374), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(G116), .B(G122), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n200), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n373), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT91), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n373), .A2(new_n380), .A3(KEYINPUT91), .A4(new_n382), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n372), .A2(G107), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n382), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT13), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n374), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n375), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n374), .A2(new_n389), .ZN(new_n392));
  OAI21_X1  g206(.A(G134), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n388), .A2(new_n393), .A3(new_n379), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n385), .A2(new_n386), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT9), .B(G234), .ZN(new_n396));
  INV_X1    g210(.A(G217), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n396), .A2(new_n397), .A3(G953), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n385), .A2(new_n386), .A3(new_n394), .A4(new_n398), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n278), .ZN(new_n403));
  INV_X1    g217(.A(G478), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(KEYINPUT15), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n403), .B(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  AND4_X1   g221(.A1(new_n283), .A2(new_n360), .A3(new_n370), .A4(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G221), .B1(new_n396), .B2(G902), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n307), .A2(G227), .ZN(new_n410));
  XOR2_X1   g224(.A(G110), .B(G140), .Z(new_n411));
  XNOR2_X1  g225(.A(new_n410), .B(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT64), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT11), .ZN(new_n415));
  INV_X1    g229(.A(G137), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n414), .A2(new_n415), .A3(new_n416), .A4(G134), .ZN(new_n417));
  OAI22_X1  g231(.A1(new_n378), .A2(G137), .B1(KEYINPUT64), .B2(KEYINPUT11), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n420), .B1(new_n416), .B2(G134), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n419), .A2(new_n309), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT65), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n421), .B1(new_n418), .B2(new_n417), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT65), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n426), .A3(new_n309), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n309), .B1(new_n419), .B2(new_n422), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT67), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT67), .ZN(new_n432));
  AOI211_X1 g246(.A(new_n432), .B(new_n429), .C1(new_n424), .C2(new_n427), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n242), .A2(G128), .B1(new_n234), .B2(new_n236), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n248), .A2(new_n234), .A3(new_n236), .ZN(new_n436));
  OAI21_X1  g250(.A(KEYINPUT10), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT82), .B1(new_n437), .B2(new_n267), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT10), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n439), .B1(new_n245), .B2(new_n249), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT82), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n213), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n242), .A2(KEYINPUT81), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT81), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n234), .A2(new_n445), .A3(KEYINPUT1), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(G128), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n436), .B1(new_n447), .B2(new_n244), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n439), .B1(new_n448), .B2(new_n267), .ZN(new_n449));
  INV_X1    g263(.A(new_n217), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(new_n240), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n223), .A2(KEYINPUT4), .A3(new_n212), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n443), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n413), .B1(new_n434), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT83), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n267), .A2(new_n245), .A3(new_n249), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n448), .B2(new_n267), .ZN(new_n458));
  AND4_X1   g272(.A1(new_n426), .A2(new_n419), .A3(new_n309), .A4(new_n422), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n426), .B1(new_n425), .B2(new_n309), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n430), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n458), .A2(new_n461), .A3(KEYINPUT12), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n432), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n428), .A2(KEYINPUT67), .A3(new_n430), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n464), .A3(new_n458), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT12), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AOI22_X1  g282(.A1(new_n438), .A2(new_n442), .B1(new_n451), .B2(new_n452), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n469), .B(new_n449), .C1(new_n431), .C2(new_n433), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT83), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n471), .A3(new_n413), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n456), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n434), .A2(new_n454), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n413), .B1(new_n474), .B2(new_n470), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AOI211_X1 g290(.A(G469), .B(G902), .C1(new_n473), .C2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n434), .A2(new_n454), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n412), .B1(new_n467), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n474), .A2(new_n470), .A3(new_n413), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(G469), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G469), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(new_n278), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n409), .B1(new_n477), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT84), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n409), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n473), .A2(new_n476), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(new_n482), .A3(new_n278), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n481), .A2(new_n484), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT84), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n408), .A2(new_n488), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n240), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n463), .A2(new_n496), .A3(new_n464), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n378), .A2(G137), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n416), .A2(G134), .ZN(new_n499));
  OAI21_X1  g313(.A(G131), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n245), .A2(new_n249), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n428), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n497), .A2(KEYINPUT30), .A3(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n218), .A2(new_n221), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n461), .A2(new_n496), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n502), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT30), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n497), .A2(new_n502), .A3(new_n504), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(KEYINPUT70), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n307), .A2(G210), .A3(new_n301), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n512), .B(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT26), .B(G101), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n512), .A2(new_n513), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n512), .A2(new_n513), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n519), .A2(new_n516), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n510), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT31), .B1(new_n509), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT71), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT28), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n510), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n504), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n506), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n497), .A2(KEYINPUT28), .A3(new_n502), .A4(new_n504), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n517), .A2(new_n521), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT73), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n510), .A2(new_n523), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n503), .A2(new_n508), .ZN(new_n538));
  XOR2_X1   g352(.A(KEYINPUT72), .B(KEYINPUT31), .Z(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n538), .A2(new_n523), .A3(new_n510), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT71), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT31), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n526), .A2(new_n536), .A3(new_n541), .A4(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(G472), .A2(G902), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT32), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n546), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(new_n548), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n545), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT29), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n553), .B1(new_n532), .B2(new_n535), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT74), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n538), .A2(new_n510), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n555), .B1(new_n556), .B2(new_n533), .ZN(new_n557));
  AOI211_X1 g371(.A(KEYINPUT74), .B(new_n523), .C1(new_n538), .C2(new_n510), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n554), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n497), .A2(new_n502), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n529), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n533), .A2(new_n553), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n528), .A2(new_n561), .A3(new_n562), .A4(new_n531), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT75), .ZN(new_n564));
  AOI21_X1  g378(.A(G902), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n565), .B1(new_n564), .B2(new_n563), .ZN(new_n566));
  OAI21_X1  g380(.A(G472), .B1(new_n559), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n549), .A2(new_n552), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n397), .B1(G234), .B2(new_n278), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT25), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT23), .B1(new_n247), .B2(G119), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT76), .ZN(new_n573));
  INV_X1    g387(.A(G119), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n573), .B1(new_n574), .B2(G128), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n572), .B(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(G110), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(KEYINPUT79), .A3(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(G119), .B(G128), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT24), .B(G110), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n578), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(KEYINPUT79), .B1(new_n576), .B2(new_n577), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n299), .B(new_n317), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n577), .B1(new_n576), .B2(KEYINPUT77), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n585), .B1(KEYINPUT77), .B2(new_n576), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n581), .A2(new_n579), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n344), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n307), .A2(G221), .A3(G234), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT22), .B(G137), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n584), .A2(new_n592), .A3(new_n588), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n571), .B1(new_n596), .B2(G902), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n594), .A2(KEYINPUT25), .A3(new_n278), .A4(new_n595), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n570), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n596), .A2(G902), .A3(new_n569), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n495), .A2(new_n568), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  AND2_X1   g417(.A1(new_n488), .A2(new_n494), .ZN(new_n604));
  INV_X1    g418(.A(G472), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n605), .A2(KEYINPUT93), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n545), .A2(new_n278), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n606), .B1(new_n545), .B2(new_n278), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n604), .A2(new_n601), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(G478), .B1(new_n402), .B2(new_n278), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT94), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n612), .A2(KEYINPUT94), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n402), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n400), .A2(KEYINPUT94), .A3(new_n612), .A4(new_n401), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n404), .A2(G902), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n611), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n355), .B2(new_n359), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n620), .A2(new_n283), .A3(new_n370), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n610), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT95), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT34), .B(G104), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  XNOR2_X1  g439(.A(new_n370), .B(KEYINPUT96), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n283), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n337), .A2(new_n338), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n339), .A2(new_n352), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n359), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n627), .A2(new_n630), .A3(new_n407), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n610), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT97), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT35), .B(G107), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  NOR2_X1   g449(.A1(new_n589), .A2(KEYINPUT98), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT98), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n584), .B2(new_n588), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n593), .A2(KEYINPUT36), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n640), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n642), .B1(new_n636), .B2(new_n638), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n569), .A2(G902), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n599), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n607), .A2(new_n608), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n495), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT37), .B(G110), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT99), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n648), .B(new_n650), .ZN(G12));
  NAND3_X1  g465(.A1(new_n641), .A2(new_n645), .A3(new_n643), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n597), .A2(new_n598), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n652), .B1(new_n653), .B2(new_n570), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n283), .ZN(new_n655));
  XOR2_X1   g469(.A(new_n365), .B(KEYINPUT100), .Z(new_n656));
  OAI21_X1  g470(.A(new_n656), .B1(G900), .B2(new_n369), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n629), .A2(new_n406), .A3(new_n359), .A4(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT101), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n655), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n604), .A2(new_n568), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  XNOR2_X1  g478(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n657), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n604), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n669));
  INV_X1    g483(.A(new_n542), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n561), .A2(new_n510), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n670), .B1(new_n671), .B2(new_n535), .ZN(new_n672));
  OAI21_X1  g486(.A(G472), .B1(new_n672), .B2(G902), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n549), .A2(new_n552), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n360), .A2(new_n407), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n280), .A2(new_n282), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NOR4_X1   g493(.A1(new_n676), .A2(new_n679), .A3(new_n188), .A4(new_n654), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n668), .A2(new_n669), .A3(new_n674), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT104), .B(G143), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G45));
  NAND2_X1  g497(.A1(new_n355), .A2(new_n359), .ZN(new_n684));
  INV_X1    g498(.A(new_n619), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n684), .A2(new_n685), .A3(new_n657), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n655), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n604), .A2(new_n568), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  AOI21_X1  g503(.A(new_n467), .B1(KEYINPUT83), .B2(new_n455), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n475), .B1(new_n690), .B2(new_n472), .ZN(new_n691));
  OAI21_X1  g505(.A(G469), .B1(new_n691), .B2(G902), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n491), .A3(new_n409), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n692), .A2(new_n491), .A3(KEYINPUT105), .A4(new_n409), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n695), .A2(new_n621), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n568), .A3(new_n601), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  AND3_X1   g514(.A1(new_n695), .A2(new_n631), .A3(new_n696), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n568), .A3(new_n601), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G116), .ZN(G18));
  NOR2_X1   g517(.A1(new_n684), .A2(new_n406), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n677), .A2(new_n187), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n693), .A2(new_n646), .A3(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n568), .A2(new_n370), .A3(new_n704), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G119), .ZN(G21));
  AND4_X1   g522(.A1(new_n283), .A2(new_n684), .A3(new_n406), .A4(new_n626), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n695), .A2(new_n696), .A3(new_n709), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n525), .A2(new_n541), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n528), .A2(new_n531), .A3(new_n561), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n535), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n550), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n545), .A2(new_n278), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n714), .B1(new_n715), .B2(G472), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n710), .A2(new_n601), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT106), .B(G122), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G24));
  NAND2_X1  g533(.A1(new_n686), .A2(KEYINPUT107), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n620), .A2(new_n721), .A3(new_n657), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n706), .A2(new_n716), .A3(new_n720), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT108), .B(G125), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G27));
  AND3_X1   g539(.A1(new_n620), .A2(new_n721), .A3(new_n657), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n721), .B1(new_n620), .B2(new_n657), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n280), .A2(new_n187), .A3(new_n282), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n409), .B(new_n728), .C1(new_n477), .C2(new_n485), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n568), .A2(new_n730), .A3(new_n601), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT42), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n280), .A2(new_n187), .A3(new_n282), .ZN(new_n734));
  AOI211_X1 g548(.A(new_n489), .B(new_n734), .C1(new_n491), .C2(new_n492), .ZN(new_n735));
  AND4_X1   g549(.A1(KEYINPUT42), .A2(new_n735), .A3(new_n720), .A4(new_n722), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT31), .ZN(new_n737));
  AOI211_X1 g551(.A(KEYINPUT71), .B(new_n737), .C1(new_n537), .C2(new_n538), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n543), .B1(new_n542), .B2(KEYINPUT31), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n536), .A2(new_n541), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n550), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT110), .B1(new_n742), .B2(KEYINPUT32), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n547), .A2(new_n744), .A3(new_n548), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n545), .A2(new_n747), .A3(new_n551), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n747), .B1(new_n545), .B2(new_n551), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n567), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n736), .B(new_n601), .C1(new_n746), .C2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n733), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n733), .A2(new_n751), .A3(KEYINPUT111), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  AND2_X1   g571(.A1(new_n568), .A2(new_n601), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n660), .A2(new_n729), .A3(new_n661), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G134), .ZN(G36));
  NAND2_X1  g575(.A1(new_n360), .A2(new_n685), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT43), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n763), .A2(new_n609), .A3(new_n646), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n764), .A2(KEYINPUT44), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n734), .B1(new_n764), .B2(KEYINPUT44), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n479), .A2(KEYINPUT45), .A3(new_n480), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT45), .B1(new_n479), .B2(new_n480), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n768), .A2(new_n769), .A3(new_n482), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n770), .A2(new_n483), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n477), .B1(new_n771), .B2(KEYINPUT46), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n772), .A2(KEYINPUT112), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(KEYINPUT46), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(KEYINPUT112), .A3(new_n491), .ZN(new_n775));
  OR3_X1    g589(.A1(new_n771), .A2(KEYINPUT113), .A3(KEYINPUT46), .ZN(new_n776));
  OAI21_X1  g590(.A(KEYINPUT113), .B1(new_n771), .B2(KEYINPUT46), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n773), .A2(new_n775), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n778), .A2(new_n409), .A3(new_n666), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n767), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT114), .B(G137), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G39));
  NAND2_X1  g596(.A1(new_n778), .A2(new_n409), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT47), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n778), .A2(KEYINPUT47), .A3(new_n409), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n568), .A2(new_n601), .A3(new_n686), .A4(new_n734), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT115), .Z(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  NAND4_X1  g605(.A1(new_n679), .A2(new_n601), .A3(new_n409), .A4(new_n187), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n692), .A2(new_n491), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  AOI211_X1 g608(.A(new_n762), .B(new_n792), .C1(KEYINPUT49), .C2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n674), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n795), .B(new_n796), .C1(KEYINPUT49), .C2(new_n794), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n602), .A2(new_n698), .A3(new_n702), .A4(new_n648), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n360), .A2(new_n685), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n800), .A2(new_n704), .A3(new_n627), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n604), .A2(new_n609), .A3(new_n601), .A4(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n707), .A2(new_n802), .A3(new_n717), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n407), .A2(new_n657), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n805), .A2(new_n630), .A3(new_n734), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n604), .A2(new_n568), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n730), .A2(new_n716), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n809), .A2(new_n654), .B1(new_n758), .B2(new_n759), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n804), .A2(new_n754), .A3(new_n755), .A4(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n676), .A2(new_n705), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n493), .A2(new_n646), .A3(new_n657), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n674), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n663), .A2(new_n688), .A3(new_n815), .A4(new_n723), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT52), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n798), .B1(new_n811), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n804), .A2(new_n810), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n816), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n663), .A2(new_n723), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT52), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n824), .A2(new_n752), .A3(KEYINPUT53), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n820), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n818), .A2(new_n819), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n824), .A2(new_n798), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n820), .A2(new_n756), .A3(new_n822), .A4(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n819), .B1(new_n829), .B2(new_n818), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n763), .A2(new_n656), .ZN(new_n832));
  INV_X1    g646(.A(new_n693), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n728), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n654), .A3(new_n716), .ZN(new_n836));
  INV_X1    g650(.A(new_n601), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n834), .A2(new_n837), .A3(new_n365), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n796), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n360), .A2(new_n619), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n836), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n716), .A2(new_n601), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n832), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n833), .A2(new_n188), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT117), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n843), .A2(new_n679), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT50), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n843), .A2(KEYINPUT50), .A3(new_n679), .A4(new_n845), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n841), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n843), .A2(new_n728), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT116), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n794), .A2(new_n409), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT118), .B1(new_n787), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n787), .A2(KEYINPUT118), .A3(new_n854), .ZN(new_n857));
  OAI211_X1 g671(.A(KEYINPUT51), .B(new_n850), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n843), .A2(new_n283), .A3(new_n833), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n838), .A2(new_n796), .A3(new_n620), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n860), .A2(new_n362), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n746), .A2(new_n750), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n837), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n835), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g678(.A(KEYINPUT119), .B(KEYINPUT48), .Z(new_n865));
  AND2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n864), .A2(new_n865), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n859), .B(new_n861), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n787), .A2(new_n854), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n850), .B1(new_n869), .B2(new_n852), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT51), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n831), .A2(new_n858), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(G952), .A2(G953), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n797), .B1(new_n873), .B2(new_n874), .ZN(G75));
  AOI21_X1  g689(.A(new_n278), .B1(new_n818), .B2(new_n826), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT56), .B1(new_n876), .B2(G210), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n232), .A2(new_n259), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT120), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT55), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(new_n257), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n877), .A2(new_n881), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n307), .A2(G952), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(G51));
  AOI21_X1  g699(.A(new_n819), .B1(new_n818), .B2(new_n826), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n827), .A2(new_n886), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n483), .B(KEYINPUT57), .Z(new_n888));
  OAI21_X1  g702(.A(new_n490), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n876), .A2(new_n770), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n884), .B1(new_n889), .B2(new_n890), .ZN(G54));
  INV_X1    g705(.A(new_n884), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n876), .A2(KEYINPUT58), .A3(G475), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n892), .B1(new_n893), .B2(new_n351), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n351), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n893), .A2(KEYINPUT121), .A3(new_n351), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(G60));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n900));
  INV_X1    g714(.A(new_n617), .ZN(new_n901));
  NAND2_X1  g715(.A1(G478), .A2(G902), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT59), .Z(new_n903));
  NOR2_X1   g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n818), .A2(new_n826), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT54), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n818), .A2(new_n826), .A3(new_n819), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n900), .B1(new_n909), .B2(new_n884), .ZN(new_n910));
  OAI211_X1 g724(.A(KEYINPUT122), .B(new_n892), .C1(new_n887), .C2(new_n905), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n901), .B1(new_n831), .B2(new_n903), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(G63));
  XNOR2_X1  g727(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n397), .A2(new_n278), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n906), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n596), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n906), .A2(new_n644), .A3(new_n916), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n892), .A3(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n918), .A2(new_n892), .A3(new_n919), .A4(new_n921), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(G66));
  OAI21_X1  g739(.A(G953), .B1(new_n366), .B2(new_n252), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n804), .B2(new_n368), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n879), .B1(G898), .B2(new_n307), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(G69));
  NAND2_X1  g743(.A1(new_n506), .A2(new_n507), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n503), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n294), .A2(new_n295), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n663), .A2(new_n688), .A3(new_n723), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n681), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n681), .A2(new_n935), .A3(KEYINPUT62), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI22_X1  g754(.A1(new_n787), .A2(new_n789), .B1(new_n767), .B2(new_n779), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n800), .A2(new_n704), .A3(new_n734), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n758), .A2(new_n942), .A3(new_n604), .A4(new_n666), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n940), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n934), .B1(new_n944), .B2(new_n368), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n307), .A2(G900), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n935), .A2(new_n760), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n863), .A2(new_n812), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n947), .B1(new_n949), .B2(new_n779), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n941), .A2(new_n756), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n934), .A2(new_n368), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n946), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n945), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(G227), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n946), .B1(new_n955), .B2(new_n368), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT125), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n954), .B(new_n958), .ZN(G72));
  NAND4_X1  g773(.A1(new_n941), .A2(new_n950), .A3(new_n756), .A4(new_n804), .ZN(new_n960));
  NAND2_X1  g774(.A1(G472), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT63), .Z(new_n962));
  AOI211_X1 g776(.A(new_n523), .B(new_n556), .C1(new_n960), .C2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n829), .A2(new_n818), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n557), .A2(new_n558), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n964), .B(new_n962), .C1(new_n670), .C2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n892), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n940), .A2(new_n941), .A3(new_n804), .A4(new_n943), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n968), .A2(KEYINPUT126), .A3(new_n962), .ZN(new_n969));
  AOI21_X1  g783(.A(KEYINPUT126), .B1(new_n968), .B2(new_n962), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n556), .A2(new_n523), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI211_X1 g786(.A(new_n963), .B(new_n967), .C1(new_n969), .C2(new_n972), .ZN(G57));
endmodule


