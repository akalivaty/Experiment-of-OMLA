

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767;

  XNOR2_X1 U369 ( .A(n572), .B(n548), .ZN(n700) );
  XOR2_X1 U370 ( .A(n529), .B(KEYINPUT16), .Z(n346) );
  XNOR2_X2 U371 ( .A(n449), .B(G469), .ZN(n564) );
  INV_X2 U372 ( .A(G128), .ZN(n442) );
  INV_X1 U373 ( .A(KEYINPUT104), .ZN(n348) );
  AND2_X1 U374 ( .A1(n397), .A2(n396), .ZN(n373) );
  NOR2_X1 U375 ( .A1(n399), .A2(n398), .ZN(n555) );
  AND2_X1 U376 ( .A1(n541), .A2(n542), .ZN(n441) );
  XNOR2_X1 U377 ( .A(n471), .B(KEYINPUT67), .ZN(n438) );
  XNOR2_X1 U378 ( .A(n483), .B(n482), .ZN(n604) );
  XNOR2_X1 U379 ( .A(n648), .B(KEYINPUT62), .ZN(n649) );
  BUF_X1 U380 ( .A(G146), .Z(n445) );
  NAND2_X1 U381 ( .A1(n375), .A2(n374), .ZN(n347) );
  NAND2_X1 U382 ( .A1(n375), .A2(n374), .ZN(n674) );
  XNOR2_X1 U383 ( .A(n348), .B(n569), .ZN(n570) );
  XNOR2_X1 U384 ( .A(n349), .B(KEYINPUT105), .ZN(n766) );
  NAND2_X1 U385 ( .A1(n400), .A2(n573), .ZN(n349) );
  NAND2_X2 U386 ( .A1(n368), .A2(n367), .ZN(n372) );
  AND2_X2 U387 ( .A1(n415), .A2(n618), .ZN(n367) );
  AND2_X1 U388 ( .A1(n388), .A2(n419), .ZN(n418) );
  AND2_X1 U389 ( .A1(n383), .A2(n394), .ZN(n350) );
  XNOR2_X2 U390 ( .A(n488), .B(n487), .ZN(n490) );
  OR2_X1 U391 ( .A1(n708), .A2(n351), .ZN(n417) );
  XNOR2_X2 U392 ( .A(n494), .B(KEYINPUT10), .ZN(n519) );
  NOR2_X2 U393 ( .A1(n628), .A2(n627), .ZN(n361) );
  XNOR2_X2 U394 ( .A(n538), .B(KEYINPUT66), .ZN(n687) );
  XNOR2_X1 U395 ( .A(n532), .B(G478), .ZN(n547) );
  INV_X1 U396 ( .A(KEYINPUT47), .ZN(n403) );
  XOR2_X1 U397 ( .A(KEYINPUT12), .B(KEYINPUT95), .Z(n512) );
  XNOR2_X1 U398 ( .A(KEYINPUT96), .B(KEYINPUT94), .ZN(n511) );
  XNOR2_X1 U399 ( .A(G113), .B(G131), .ZN(n514) );
  NOR2_X1 U400 ( .A1(n370), .A2(n376), .ZN(n369) );
  INV_X1 U401 ( .A(n763), .ZN(n376) );
  NOR2_X1 U402 ( .A1(n397), .A2(n396), .ZN(n370) );
  XNOR2_X1 U403 ( .A(n474), .B(G140), .ZN(n450) );
  XNOR2_X1 U404 ( .A(G131), .B(KEYINPUT4), .ZN(n444) );
  INV_X1 U405 ( .A(G122), .ZN(n489) );
  XNOR2_X1 U406 ( .A(n549), .B(n427), .ZN(n704) );
  INV_X1 U407 ( .A(KEYINPUT108), .ZN(n427) );
  BUF_X1 U408 ( .A(n564), .Z(n539) );
  INV_X1 U409 ( .A(n450), .ZN(n421) );
  INV_X1 U410 ( .A(KEYINPUT33), .ZN(n389) );
  NOR2_X1 U411 ( .A1(n664), .A2(n508), .ZN(n411) );
  INV_X1 U412 ( .A(KEYINPUT19), .ZN(n412) );
  INV_X1 U413 ( .A(n539), .ZN(n439) );
  XNOR2_X1 U414 ( .A(n525), .B(n408), .ZN(n546) );
  XNOR2_X1 U415 ( .A(n524), .B(G475), .ZN(n408) );
  XNOR2_X1 U416 ( .A(n631), .B(n630), .ZN(n632) );
  XOR2_X1 U417 ( .A(KEYINPUT88), .B(n634), .Z(n721) );
  INV_X1 U418 ( .A(KEYINPUT40), .ZN(n557) );
  XNOR2_X1 U419 ( .A(n404), .B(n403), .ZN(n545) );
  XOR2_X1 U420 ( .A(n672), .B(KEYINPUT82), .Z(n567) );
  NAND2_X1 U421 ( .A1(n567), .A2(n355), .ZN(n395) );
  OR2_X1 U422 ( .A1(G237), .A2(G902), .ZN(n443) );
  XNOR2_X1 U423 ( .A(KEYINPUT15), .B(G902), .ZN(n625) );
  XNOR2_X1 U424 ( .A(n519), .B(n450), .ZN(n748) );
  XOR2_X1 U425 ( .A(G119), .B(G110), .Z(n451) );
  XNOR2_X1 U426 ( .A(n431), .B(n430), .ZN(n526) );
  INV_X1 U427 ( .A(KEYINPUT8), .ZN(n430) );
  NOR2_X1 U428 ( .A1(G953), .A2(G237), .ZN(n518) );
  XNOR2_X1 U429 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U430 ( .A(G143), .B(G104), .ZN(n509) );
  XOR2_X1 U431 ( .A(G140), .B(G122), .Z(n510) );
  XNOR2_X1 U432 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n495) );
  XNOR2_X1 U433 ( .A(n391), .B(KEYINPUT17), .ZN(n496) );
  INV_X1 U434 ( .A(KEYINPUT18), .ZN(n391) );
  XNOR2_X1 U435 ( .A(KEYINPUT72), .B(KEYINPUT4), .ZN(n492) );
  INV_X1 U436 ( .A(KEYINPUT101), .ZN(n356) );
  NAND2_X1 U437 ( .A1(G234), .A2(G237), .ZN(n461) );
  XNOR2_X1 U438 ( .A(n458), .B(n457), .ZN(n459) );
  INV_X1 U439 ( .A(G902), .ZN(n481) );
  XNOR2_X1 U440 ( .A(G116), .B(KEYINPUT5), .ZN(n475) );
  NAND2_X1 U441 ( .A1(n350), .A2(KEYINPUT80), .ZN(n374) );
  XOR2_X1 U442 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n528) );
  XNOR2_X1 U443 ( .A(n426), .B(KEYINPUT41), .ZN(n682) );
  NAND2_X1 U444 ( .A1(n704), .A2(n550), .ZN(n426) );
  INV_X1 U445 ( .A(KEYINPUT39), .ZN(n556) );
  BUF_X1 U446 ( .A(n604), .Z(n405) );
  XNOR2_X1 U447 ( .A(n435), .B(n433), .ZN(n728) );
  XNOR2_X1 U448 ( .A(n527), .B(n436), .ZN(n435) );
  XNOR2_X1 U449 ( .A(n434), .B(n530), .ZN(n433) );
  XNOR2_X1 U450 ( .A(n528), .B(KEYINPUT98), .ZN(n436) );
  XNOR2_X1 U451 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U452 ( .A(n422), .B(n421), .ZN(n447) );
  XNOR2_X1 U453 ( .A(n446), .B(G101), .ZN(n422) );
  XNOR2_X1 U454 ( .A(n588), .B(KEYINPUT35), .ZN(n440) );
  NAND2_X1 U455 ( .A1(n418), .A2(n417), .ZN(n587) );
  XNOR2_X1 U456 ( .A(n386), .B(KEYINPUT74), .ZN(n662) );
  INV_X1 U457 ( .A(n546), .ZN(n432) );
  INV_X1 U458 ( .A(KEYINPUT56), .ZN(n359) );
  INV_X1 U459 ( .A(G143), .ZN(n645) );
  OR2_X1 U460 ( .A1(n585), .A2(KEYINPUT34), .ZN(n351) );
  NAND2_X1 U461 ( .A1(n547), .A2(n432), .ZN(n664) );
  INV_X1 U462 ( .A(G137), .ZN(n474) );
  AND2_X1 U463 ( .A1(n439), .A2(n382), .ZN(n352) );
  NAND2_X1 U464 ( .A1(n507), .A2(G214), .ZN(n699) );
  XNOR2_X1 U465 ( .A(n557), .B(KEYINPUT107), .ZN(n353) );
  OR2_X1 U466 ( .A1(KEYINPUT65), .A2(KEYINPUT44), .ZN(n354) );
  XNOR2_X1 U467 ( .A(KEYINPUT48), .B(KEYINPUT81), .ZN(n355) );
  INV_X1 U468 ( .A(KEYINPUT80), .ZN(n396) );
  INV_X1 U469 ( .A(n700), .ZN(n398) );
  NOR2_X1 U470 ( .A1(n574), .A2(n664), .ZN(n377) );
  XNOR2_X1 U471 ( .A(n357), .B(n356), .ZN(n577) );
  NOR2_X1 U472 ( .A1(n687), .A2(n576), .ZN(n357) );
  NOR2_X1 U473 ( .A1(n767), .A2(n765), .ZN(n558) );
  NAND2_X1 U474 ( .A1(n373), .A2(n385), .ZN(n371) );
  XNOR2_X1 U475 ( .A(n595), .B(n594), .ZN(n379) );
  XNOR2_X1 U476 ( .A(n359), .B(n636), .ZN(G51) );
  NAND2_X1 U477 ( .A1(n379), .A2(n597), .ZN(n598) );
  OR2_X1 U478 ( .A1(n687), .A2(n576), .ZN(n360) );
  AND2_X2 U479 ( .A1(n371), .A2(n369), .ZN(n375) );
  OR2_X2 U480 ( .A1(n687), .A2(n539), .ZN(n399) );
  INV_X1 U481 ( .A(n531), .ZN(n434) );
  XNOR2_X1 U482 ( .A(n480), .B(n448), .ZN(n726) );
  XNOR2_X1 U483 ( .A(n480), .B(n479), .ZN(n648) );
  BUF_X1 U484 ( .A(n606), .Z(n362) );
  BUF_X1 U485 ( .A(n675), .Z(n737) );
  NAND2_X1 U486 ( .A1(n759), .A2(G234), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n380), .B(n381), .ZN(n363) );
  XNOR2_X1 U488 ( .A(n380), .B(n381), .ZN(n629) );
  BUF_X1 U489 ( .A(n767), .Z(n364) );
  BUF_X1 U490 ( .A(n732), .Z(n365) );
  XNOR2_X1 U491 ( .A(n377), .B(n353), .ZN(n767) );
  XNOR2_X1 U492 ( .A(n402), .B(n455), .ZN(n732) );
  XNOR2_X1 U493 ( .A(n748), .B(n452), .ZN(n402) );
  BUF_X1 U494 ( .A(G107), .Z(n409) );
  NOR2_X1 U495 ( .A1(n675), .A2(n347), .ZN(n366) );
  NAND2_X1 U496 ( .A1(n562), .A2(n411), .ZN(n569) );
  BUF_X1 U497 ( .A(n361), .Z(n731) );
  BUF_X1 U498 ( .A(n572), .Z(n400) );
  OR2_X2 U499 ( .A1(n675), .A2(n674), .ZN(n624) );
  NAND2_X1 U500 ( .A1(n401), .A2(KEYINPUT44), .ZN(n368) );
  XNOR2_X2 U501 ( .A(n372), .B(n623), .ZN(n675) );
  XNOR2_X2 U502 ( .A(n378), .B(n556), .ZN(n574) );
  NAND2_X1 U503 ( .A1(n555), .A2(n441), .ZN(n378) );
  AND2_X1 U504 ( .A1(n379), .A2(n576), .ZN(n611) );
  XNOR2_X2 U505 ( .A(n490), .B(n346), .ZN(n381) );
  INV_X1 U506 ( .A(n501), .ZN(n380) );
  XNOR2_X1 U507 ( .A(n381), .B(KEYINPUT120), .ZN(n744) );
  NAND2_X1 U508 ( .A1(n382), .A2(n582), .ZN(n584) );
  XNOR2_X1 U509 ( .A(n413), .B(n412), .ZN(n382) );
  NAND2_X1 U510 ( .A1(n383), .A2(n394), .ZN(n385) );
  AND2_X2 U511 ( .A1(n384), .A2(n395), .ZN(n383) );
  NAND2_X1 U512 ( .A1(n568), .A2(n355), .ZN(n384) );
  NOR2_X1 U513 ( .A1(n662), .A2(n534), .ZN(n404) );
  NAND2_X1 U514 ( .A1(n387), .A2(n352), .ZN(n386) );
  INV_X1 U515 ( .A(n486), .ZN(n387) );
  NAND2_X1 U516 ( .A1(n708), .A2(KEYINPUT34), .ZN(n388) );
  XNOR2_X2 U517 ( .A(n390), .B(n389), .ZN(n708) );
  NAND2_X1 U518 ( .A1(n577), .A2(n609), .ZN(n390) );
  NAND2_X1 U519 ( .A1(n393), .A2(n392), .ZN(n394) );
  NOR2_X1 U520 ( .A1(n567), .A2(n355), .ZN(n392) );
  INV_X1 U521 ( .A(n568), .ZN(n393) );
  INV_X1 U522 ( .A(n766), .ZN(n397) );
  INV_X1 U523 ( .A(n399), .ZN(n605) );
  INV_X2 U524 ( .A(G146), .ZN(n437) );
  NAND2_X1 U525 ( .A1(n622), .A2(n414), .ZN(n401) );
  OR2_X2 U526 ( .A1(n764), .A2(n354), .ZN(n590) );
  NAND2_X1 U527 ( .A1(n606), .A2(n593), .ZN(n595) );
  XNOR2_X2 U528 ( .A(n584), .B(n583), .ZN(n606) );
  NAND2_X1 U529 ( .A1(n682), .A2(n551), .ZN(n554) );
  NAND2_X1 U530 ( .A1(n406), .A2(n699), .ZN(n410) );
  INV_X1 U531 ( .A(n604), .ZN(n406) );
  XNOR2_X1 U532 ( .A(n407), .B(n517), .ZN(n523) );
  XNOR2_X1 U533 ( .A(n516), .B(n515), .ZN(n407) );
  XNOR2_X1 U534 ( .A(n410), .B(n540), .ZN(n541) );
  BUF_X2 U535 ( .A(n535), .Z(n599) );
  XNOR2_X1 U536 ( .A(n604), .B(KEYINPUT6), .ZN(n609) );
  NOR2_X2 U537 ( .A1(n572), .A2(n508), .ZN(n413) );
  AND2_X1 U538 ( .A1(n621), .A2(n620), .ZN(n414) );
  NAND2_X1 U539 ( .A1(n416), .A2(n429), .ZN(n415) );
  NAND2_X1 U540 ( .A1(n590), .A2(n589), .ZN(n416) );
  AND2_X1 U541 ( .A1(n420), .A2(n586), .ZN(n419) );
  NAND2_X1 U542 ( .A1(n585), .A2(KEYINPUT34), .ZN(n420) );
  XNOR2_X2 U543 ( .A(n423), .B(G104), .ZN(n487) );
  XNOR2_X2 U544 ( .A(G110), .B(G107), .ZN(n423) );
  XNOR2_X2 U545 ( .A(n425), .B(n424), .ZN(n488) );
  XNOR2_X2 U546 ( .A(G119), .B(KEYINPUT3), .ZN(n424) );
  XNOR2_X2 U547 ( .A(G113), .B(G101), .ZN(n425) );
  NAND2_X2 U548 ( .A1(n647), .A2(n428), .ZN(n601) );
  XNOR2_X1 U549 ( .A(n428), .B(G110), .ZN(G12) );
  NAND2_X1 U550 ( .A1(n611), .A2(n600), .ZN(n428) );
  NAND2_X1 U551 ( .A1(n429), .A2(KEYINPUT65), .ZN(n622) );
  XNOR2_X1 U552 ( .A(n620), .B(KEYINPUT84), .ZN(n429) );
  INV_X4 U553 ( .A(G953), .ZN(n759) );
  INV_X1 U554 ( .A(n547), .ZN(n533) );
  XNOR2_X2 U555 ( .A(n437), .B(G125), .ZN(n494) );
  NAND2_X1 U556 ( .A1(n438), .A2(n609), .ZN(n561) );
  NAND2_X1 U557 ( .A1(n438), .A2(n406), .ZN(n485) );
  NOR2_X1 U558 ( .A1(n486), .A2(n539), .ZN(n551) );
  XNOR2_X2 U559 ( .A(n587), .B(n440), .ZN(n764) );
  AND2_X1 U560 ( .A1(n605), .A2(n441), .ZN(n543) );
  XNOR2_X2 U561 ( .A(n442), .B(G143), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n460), .B(n459), .ZN(n535) );
  INV_X1 U563 ( .A(KEYINPUT11), .ZN(n513) );
  XNOR2_X1 U564 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U565 ( .A(n477), .B(n476), .ZN(n478) );
  INV_X1 U566 ( .A(KEYINPUT25), .ZN(n457) );
  XNOR2_X1 U567 ( .A(n451), .B(KEYINPUT23), .ZN(n452) );
  XNOR2_X1 U568 ( .A(KEYINPUT106), .B(KEYINPUT28), .ZN(n484) );
  XNOR2_X1 U569 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U570 ( .A(n633), .B(n632), .ZN(n635) );
  INV_X1 U571 ( .A(KEYINPUT60), .ZN(n642) );
  XNOR2_X2 U572 ( .A(n498), .B(G134), .ZN(n531) );
  XNOR2_X2 U573 ( .A(n531), .B(n444), .ZN(n749) );
  XNOR2_X2 U574 ( .A(n749), .B(n445), .ZN(n480) );
  NAND2_X1 U575 ( .A1(G227), .A2(n759), .ZN(n446) );
  XNOR2_X1 U576 ( .A(n487), .B(n447), .ZN(n448) );
  NOR2_X1 U577 ( .A1(n726), .A2(G902), .ZN(n449) );
  XOR2_X1 U578 ( .A(G128), .B(KEYINPUT24), .Z(n454) );
  NAND2_X1 U579 ( .A1(G221), .A2(n526), .ZN(n453) );
  XNOR2_X1 U580 ( .A(n454), .B(n453), .ZN(n455) );
  NOR2_X1 U581 ( .A1(n732), .A2(G902), .ZN(n460) );
  NAND2_X1 U582 ( .A1(n625), .A2(G234), .ZN(n456) );
  XNOR2_X1 U583 ( .A(n456), .B(KEYINPUT20), .ZN(n468) );
  NAND2_X1 U584 ( .A1(n468), .A2(G217), .ZN(n458) );
  XNOR2_X1 U585 ( .A(n461), .B(KEYINPUT14), .ZN(n580) );
  INV_X1 U586 ( .A(n580), .ZN(n713) );
  NAND2_X1 U587 ( .A1(n759), .A2(G952), .ZN(n578) );
  NOR2_X1 U588 ( .A1(n713), .A2(n578), .ZN(n466) );
  NAND2_X1 U589 ( .A1(G902), .A2(n580), .ZN(n462) );
  NOR2_X1 U590 ( .A1(G900), .A2(n462), .ZN(n463) );
  NAND2_X1 U591 ( .A1(G953), .A2(n463), .ZN(n464) );
  XOR2_X1 U592 ( .A(KEYINPUT102), .B(n464), .Z(n465) );
  NOR2_X1 U593 ( .A1(n466), .A2(n465), .ZN(n467) );
  XOR2_X1 U594 ( .A(KEYINPUT76), .B(n467), .Z(n542) );
  NAND2_X1 U595 ( .A1(G221), .A2(n468), .ZN(n469) );
  XNOR2_X1 U596 ( .A(KEYINPUT21), .B(n469), .ZN(n683) );
  INV_X1 U597 ( .A(n683), .ZN(n536) );
  AND2_X1 U598 ( .A1(n542), .A2(n536), .ZN(n470) );
  NAND2_X1 U599 ( .A1(n599), .A2(n470), .ZN(n471) );
  XOR2_X1 U600 ( .A(KEYINPUT71), .B(KEYINPUT93), .Z(n473) );
  NAND2_X1 U601 ( .A1(n518), .A2(G210), .ZN(n472) );
  XNOR2_X1 U602 ( .A(n473), .B(n472), .ZN(n477) );
  XNOR2_X1 U603 ( .A(n488), .B(n478), .ZN(n479) );
  NAND2_X1 U604 ( .A1(n648), .A2(n481), .ZN(n483) );
  XOR2_X1 U605 ( .A(G472), .B(KEYINPUT68), .Z(n482) );
  XNOR2_X1 U606 ( .A(n489), .B(G116), .ZN(n529) );
  NAND2_X1 U607 ( .A1(n759), .A2(G224), .ZN(n491) );
  XNOR2_X1 U608 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U609 ( .A(n494), .B(n493), .ZN(n500) );
  XNOR2_X1 U610 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U611 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U612 ( .A(n500), .B(n499), .ZN(n501) );
  NAND2_X1 U613 ( .A1(n629), .A2(n625), .ZN(n506) );
  XNOR2_X1 U614 ( .A(KEYINPUT75), .B(KEYINPUT91), .ZN(n502) );
  XNOR2_X1 U615 ( .A(n502), .B(KEYINPUT92), .ZN(n504) );
  XNOR2_X1 U616 ( .A(KEYINPUT70), .B(n443), .ZN(n507) );
  NAND2_X1 U617 ( .A1(n507), .A2(G210), .ZN(n503) );
  XNOR2_X1 U618 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X2 U619 ( .A(n506), .B(n505), .ZN(n572) );
  INV_X1 U620 ( .A(n699), .ZN(n508) );
  XNOR2_X1 U621 ( .A(n510), .B(n509), .ZN(n517) );
  XNOR2_X1 U622 ( .A(n512), .B(n511), .ZN(n516) );
  NAND2_X1 U623 ( .A1(G214), .A2(n518), .ZN(n521) );
  BUF_X1 U624 ( .A(n519), .Z(n520) );
  XNOR2_X1 U625 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U626 ( .A(n523), .B(n522), .ZN(n638) );
  NOR2_X1 U627 ( .A1(G902), .A2(n638), .ZN(n525) );
  XNOR2_X1 U628 ( .A(KEYINPUT13), .B(KEYINPUT97), .ZN(n524) );
  NAND2_X1 U629 ( .A1(G217), .A2(n526), .ZN(n527) );
  XNOR2_X1 U630 ( .A(n409), .B(n529), .ZN(n530) );
  NOR2_X1 U631 ( .A1(n728), .A2(G902), .ZN(n532) );
  NAND2_X1 U632 ( .A1(n546), .A2(n533), .ZN(n668) );
  NAND2_X1 U633 ( .A1(n668), .A2(n664), .ZN(n703) );
  INV_X1 U634 ( .A(n703), .ZN(n534) );
  INV_X1 U635 ( .A(n535), .ZN(n537) );
  NAND2_X1 U636 ( .A1(n537), .A2(n536), .ZN(n538) );
  INV_X1 U637 ( .A(KEYINPUT30), .ZN(n540) );
  NOR2_X1 U638 ( .A1(n547), .A2(n546), .ZN(n586) );
  NAND2_X1 U639 ( .A1(n543), .A2(n586), .ZN(n544) );
  NOR2_X1 U640 ( .A1(n544), .A2(n400), .ZN(n644) );
  NOR2_X1 U641 ( .A1(n545), .A2(n644), .ZN(n560) );
  NAND2_X1 U642 ( .A1(n547), .A2(n546), .ZN(n702) );
  INV_X1 U643 ( .A(n702), .ZN(n550) );
  XOR2_X1 U644 ( .A(KEYINPUT69), .B(KEYINPUT38), .Z(n548) );
  NAND2_X1 U645 ( .A1(n700), .A2(n699), .ZN(n549) );
  XNOR2_X1 U646 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n552) );
  XNOR2_X1 U647 ( .A(n552), .B(KEYINPUT42), .ZN(n553) );
  XNOR2_X1 U648 ( .A(n554), .B(n553), .ZN(n765) );
  XNOR2_X1 U649 ( .A(n558), .B(KEYINPUT46), .ZN(n559) );
  NAND2_X1 U650 ( .A1(n559), .A2(n560), .ZN(n568) );
  XNOR2_X1 U651 ( .A(n561), .B(KEYINPUT103), .ZN(n562) );
  NOR2_X1 U652 ( .A1(n569), .A2(n400), .ZN(n563) );
  XNOR2_X1 U653 ( .A(n563), .B(KEYINPUT36), .ZN(n566) );
  XNOR2_X2 U654 ( .A(n564), .B(KEYINPUT1), .ZN(n576) );
  INV_X1 U655 ( .A(n576), .ZN(n565) );
  NAND2_X1 U656 ( .A1(n566), .A2(n565), .ZN(n672) );
  NAND2_X1 U657 ( .A1(n570), .A2(n576), .ZN(n571) );
  XNOR2_X1 U658 ( .A(KEYINPUT43), .B(n571), .ZN(n573) );
  NOR2_X1 U659 ( .A1(n668), .A2(n574), .ZN(n575) );
  XNOR2_X1 U660 ( .A(n575), .B(KEYINPUT111), .ZN(n763) );
  NOR2_X1 U661 ( .A1(G898), .A2(n759), .ZN(n743) );
  NAND2_X1 U662 ( .A1(n743), .A2(G902), .ZN(n579) );
  NAND2_X1 U663 ( .A1(n579), .A2(n578), .ZN(n581) );
  AND2_X1 U664 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U665 ( .A(KEYINPUT87), .B(KEYINPUT0), .ZN(n583) );
  INV_X1 U666 ( .A(n606), .ZN(n585) );
  INV_X1 U667 ( .A(KEYINPUT73), .ZN(n588) );
  NAND2_X1 U668 ( .A1(n764), .A2(KEYINPUT65), .ZN(n589) );
  NOR2_X1 U669 ( .A1(n702), .A2(n683), .ZN(n592) );
  INV_X1 U670 ( .A(KEYINPUT99), .ZN(n591) );
  XNOR2_X1 U671 ( .A(n592), .B(n591), .ZN(n593) );
  INV_X1 U672 ( .A(KEYINPUT22), .ZN(n594) );
  XNOR2_X1 U673 ( .A(n599), .B(KEYINPUT100), .ZN(n684) );
  NOR2_X1 U674 ( .A1(n576), .A2(n609), .ZN(n596) );
  AND2_X1 U675 ( .A1(n684), .A2(n596), .ZN(n597) );
  XNOR2_X2 U676 ( .A(n598), .B(KEYINPUT32), .ZN(n647) );
  AND2_X1 U677 ( .A1(n405), .A2(n599), .ZN(n600) );
  XNOR2_X2 U678 ( .A(n601), .B(KEYINPUT85), .ZN(n620) );
  NOR2_X1 U679 ( .A1(n360), .A2(n405), .ZN(n695) );
  NAND2_X1 U680 ( .A1(n695), .A2(n362), .ZN(n603) );
  INV_X1 U681 ( .A(KEYINPUT31), .ZN(n602) );
  XNOR2_X1 U682 ( .A(n603), .B(n602), .ZN(n667) );
  AND2_X1 U683 ( .A1(n605), .A2(n405), .ZN(n607) );
  NAND2_X1 U684 ( .A1(n607), .A2(n362), .ZN(n655) );
  NAND2_X1 U685 ( .A1(n667), .A2(n655), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n608), .A2(n703), .ZN(n612) );
  NOR2_X1 U687 ( .A1(n684), .A2(n609), .ZN(n610) );
  NAND2_X1 U688 ( .A1(n611), .A2(n610), .ZN(n653) );
  AND2_X1 U689 ( .A1(n612), .A2(n653), .ZN(n614) );
  AND2_X1 U690 ( .A1(KEYINPUT44), .A2(n614), .ZN(n613) );
  NAND2_X1 U691 ( .A1(n764), .A2(n613), .ZN(n617) );
  INV_X1 U692 ( .A(n614), .ZN(n615) );
  OR2_X1 U693 ( .A1(n615), .A2(KEYINPUT83), .ZN(n616) );
  NAND2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n618) );
  INV_X1 U695 ( .A(KEYINPUT83), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n764), .A2(n619), .ZN(n621) );
  INV_X1 U697 ( .A(KEYINPUT45), .ZN(n623) );
  XNOR2_X1 U698 ( .A(n366), .B(KEYINPUT2), .ZN(n628) );
  NAND2_X1 U699 ( .A1(n624), .A2(KEYINPUT79), .ZN(n626) );
  XNOR2_X1 U700 ( .A(n626), .B(n625), .ZN(n627) );
  NOR2_X2 U701 ( .A1(n628), .A2(n627), .ZN(n722) );
  NAND2_X1 U702 ( .A1(n722), .A2(G210), .ZN(n633) );
  XNOR2_X1 U703 ( .A(n363), .B(KEYINPUT54), .ZN(n631) );
  XOR2_X1 U704 ( .A(KEYINPUT55), .B(KEYINPUT86), .Z(n630) );
  NOR2_X1 U705 ( .A1(n759), .A2(G952), .ZN(n634) );
  NAND2_X1 U706 ( .A1(n635), .A2(n721), .ZN(n636) );
  NAND2_X1 U707 ( .A1(n361), .A2(G475), .ZN(n640) );
  XNOR2_X1 U708 ( .A(KEYINPUT64), .B(KEYINPUT59), .ZN(n637) );
  XNOR2_X1 U709 ( .A(n640), .B(n639), .ZN(n641) );
  NAND2_X1 U710 ( .A1(n641), .A2(n721), .ZN(n643) );
  XNOR2_X1 U711 ( .A(n643), .B(n642), .ZN(G60) );
  XNOR2_X1 U712 ( .A(n645), .B(n644), .ZN(G45) );
  XOR2_X1 U713 ( .A(G119), .B(KEYINPUT127), .Z(n646) );
  XNOR2_X1 U714 ( .A(n647), .B(n646), .ZN(G21) );
  NAND2_X1 U715 ( .A1(n361), .A2(G472), .ZN(n650) );
  XNOR2_X1 U716 ( .A(n650), .B(n649), .ZN(n651) );
  NAND2_X1 U717 ( .A1(n651), .A2(n721), .ZN(n652) );
  XNOR2_X1 U718 ( .A(n652), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U719 ( .A(G101), .B(n653), .ZN(G3) );
  NOR2_X1 U720 ( .A1(n664), .A2(n655), .ZN(n654) );
  XOR2_X1 U721 ( .A(G104), .B(n654), .Z(G6) );
  NOR2_X1 U722 ( .A1(n668), .A2(n655), .ZN(n657) );
  XNOR2_X1 U723 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n656) );
  XNOR2_X1 U724 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U725 ( .A(n409), .B(n658), .ZN(G9) );
  NOR2_X1 U726 ( .A1(n662), .A2(n668), .ZN(n660) );
  XNOR2_X1 U727 ( .A(KEYINPUT112), .B(KEYINPUT29), .ZN(n659) );
  XNOR2_X1 U728 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U729 ( .A(G128), .B(n661), .ZN(G30) );
  NOR2_X1 U730 ( .A1(n662), .A2(n664), .ZN(n663) );
  XOR2_X1 U731 ( .A(n445), .B(n663), .Z(G48) );
  NOR2_X1 U732 ( .A1(n664), .A2(n667), .ZN(n666) );
  XNOR2_X1 U733 ( .A(G113), .B(KEYINPUT113), .ZN(n665) );
  XNOR2_X1 U734 ( .A(n666), .B(n665), .ZN(G15) );
  NOR2_X1 U735 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U736 ( .A(KEYINPUT114), .B(n669), .Z(n670) );
  XNOR2_X1 U737 ( .A(G116), .B(n670), .ZN(G18) );
  XOR2_X1 U738 ( .A(G125), .B(KEYINPUT37), .Z(n671) );
  XNOR2_X1 U739 ( .A(n672), .B(n671), .ZN(G27) );
  NOR2_X1 U740 ( .A1(n366), .A2(KEYINPUT77), .ZN(n673) );
  XNOR2_X1 U741 ( .A(n673), .B(KEYINPUT2), .ZN(n679) );
  INV_X1 U742 ( .A(n347), .ZN(n676) );
  NAND2_X1 U743 ( .A1(n676), .A2(n737), .ZN(n677) );
  NAND2_X1 U744 ( .A1(n677), .A2(KEYINPUT77), .ZN(n678) );
  NAND2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U746 ( .A(n680), .B(KEYINPUT78), .ZN(n681) );
  NAND2_X1 U747 ( .A1(n681), .A2(n759), .ZN(n719) );
  INV_X1 U748 ( .A(n682), .ZN(n698) );
  OR2_X1 U749 ( .A1(n708), .A2(n698), .ZN(n716) );
  NAND2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U751 ( .A(n685), .B(KEYINPUT49), .ZN(n686) );
  XNOR2_X1 U752 ( .A(KEYINPUT115), .B(n686), .ZN(n692) );
  BUF_X1 U753 ( .A(n687), .Z(n688) );
  NAND2_X1 U754 ( .A1(n576), .A2(n688), .ZN(n689) );
  XNOR2_X1 U755 ( .A(n689), .B(KEYINPUT116), .ZN(n690) );
  XNOR2_X1 U756 ( .A(KEYINPUT50), .B(n690), .ZN(n691) );
  NAND2_X1 U757 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U758 ( .A1(n406), .A2(n693), .ZN(n694) );
  NOR2_X1 U759 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U760 ( .A(KEYINPUT51), .B(n696), .Z(n697) );
  NOR2_X1 U761 ( .A1(n698), .A2(n697), .ZN(n710) );
  NOR2_X1 U762 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U763 ( .A1(n702), .A2(n701), .ZN(n706) );
  AND2_X1 U764 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U765 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U766 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U767 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U768 ( .A(n711), .B(KEYINPUT52), .ZN(n712) );
  NOR2_X1 U769 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U770 ( .A1(n714), .A2(G952), .ZN(n715) );
  NAND2_X1 U771 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U772 ( .A(KEYINPUT117), .B(n717), .Z(n718) );
  NOR2_X1 U773 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U774 ( .A(KEYINPUT53), .B(n720), .ZN(G75) );
  INV_X1 U775 ( .A(n721), .ZN(n735) );
  NAND2_X1 U776 ( .A1(n722), .A2(G469), .ZN(n724) );
  XOR2_X1 U777 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n723) );
  XNOR2_X1 U778 ( .A(n724), .B(n723), .ZN(n725) );
  XNOR2_X1 U779 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U780 ( .A1(n735), .A2(n727), .ZN(G54) );
  NAND2_X1 U781 ( .A1(n731), .A2(G478), .ZN(n729) );
  XNOR2_X1 U782 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X1 U783 ( .A1(n730), .A2(n735), .ZN(G63) );
  NAND2_X1 U784 ( .A1(n731), .A2(G217), .ZN(n734) );
  XNOR2_X1 U785 ( .A(n365), .B(KEYINPUT118), .ZN(n733) );
  XNOR2_X1 U786 ( .A(n734), .B(n733), .ZN(n736) );
  NOR2_X1 U787 ( .A1(n736), .A2(n735), .ZN(G66) );
  INV_X1 U788 ( .A(n737), .ZN(n738) );
  NAND2_X1 U789 ( .A1(n738), .A2(n759), .ZN(n742) );
  NAND2_X1 U790 ( .A1(G953), .A2(G224), .ZN(n739) );
  XNOR2_X1 U791 ( .A(KEYINPUT61), .B(n739), .ZN(n740) );
  NAND2_X1 U792 ( .A1(n740), .A2(G898), .ZN(n741) );
  NAND2_X1 U793 ( .A1(n742), .A2(n741), .ZN(n747) );
  NOR2_X1 U794 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U795 ( .A(KEYINPUT119), .B(n745), .Z(n746) );
  XNOR2_X1 U796 ( .A(n747), .B(n746), .ZN(G69) );
  XNOR2_X1 U797 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n751) );
  XNOR2_X1 U798 ( .A(n748), .B(n749), .ZN(n750) );
  XOR2_X1 U799 ( .A(n751), .B(n750), .Z(n755) );
  XNOR2_X1 U800 ( .A(n347), .B(n755), .ZN(n752) );
  XNOR2_X1 U801 ( .A(KEYINPUT123), .B(n752), .ZN(n753) );
  NOR2_X1 U802 ( .A1(G953), .A2(n753), .ZN(n754) );
  XNOR2_X1 U803 ( .A(n754), .B(KEYINPUT124), .ZN(n761) );
  XNOR2_X1 U804 ( .A(G227), .B(n755), .ZN(n756) );
  NAND2_X1 U805 ( .A1(n756), .A2(G900), .ZN(n757) );
  XNOR2_X1 U806 ( .A(KEYINPUT125), .B(n757), .ZN(n758) );
  NOR2_X1 U807 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U808 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U809 ( .A(KEYINPUT126), .B(n762), .Z(G72) );
  XNOR2_X1 U810 ( .A(G134), .B(n763), .ZN(G36) );
  XOR2_X1 U811 ( .A(n764), .B(G122), .Z(G24) );
  XOR2_X1 U812 ( .A(n765), .B(G137), .Z(G39) );
  XOR2_X1 U813 ( .A(G140), .B(n766), .Z(G42) );
  XOR2_X1 U814 ( .A(n364), .B(G131), .Z(G33) );
endmodule

