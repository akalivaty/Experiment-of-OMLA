

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771;

  XNOR2_X1 U371 ( .A(n408), .B(n750), .ZN(n451) );
  INV_X2 U372 ( .A(G953), .ZN(n452) );
  NOR2_X1 U373 ( .A1(G953), .A2(G237), .ZN(n472) );
  XNOR2_X1 U374 ( .A(n502), .B(n501), .ZN(n521) );
  XNOR2_X2 U375 ( .A(n470), .B(n418), .ZN(n611) );
  NOR2_X2 U376 ( .A1(n759), .A2(n582), .ZN(n625) );
  NOR2_X1 U377 ( .A1(n583), .A2(n539), .ZN(n695) );
  OR2_X2 U378 ( .A1(n550), .A2(n536), .ZN(n538) );
  XNOR2_X2 U379 ( .A(n392), .B(KEYINPUT107), .ZN(n550) );
  NAND2_X2 U380 ( .A1(n415), .A2(n412), .ZN(n554) );
  NOR2_X2 U381 ( .A1(n699), .A2(n607), .ZN(n609) );
  XNOR2_X2 U382 ( .A(KEYINPUT71), .B(G101), .ZN(n443) );
  XNOR2_X2 U383 ( .A(n447), .B(n446), .ZN(n659) );
  XNOR2_X2 U384 ( .A(n593), .B(n390), .ZN(n393) );
  NOR2_X1 U385 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X2 U386 ( .A1(n669), .A2(n590), .ZN(n591) );
  XNOR2_X2 U387 ( .A(G119), .B(G110), .ZN(n512) );
  INV_X1 U388 ( .A(G137), .ZN(n433) );
  AND2_X2 U389 ( .A1(n638), .A2(n639), .ZN(n670) );
  NAND2_X1 U390 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U391 ( .A1(n623), .A2(n624), .ZN(n368) );
  OR2_X1 U392 ( .A1(n769), .A2(KEYINPUT88), .ZN(n355) );
  NAND2_X1 U393 ( .A1(n397), .A2(n394), .ZN(n580) );
  AND2_X1 U394 ( .A1(n399), .A2(n398), .ZN(n397) );
  AND2_X1 U395 ( .A1(n385), .A2(n554), .ZN(n724) );
  AND2_X1 U396 ( .A1(n406), .A2(n405), .ZN(n361) );
  NAND2_X2 U397 ( .A1(n383), .A2(n381), .ZN(n392) );
  AND2_X1 U398 ( .A1(n417), .A2(n416), .ZN(n415) );
  XNOR2_X1 U399 ( .A(n410), .B(G113), .ZN(n450) );
  XNOR2_X1 U400 ( .A(KEYINPUT3), .B(G116), .ZN(n410) );
  INV_X1 U401 ( .A(KEYINPUT81), .ZN(n423) );
  BUF_X1 U402 ( .A(n743), .Z(n349) );
  XNOR2_X1 U403 ( .A(n591), .B(KEYINPUT90), .ZN(n350) );
  INV_X1 U404 ( .A(n607), .ZN(n351) );
  XNOR2_X1 U405 ( .A(n591), .B(KEYINPUT90), .ZN(n620) );
  NAND2_X1 U406 ( .A1(n569), .A2(n724), .ZN(n571) );
  INV_X1 U407 ( .A(KEYINPUT80), .ZN(n390) );
  INV_X1 U408 ( .A(G143), .ZN(n424) );
  XNOR2_X1 U409 ( .A(n407), .B(G104), .ZN(n750) );
  INV_X1 U410 ( .A(G107), .ZN(n407) );
  XNOR2_X1 U411 ( .A(n379), .B(KEYINPUT77), .ZN(n378) );
  NAND2_X1 U412 ( .A1(n572), .A2(n573), .ZN(n379) );
  XOR2_X1 U413 ( .A(G113), .B(G104), .Z(n475) );
  XNOR2_X1 U414 ( .A(G143), .B(G122), .ZN(n474) );
  XOR2_X1 U415 ( .A(G131), .B(G140), .Z(n479) );
  NAND2_X1 U416 ( .A1(n452), .A2(G224), .ZN(n453) );
  INV_X1 U417 ( .A(KEYINPUT64), .ZN(n432) );
  XNOR2_X1 U418 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n456) );
  INV_X1 U419 ( .A(KEYINPUT111), .ZN(n387) );
  XNOR2_X1 U420 ( .A(n482), .B(n481), .ZN(n483) );
  NAND2_X1 U421 ( .A1(n414), .A2(n515), .ZN(n413) );
  OR2_X1 U422 ( .A1(n659), .A2(n382), .ZN(n381) );
  AND2_X1 U423 ( .A1(n380), .A2(n384), .ZN(n383) );
  OR2_X1 U424 ( .A1(n354), .A2(G902), .ZN(n382) );
  XNOR2_X1 U425 ( .A(n409), .B(n450), .ZN(n752) );
  XNOR2_X1 U426 ( .A(KEYINPUT16), .B(G122), .ZN(n449) );
  XOR2_X1 U427 ( .A(KEYINPUT24), .B(G140), .Z(n508) );
  XNOR2_X1 U428 ( .A(G128), .B(G137), .ZN(n507) );
  XOR2_X1 U429 ( .A(KEYINPUT72), .B(KEYINPUT8), .Z(n491) );
  XNOR2_X1 U430 ( .A(KEYINPUT74), .B(KEYINPUT75), .ZN(n437) );
  NAND2_X1 U431 ( .A1(n404), .A2(n403), .ZN(n402) );
  NOR2_X1 U432 ( .A1(n353), .A2(n536), .ZN(n403) );
  XNOR2_X1 U433 ( .A(n519), .B(n518), .ZN(n583) );
  NOR2_X1 U434 ( .A1(n376), .A2(n375), .ZN(n374) );
  INV_X1 U435 ( .A(n740), .ZN(n375) );
  INV_X1 U436 ( .A(G237), .ZN(n459) );
  INV_X1 U437 ( .A(G469), .ZN(n414) );
  NAND2_X1 U438 ( .A1(G902), .A2(G469), .ZN(n416) );
  NAND2_X1 U439 ( .A1(n354), .A2(G902), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n401), .B(n400), .ZN(n628) );
  INV_X1 U441 ( .A(KEYINPUT48), .ZN(n400) );
  NAND2_X1 U442 ( .A1(n377), .A2(n373), .ZN(n401) );
  AND2_X1 U443 ( .A1(n378), .A2(n374), .ZN(n373) );
  XNOR2_X1 U444 ( .A(n554), .B(KEYINPUT1), .ZN(n592) );
  INV_X1 U445 ( .A(n594), .ZN(n389) );
  NAND2_X1 U446 ( .A1(n353), .A2(n536), .ZN(n405) );
  XOR2_X1 U447 ( .A(G131), .B(G119), .Z(n441) );
  XNOR2_X1 U448 ( .A(G107), .B(G116), .ZN(n485) );
  XNOR2_X1 U449 ( .A(n477), .B(n476), .ZN(n480) );
  XNOR2_X1 U450 ( .A(n473), .B(n428), .ZN(n477) );
  XNOR2_X1 U451 ( .A(n421), .B(n419), .ZN(n653) );
  XNOR2_X1 U452 ( .A(n458), .B(n420), .ZN(n419) );
  XNOR2_X1 U453 ( .A(n752), .B(n451), .ZN(n421) );
  NAND2_X1 U454 ( .A1(n396), .A2(n395), .ZN(n394) );
  BUF_X1 U455 ( .A(n592), .Z(n578) );
  XNOR2_X1 U456 ( .A(n553), .B(n386), .ZN(n385) );
  XNOR2_X1 U457 ( .A(n552), .B(n387), .ZN(n386) );
  INV_X1 U458 ( .A(KEYINPUT0), .ZN(n418) );
  XNOR2_X1 U459 ( .A(n365), .B(n510), .ZN(n641) );
  XNOR2_X1 U460 ( .A(n511), .B(n514), .ZN(n365) );
  XNOR2_X1 U461 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U462 ( .A(n447), .B(n439), .ZN(n388) );
  INV_X1 U463 ( .A(n597), .ZN(n363) );
  BUF_X1 U464 ( .A(n732), .Z(n735) );
  NOR2_X1 U465 ( .A1(n548), .A2(n597), .ZN(n545) );
  AND2_X1 U466 ( .A1(n563), .A2(n562), .ZN(n736) );
  NOR2_X1 U467 ( .A1(n422), .A2(n679), .ZN(n717) );
  XNOR2_X1 U468 ( .A(KEYINPUT46), .B(KEYINPUT85), .ZN(n352) );
  XNOR2_X1 U469 ( .A(KEYINPUT70), .B(KEYINPUT19), .ZN(n353) );
  XNOR2_X1 U470 ( .A(n448), .B(G472), .ZN(n354) );
  NAND2_X1 U471 ( .A1(n768), .A2(n352), .ZN(n356) );
  XOR2_X1 U472 ( .A(n549), .B(KEYINPUT39), .Z(n357) );
  XOR2_X1 U473 ( .A(KEYINPUT108), .B(KEYINPUT33), .Z(n358) );
  XNOR2_X1 U474 ( .A(KEYINPUT84), .B(KEYINPUT35), .ZN(n359) );
  XOR2_X1 U475 ( .A(KEYINPUT76), .B(KEYINPUT34), .Z(n360) );
  NAND2_X1 U476 ( .A1(n361), .A2(n402), .ZN(n567) );
  XNOR2_X2 U477 ( .A(n589), .B(n588), .ZN(n669) );
  XNOR2_X2 U478 ( .A(n362), .B(n359), .ZN(n769) );
  NAND2_X1 U479 ( .A1(n364), .A2(n363), .ZN(n362) );
  XNOR2_X1 U480 ( .A(n369), .B(n358), .ZN(n680) );
  NAND2_X1 U481 ( .A1(n393), .A2(n389), .ZN(n369) );
  XNOR2_X1 U482 ( .A(n596), .B(n360), .ZN(n364) );
  NAND2_X1 U483 ( .A1(n586), .A2(n585), .ZN(n589) );
  XNOR2_X1 U484 ( .A(n512), .B(n449), .ZN(n409) );
  NAND2_X1 U485 ( .A1(n567), .A2(n469), .ZN(n470) );
  OR2_X2 U486 ( .A1(n574), .A2(n546), .ZN(n572) );
  XNOR2_X1 U487 ( .A(n443), .B(n437), .ZN(n408) );
  NAND2_X1 U488 ( .A1(n542), .A2(n366), .ZN(n543) );
  AND2_X1 U489 ( .A1(n610), .A2(n541), .ZN(n366) );
  NAND2_X1 U490 ( .A1(n372), .A2(n352), .ZN(n371) );
  XNOR2_X2 U491 ( .A(n367), .B(KEYINPUT40), .ZN(n771) );
  NAND2_X1 U492 ( .A1(n580), .A2(n733), .ZN(n367) );
  XNOR2_X2 U493 ( .A(n368), .B(KEYINPUT45), .ZN(n743) );
  NAND2_X1 U494 ( .A1(n670), .A2(G478), .ZN(n665) );
  NAND2_X1 U495 ( .A1(n371), .A2(n370), .ZN(n377) );
  NAND2_X1 U496 ( .A1(n771), .A2(n356), .ZN(n370) );
  INV_X1 U497 ( .A(n771), .ZN(n372) );
  NOR2_X1 U498 ( .A1(n768), .A2(n352), .ZN(n376) );
  NAND2_X1 U499 ( .A1(n659), .A2(n354), .ZN(n380) );
  NAND2_X1 U500 ( .A1(n388), .A2(G469), .ZN(n417) );
  OR2_X1 U501 ( .A1(n388), .A2(n413), .ZN(n412) );
  XNOR2_X1 U502 ( .A(n388), .B(n672), .ZN(n673) );
  XNOR2_X1 U503 ( .A(n392), .B(KEYINPUT6), .ZN(n594) );
  NAND2_X1 U504 ( .A1(n693), .A2(n391), .ZN(n694) );
  AND2_X1 U505 ( .A1(n610), .A2(n391), .ZN(n612) );
  INV_X1 U506 ( .A(n392), .ZN(n391) );
  NAND2_X1 U507 ( .A1(n393), .A2(n392), .ZN(n699) );
  NOR2_X1 U508 ( .A1(n556), .A2(n357), .ZN(n395) );
  INV_X1 U509 ( .A(n548), .ZN(n396) );
  NAND2_X1 U510 ( .A1(n556), .A2(n357), .ZN(n398) );
  NAND2_X1 U511 ( .A1(n548), .A2(n357), .ZN(n399) );
  NAND2_X1 U512 ( .A1(n628), .A2(n627), .ZN(n759) );
  INV_X1 U513 ( .A(n534), .ZN(n404) );
  NAND2_X1 U514 ( .A1(n534), .A2(n353), .ZN(n406) );
  XNOR2_X2 U515 ( .A(n461), .B(n460), .ZN(n534) );
  XNOR2_X2 U516 ( .A(n411), .B(G134), .ZN(n495) );
  XNOR2_X1 U517 ( .A(n411), .B(n457), .ZN(n420) );
  XNOR2_X2 U518 ( .A(n431), .B(n424), .ZN(n411) );
  INV_X1 U519 ( .A(n578), .ZN(n577) );
  NAND2_X1 U520 ( .A1(n653), .A2(n632), .ZN(n461) );
  XNOR2_X1 U521 ( .A(n586), .B(KEYINPUT87), .ZN(n523) );
  AND2_X2 U522 ( .A1(n521), .A2(n594), .ZN(n586) );
  INV_X1 U523 ( .A(n639), .ZN(n422) );
  XNOR2_X2 U524 ( .A(n626), .B(n423), .ZN(n639) );
  XNOR2_X2 U525 ( .A(n495), .B(n434), .ZN(n758) );
  AND2_X1 U526 ( .A1(n351), .A2(n612), .ZN(n425) );
  XOR2_X1 U527 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n426) );
  AND2_X1 U528 ( .A1(n601), .A2(KEYINPUT88), .ZN(n427) );
  AND2_X1 U529 ( .A1(n472), .A2(G214), .ZN(n428) );
  AND2_X1 U530 ( .A1(n555), .A2(n690), .ZN(n429) );
  AND2_X1 U531 ( .A1(n603), .A2(KEYINPUT44), .ZN(n430) );
  INV_X1 U532 ( .A(KEYINPUT47), .ZN(n570) );
  NOR2_X1 U533 ( .A1(n613), .A2(n686), .ZN(n614) );
  INV_X1 U534 ( .A(KEYINPUT105), .ZN(n617) );
  INV_X1 U535 ( .A(KEYINPUT30), .ZN(n537) );
  XNOR2_X1 U536 ( .A(n455), .B(n433), .ZN(n434) );
  BUF_X1 U537 ( .A(n759), .Z(n760) );
  INV_X1 U538 ( .A(KEYINPUT86), .ZN(n549) );
  XNOR2_X1 U539 ( .A(n484), .B(n483), .ZN(n544) );
  BUF_X1 U540 ( .A(n567), .Z(n728) );
  BUF_X1 U541 ( .A(n534), .Z(n574) );
  XNOR2_X2 U542 ( .A(G128), .B(KEYINPUT65), .ZN(n431) );
  XNOR2_X1 U543 ( .A(n432), .B(KEYINPUT4), .ZN(n455) );
  XNOR2_X2 U544 ( .A(n758), .B(G146), .ZN(n447) );
  XOR2_X1 U545 ( .A(G110), .B(n479), .Z(n436) );
  NAND2_X1 U546 ( .A1(G227), .A2(n452), .ZN(n435) );
  XNOR2_X1 U547 ( .A(n436), .B(n435), .ZN(n438) );
  XNOR2_X1 U548 ( .A(n451), .B(n438), .ZN(n439) );
  NAND2_X1 U549 ( .A1(n472), .A2(G210), .ZN(n440) );
  XNOR2_X1 U550 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U551 ( .A(KEYINPUT5), .B(n442), .ZN(n444) );
  XNOR2_X1 U552 ( .A(n443), .B(n444), .ZN(n445) );
  XNOR2_X1 U553 ( .A(n445), .B(n450), .ZN(n446) );
  INV_X1 U554 ( .A(KEYINPUT95), .ZN(n448) );
  AND2_X1 U555 ( .A1(n550), .A2(n577), .ZN(n503) );
  XNOR2_X1 U556 ( .A(n453), .B(KEYINPUT83), .ZN(n454) );
  XNOR2_X1 U557 ( .A(n455), .B(n454), .ZN(n458) );
  XNOR2_X2 U558 ( .A(G146), .B(G125), .ZN(n478) );
  XNOR2_X1 U559 ( .A(n478), .B(n456), .ZN(n457) );
  XNOR2_X1 U560 ( .A(G902), .B(KEYINPUT15), .ZN(n632) );
  INV_X1 U561 ( .A(G902), .ZN(n515) );
  NAND2_X1 U562 ( .A1(n515), .A2(n459), .ZN(n462) );
  NAND2_X1 U563 ( .A1(n462), .A2(G210), .ZN(n460) );
  NAND2_X1 U564 ( .A1(n462), .A2(G214), .ZN(n681) );
  INV_X1 U565 ( .A(n681), .ZN(n536) );
  NAND2_X1 U566 ( .A1(G237), .A2(G234), .ZN(n463) );
  XNOR2_X1 U567 ( .A(n463), .B(KEYINPUT14), .ZN(n464) );
  XNOR2_X1 U568 ( .A(KEYINPUT78), .B(n464), .ZN(n466) );
  AND2_X1 U569 ( .A1(n466), .A2(G953), .ZN(n465) );
  NAND2_X1 U570 ( .A1(G902), .A2(n465), .ZN(n524) );
  NOR2_X1 U571 ( .A1(n524), .A2(G898), .ZN(n468) );
  NAND2_X1 U572 ( .A1(G952), .A2(n466), .ZN(n709) );
  NOR2_X1 U573 ( .A1(G953), .A2(n709), .ZN(n467) );
  XNOR2_X1 U574 ( .A(n467), .B(KEYINPUT92), .ZN(n527) );
  OR2_X1 U575 ( .A1(n468), .A2(n527), .ZN(n469) );
  XNOR2_X1 U576 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n471) );
  XNOR2_X1 U577 ( .A(n426), .B(n471), .ZN(n473) );
  XNOR2_X1 U578 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U579 ( .A(n478), .B(KEYINPUT10), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n479), .B(n513), .ZN(n757) );
  XNOR2_X1 U581 ( .A(n480), .B(n757), .ZN(n645) );
  NOR2_X1 U582 ( .A1(G902), .A2(n645), .ZN(n484) );
  XNOR2_X1 U583 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n482) );
  INV_X1 U584 ( .A(G475), .ZN(n481) );
  XNOR2_X1 U585 ( .A(n485), .B(KEYINPUT101), .ZN(n489) );
  XOR2_X1 U586 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n487) );
  XNOR2_X1 U587 ( .A(G122), .B(KEYINPUT102), .ZN(n486) );
  XNOR2_X1 U588 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U589 ( .A(n489), .B(n488), .Z(n493) );
  NAND2_X1 U590 ( .A1(G234), .A2(n452), .ZN(n490) );
  XNOR2_X1 U591 ( .A(n491), .B(n490), .ZN(n506) );
  NAND2_X1 U592 ( .A1(G217), .A2(n506), .ZN(n492) );
  XNOR2_X1 U593 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U594 ( .A(n495), .B(n494), .ZN(n664) );
  NAND2_X1 U595 ( .A1(n664), .A2(n515), .ZN(n496) );
  XNOR2_X1 U596 ( .A(n496), .B(G478), .ZN(n562) );
  NOR2_X1 U597 ( .A1(n544), .A2(n562), .ZN(n555) );
  XOR2_X1 U598 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n498) );
  NAND2_X1 U599 ( .A1(G234), .A2(n632), .ZN(n497) );
  XNOR2_X1 U600 ( .A(n498), .B(n497), .ZN(n516) );
  AND2_X1 U601 ( .A1(n516), .A2(G221), .ZN(n500) );
  INV_X1 U602 ( .A(KEYINPUT21), .ZN(n499) );
  XNOR2_X1 U603 ( .A(n500), .B(n499), .ZN(n539) );
  INV_X1 U604 ( .A(n539), .ZN(n690) );
  NAND2_X1 U605 ( .A1(n611), .A2(n429), .ZN(n502) );
  INV_X1 U606 ( .A(KEYINPUT22), .ZN(n501) );
  NAND2_X1 U607 ( .A1(n503), .A2(n521), .ZN(n505) );
  INV_X1 U608 ( .A(KEYINPUT68), .ZN(n504) );
  XNOR2_X1 U609 ( .A(n505), .B(n504), .ZN(n520) );
  AND2_X1 U610 ( .A1(n506), .A2(G221), .ZN(n511) );
  XOR2_X1 U611 ( .A(n509), .B(KEYINPUT23), .Z(n510) );
  XNOR2_X1 U612 ( .A(n513), .B(n512), .ZN(n514) );
  NAND2_X1 U613 ( .A1(n641), .A2(n515), .ZN(n519) );
  NAND2_X1 U614 ( .A1(G217), .A2(n516), .ZN(n517) );
  XNOR2_X1 U615 ( .A(KEYINPUT25), .B(n517), .ZN(n518) );
  NAND2_X1 U616 ( .A1(n520), .A2(n583), .ZN(n590) );
  XNOR2_X1 U617 ( .A(n590), .B(G110), .ZN(G12) );
  INV_X1 U618 ( .A(n583), .ZN(n691) );
  NAND2_X1 U619 ( .A1(n691), .A2(n577), .ZN(n522) );
  NOR2_X1 U620 ( .A1(n523), .A2(n522), .ZN(n615) );
  XOR2_X1 U621 ( .A(G101), .B(n615), .Z(G3) );
  XOR2_X1 U622 ( .A(KEYINPUT100), .B(n544), .Z(n563) );
  NOR2_X2 U623 ( .A1(n563), .A2(n562), .ZN(n733) );
  INV_X1 U624 ( .A(n733), .ZN(n564) );
  NOR2_X1 U625 ( .A1(G900), .A2(n524), .ZN(n525) );
  XOR2_X1 U626 ( .A(KEYINPUT109), .B(n525), .Z(n526) );
  OR2_X1 U627 ( .A1(n527), .A2(n526), .ZN(n541) );
  NAND2_X1 U628 ( .A1(n690), .A2(n541), .ZN(n528) );
  XNOR2_X1 U629 ( .A(KEYINPUT73), .B(n528), .ZN(n529) );
  NAND2_X1 U630 ( .A1(n529), .A2(n583), .ZN(n551) );
  OR2_X1 U631 ( .A1(n564), .A2(n551), .ZN(n530) );
  NOR2_X1 U632 ( .A1(n594), .A2(n530), .ZN(n531) );
  NAND2_X1 U633 ( .A1(n531), .A2(n681), .ZN(n575) );
  XOR2_X1 U634 ( .A(n575), .B(KEYINPUT110), .Z(n532) );
  NAND2_X1 U635 ( .A1(n532), .A2(n577), .ZN(n533) );
  XNOR2_X1 U636 ( .A(n533), .B(KEYINPUT43), .ZN(n535) );
  AND2_X1 U637 ( .A1(n535), .A2(n574), .ZN(n581) );
  XOR2_X1 U638 ( .A(n581), .B(G140), .Z(G42) );
  XNOR2_X1 U639 ( .A(n538), .B(n537), .ZN(n542) );
  NAND2_X1 U640 ( .A1(n695), .A2(n554), .ZN(n540) );
  XOR2_X1 U641 ( .A(n540), .B(KEYINPUT94), .Z(n610) );
  XNOR2_X2 U642 ( .A(n543), .B(KEYINPUT82), .ZN(n548) );
  NAND2_X1 U643 ( .A1(n544), .A2(n562), .ZN(n597) );
  INV_X1 U644 ( .A(n545), .ZN(n546) );
  XNOR2_X1 U645 ( .A(n572), .B(G143), .ZN(G45) );
  XOR2_X1 U646 ( .A(KEYINPUT38), .B(KEYINPUT79), .Z(n547) );
  XOR2_X1 U647 ( .A(n547), .B(n574), .Z(n556) );
  NOR2_X1 U648 ( .A1(n551), .A2(n550), .ZN(n553) );
  XNOR2_X1 U649 ( .A(KEYINPUT28), .B(KEYINPUT112), .ZN(n552) );
  INV_X1 U650 ( .A(n555), .ZN(n684) );
  INV_X1 U651 ( .A(n556), .ZN(n682) );
  NAND2_X1 U652 ( .A1(n682), .A2(n681), .ZN(n685) );
  NOR2_X1 U653 ( .A1(n684), .A2(n685), .ZN(n558) );
  XNOR2_X1 U654 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n557) );
  XNOR2_X1 U655 ( .A(n558), .B(n557), .ZN(n702) );
  NAND2_X1 U656 ( .A1(n724), .A2(n702), .ZN(n561) );
  XOR2_X1 U657 ( .A(KEYINPUT115), .B(KEYINPUT42), .Z(n559) );
  XNOR2_X1 U658 ( .A(KEYINPUT114), .B(n559), .ZN(n560) );
  XNOR2_X1 U659 ( .A(n561), .B(n560), .ZN(n768) );
  INV_X1 U660 ( .A(n736), .ZN(n565) );
  NAND2_X1 U661 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U662 ( .A(n566), .B(KEYINPUT103), .ZN(n686) );
  INV_X1 U663 ( .A(n728), .ZN(n568) );
  NOR2_X1 U664 ( .A1(n686), .A2(n568), .ZN(n569) );
  XNOR2_X1 U665 ( .A(n571), .B(n570), .ZN(n573) );
  NOR2_X1 U666 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U667 ( .A(n576), .B(KEYINPUT36), .ZN(n579) );
  NAND2_X1 U668 ( .A1(n579), .A2(n578), .ZN(n740) );
  AND2_X1 U669 ( .A1(n580), .A2(n736), .ZN(n742) );
  NOR2_X1 U670 ( .A1(n742), .A2(n581), .ZN(n627) );
  INV_X1 U671 ( .A(KEYINPUT2), .ZN(n582) );
  AND2_X1 U672 ( .A1(n583), .A2(n578), .ZN(n584) );
  XNOR2_X1 U673 ( .A(n584), .B(KEYINPUT106), .ZN(n585) );
  INV_X1 U674 ( .A(KEYINPUT67), .ZN(n587) );
  XNOR2_X1 U675 ( .A(n587), .B(KEYINPUT32), .ZN(n588) );
  XNOR2_X1 U676 ( .A(n620), .B(KEYINPUT89), .ZN(n599) );
  NAND2_X1 U677 ( .A1(n592), .A2(n695), .ZN(n593) );
  INV_X1 U678 ( .A(n680), .ZN(n595) );
  NAND2_X1 U679 ( .A1(n595), .A2(n351), .ZN(n596) );
  INV_X1 U680 ( .A(n769), .ZN(n598) );
  NAND2_X1 U681 ( .A1(n599), .A2(n598), .ZN(n602) );
  INV_X1 U682 ( .A(KEYINPUT66), .ZN(n600) );
  NOR2_X1 U683 ( .A1(n600), .A2(KEYINPUT44), .ZN(n601) );
  NAND2_X1 U684 ( .A1(n602), .A2(n427), .ZN(n606) );
  NAND2_X1 U685 ( .A1(n769), .A2(KEYINPUT88), .ZN(n604) );
  NAND2_X1 U686 ( .A1(n350), .A2(KEYINPUT66), .ZN(n603) );
  NAND2_X1 U687 ( .A1(n604), .A2(n430), .ZN(n605) );
  NAND2_X1 U688 ( .A1(n606), .A2(n605), .ZN(n624) );
  INV_X1 U689 ( .A(n611), .ZN(n607) );
  XOR2_X1 U690 ( .A(KEYINPUT31), .B(KEYINPUT96), .Z(n608) );
  XNOR2_X1 U691 ( .A(n609), .B(n608), .ZN(n732) );
  NOR2_X1 U692 ( .A1(n732), .A2(n425), .ZN(n613) );
  XNOR2_X1 U693 ( .A(n614), .B(KEYINPUT104), .ZN(n616) );
  NOR2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n618) );
  XNOR2_X1 U695 ( .A(n618), .B(n617), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n619), .A2(n355), .ZN(n622) );
  NOR2_X1 U697 ( .A1(n350), .A2(KEYINPUT66), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n625), .A2(n743), .ZN(n626) );
  AND2_X1 U699 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U700 ( .A1(n629), .A2(n743), .ZN(n677) );
  INV_X1 U701 ( .A(KEYINPUT69), .ZN(n630) );
  NAND2_X1 U702 ( .A1(n630), .A2(KEYINPUT2), .ZN(n631) );
  NAND2_X1 U703 ( .A1(n677), .A2(n631), .ZN(n633) );
  INV_X1 U704 ( .A(n632), .ZN(n634) );
  NAND2_X1 U705 ( .A1(n633), .A2(n634), .ZN(n637) );
  NAND2_X1 U706 ( .A1(n634), .A2(KEYINPUT2), .ZN(n635) );
  NAND2_X1 U707 ( .A1(n635), .A2(KEYINPUT69), .ZN(n636) );
  NAND2_X1 U708 ( .A1(n670), .A2(G217), .ZN(n640) );
  XOR2_X1 U709 ( .A(n641), .B(n640), .Z(n643) );
  INV_X1 U710 ( .A(G952), .ZN(n642) );
  NAND2_X1 U711 ( .A1(n642), .A2(G953), .ZN(n666) );
  INV_X1 U712 ( .A(n666), .ZN(n675) );
  NOR2_X1 U713 ( .A1(n643), .A2(n675), .ZN(G66) );
  NAND2_X1 U714 ( .A1(n670), .A2(G475), .ZN(n647) );
  XNOR2_X1 U715 ( .A(KEYINPUT124), .B(KEYINPUT59), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U717 ( .A(n647), .B(n646), .ZN(n648) );
  NAND2_X1 U718 ( .A1(n648), .A2(n666), .ZN(n650) );
  INV_X1 U719 ( .A(KEYINPUT60), .ZN(n649) );
  XNOR2_X1 U720 ( .A(n650), .B(n649), .ZN(G60) );
  NAND2_X1 U721 ( .A1(n670), .A2(G210), .ZN(n655) );
  XNOR2_X1 U722 ( .A(KEYINPUT91), .B(KEYINPUT54), .ZN(n651) );
  XNOR2_X1 U723 ( .A(n651), .B(KEYINPUT55), .ZN(n652) );
  XNOR2_X1 U724 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U725 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U726 ( .A1(n656), .A2(n666), .ZN(n658) );
  XOR2_X1 U727 ( .A(KEYINPUT122), .B(KEYINPUT56), .Z(n657) );
  XNOR2_X1 U728 ( .A(n658), .B(n657), .ZN(G51) );
  NAND2_X1 U729 ( .A1(n670), .A2(G472), .ZN(n661) );
  XOR2_X1 U730 ( .A(n659), .B(KEYINPUT62), .Z(n660) );
  XNOR2_X1 U731 ( .A(n661), .B(n660), .ZN(n662) );
  NAND2_X1 U732 ( .A1(n662), .A2(n666), .ZN(n663) );
  XNOR2_X1 U733 ( .A(n663), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U734 ( .A(n665), .B(n664), .ZN(n667) );
  NAND2_X1 U735 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U736 ( .A(n668), .B(KEYINPUT125), .ZN(G63) );
  XNOR2_X1 U737 ( .A(n669), .B(G119), .ZN(G21) );
  NAND2_X1 U738 ( .A1(n670), .A2(G469), .ZN(n674) );
  XNOR2_X1 U739 ( .A(KEYINPUT123), .B(KEYINPUT57), .ZN(n671) );
  XNOR2_X1 U740 ( .A(n671), .B(KEYINPUT58), .ZN(n672) );
  XNOR2_X1 U741 ( .A(n674), .B(n673), .ZN(n676) );
  NOR2_X1 U742 ( .A1(n676), .A2(n675), .ZN(G54) );
  INV_X1 U743 ( .A(n677), .ZN(n678) );
  NOR2_X1 U744 ( .A1(n678), .A2(KEYINPUT2), .ZN(n679) );
  BUF_X1 U745 ( .A(n680), .Z(n711) );
  NOR2_X1 U746 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U747 ( .A1(n684), .A2(n683), .ZN(n688) );
  NOR2_X1 U748 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U749 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U750 ( .A1(n711), .A2(n689), .ZN(n705) );
  NOR2_X1 U751 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U752 ( .A(n692), .B(KEYINPUT49), .ZN(n693) );
  XNOR2_X1 U753 ( .A(n694), .B(KEYINPUT119), .ZN(n698) );
  NOR2_X1 U754 ( .A1(n695), .A2(n578), .ZN(n696) );
  XOR2_X1 U755 ( .A(KEYINPUT50), .B(n696), .Z(n697) );
  NAND2_X1 U756 ( .A1(n698), .A2(n697), .ZN(n700) );
  NAND2_X1 U757 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U758 ( .A(KEYINPUT51), .B(n701), .ZN(n703) );
  INV_X1 U759 ( .A(n702), .ZN(n710) );
  NOR2_X1 U760 ( .A1(n703), .A2(n710), .ZN(n704) );
  NOR2_X1 U761 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U762 ( .A(n706), .B(KEYINPUT120), .ZN(n707) );
  XNOR2_X1 U763 ( .A(KEYINPUT52), .B(n707), .ZN(n708) );
  NOR2_X1 U764 ( .A1(n709), .A2(n708), .ZN(n713) );
  NOR2_X1 U765 ( .A1(n711), .A2(n710), .ZN(n712) );
  OR2_X1 U766 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U767 ( .A(n714), .B(KEYINPUT121), .ZN(n715) );
  NAND2_X1 U768 ( .A1(n715), .A2(n452), .ZN(n716) );
  NOR2_X1 U769 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U770 ( .A(n718), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U771 ( .A1(n425), .A2(n733), .ZN(n719) );
  XNOR2_X1 U772 ( .A(n719), .B(G104), .ZN(G6) );
  XNOR2_X1 U773 ( .A(G107), .B(KEYINPUT27), .ZN(n723) );
  XOR2_X1 U774 ( .A(KEYINPUT116), .B(KEYINPUT26), .Z(n721) );
  NAND2_X1 U775 ( .A1(n425), .A2(n736), .ZN(n720) );
  XNOR2_X1 U776 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U777 ( .A(n723), .B(n722), .ZN(G9) );
  INV_X1 U778 ( .A(n724), .ZN(n730) );
  NAND2_X1 U779 ( .A1(n736), .A2(n728), .ZN(n725) );
  NOR2_X1 U780 ( .A1(n730), .A2(n725), .ZN(n727) );
  XNOR2_X1 U781 ( .A(G128), .B(KEYINPUT29), .ZN(n726) );
  XNOR2_X1 U782 ( .A(n727), .B(n726), .ZN(G30) );
  NAND2_X1 U783 ( .A1(n733), .A2(n728), .ZN(n729) );
  NOR2_X1 U784 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U785 ( .A(G146), .B(n731), .Z(G48) );
  NAND2_X1 U786 ( .A1(n735), .A2(n733), .ZN(n734) );
  XNOR2_X1 U787 ( .A(n734), .B(G113), .ZN(G15) );
  XOR2_X1 U788 ( .A(G116), .B(KEYINPUT117), .Z(n738) );
  NAND2_X1 U789 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U790 ( .A(n738), .B(n737), .ZN(G18) );
  XOR2_X1 U791 ( .A(KEYINPUT118), .B(KEYINPUT37), .Z(n739) );
  XNOR2_X1 U792 ( .A(n740), .B(n739), .ZN(n741) );
  XNOR2_X1 U793 ( .A(G125), .B(n741), .ZN(G27) );
  XOR2_X1 U794 ( .A(G134), .B(n742), .Z(G36) );
  INV_X1 U795 ( .A(n349), .ZN(n744) );
  NOR2_X1 U796 ( .A1(n744), .A2(G953), .ZN(n749) );
  INV_X1 U797 ( .A(G898), .ZN(n747) );
  NAND2_X1 U798 ( .A1(G953), .A2(G224), .ZN(n745) );
  XOR2_X1 U799 ( .A(KEYINPUT61), .B(n745), .Z(n746) );
  NOR2_X1 U800 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U801 ( .A1(n749), .A2(n748), .ZN(n756) );
  XOR2_X1 U802 ( .A(n750), .B(G101), .Z(n751) );
  XNOR2_X1 U803 ( .A(n752), .B(n751), .ZN(n754) );
  NOR2_X1 U804 ( .A1(G898), .A2(n452), .ZN(n753) );
  NOR2_X1 U805 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U806 ( .A(n756), .B(n755), .Z(G69) );
  XNOR2_X1 U807 ( .A(n758), .B(n757), .ZN(n763) );
  XNOR2_X1 U808 ( .A(n763), .B(n760), .ZN(n761) );
  NAND2_X1 U809 ( .A1(n761), .A2(n452), .ZN(n762) );
  XNOR2_X1 U810 ( .A(n762), .B(KEYINPUT126), .ZN(n767) );
  XNOR2_X1 U811 ( .A(G227), .B(n763), .ZN(n764) );
  NAND2_X1 U812 ( .A1(n764), .A2(G900), .ZN(n765) );
  NAND2_X1 U813 ( .A1(G953), .A2(n765), .ZN(n766) );
  NAND2_X1 U814 ( .A1(n767), .A2(n766), .ZN(G72) );
  XNOR2_X1 U815 ( .A(G137), .B(n768), .ZN(G39) );
  XNOR2_X1 U816 ( .A(G122), .B(KEYINPUT127), .ZN(n770) );
  XNOR2_X1 U817 ( .A(n770), .B(n769), .ZN(G24) );
  XNOR2_X1 U818 ( .A(n771), .B(G131), .ZN(G33) );
endmodule

