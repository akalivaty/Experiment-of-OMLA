//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n201), .A2(G77), .A3(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  INV_X1    g0010(.A(G77), .ZN(new_n211));
  INV_X1    g0011(.A(G244), .ZN(new_n212));
  INV_X1    g0012(.A(G107), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n211), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT65), .Z(new_n217));
  AOI211_X1 g0017(.A(new_n215), .B(new_n217), .C1(G50), .C2(G226), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G116), .A2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n218), .B(new_n219), .C1(new_n202), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n203), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n207), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n204), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n210), .B(new_n225), .C1(new_n228), .C2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G1), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT66), .B(G45), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  OAI211_X1 g0049(.A(new_n247), .B(G274), .C1(new_n249), .C2(G41), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  OAI21_X1  g0052(.A(KEYINPUT67), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n226), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT67), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G33), .A3(G41), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n253), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n247), .B1(G41), .B2(G45), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G226), .A2(G1698), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n264), .B1(new_n220), .B2(G1698), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n263), .A2(new_n265), .B1(G33), .B2(G97), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  OAI221_X1 g0068(.A(new_n250), .B1(new_n259), .B2(new_n222), .C1(new_n266), .C2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT13), .ZN(new_n270));
  OR2_X1    g0070(.A1(new_n266), .A2(new_n268), .ZN(new_n271));
  INV_X1    g0071(.A(new_n259), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G238), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT13), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n271), .A2(new_n273), .A3(new_n274), .A4(new_n250), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n270), .A2(KEYINPUT69), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT69), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n269), .A2(new_n277), .A3(KEYINPUT13), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(G169), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT74), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n279), .B1(new_n280), .B2(KEYINPUT14), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT70), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n270), .A2(new_n282), .A3(new_n275), .ZN(new_n283));
  OR3_X1    g0083(.A1(new_n269), .A2(new_n282), .A3(KEYINPUT13), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G179), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n280), .A2(KEYINPUT14), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n280), .A2(KEYINPUT14), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n276), .A2(G169), .A3(new_n288), .A4(new_n278), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n281), .A2(new_n286), .A3(new_n287), .A4(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(KEYINPUT73), .A2(KEYINPUT12), .ZN(new_n291));
  OR2_X1    g0091(.A1(KEYINPUT73), .A2(KEYINPUT12), .ZN(new_n292));
  INV_X1    g0092(.A(G13), .ZN(new_n293));
  NOR3_X1   g0093(.A1(new_n293), .A2(new_n227), .A3(G1), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n291), .B(new_n292), .C1(new_n295), .C2(G68), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n203), .ZN(new_n297));
  NAND3_X1  g0097(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n226), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(new_n247), .B2(G20), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OAI221_X1 g0101(.A(new_n296), .B1(new_n297), .B2(new_n291), .C1(new_n301), .C2(new_n203), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n227), .A2(G33), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n303), .A2(new_n211), .B1(new_n227), .B2(G68), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n227), .A2(new_n251), .ZN(new_n305));
  INV_X1    g0105(.A(G50), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n299), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT72), .B(KEYINPUT11), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n308), .B(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n302), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n290), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G190), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n283), .B2(new_n284), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n315), .A2(KEYINPUT71), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n276), .A2(G200), .A3(new_n278), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n317), .A2(new_n311), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(KEYINPUT71), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(G20), .B1(new_n201), .B2(new_n204), .ZN(new_n322));
  INV_X1    g0122(.A(G150), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT8), .B(G58), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n322), .B1(new_n323), .B2(new_n305), .C1(new_n303), .C2(new_n324), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n325), .A2(new_n299), .B1(new_n306), .B2(new_n294), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n306), .B2(new_n301), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT9), .ZN(new_n328));
  NOR2_X1   g0128(.A1(G222), .A2(G1698), .ZN(new_n329));
  INV_X1    g0129(.A(G1698), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(G223), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n263), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n332), .B(new_n267), .C1(G77), .C2(new_n263), .ZN(new_n333));
  INV_X1    g0133(.A(G226), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n333), .B(new_n250), .C1(new_n334), .C2(new_n259), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G200), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n328), .B(new_n336), .C1(new_n314), .C2(new_n335), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT10), .ZN(new_n338));
  INV_X1    g0138(.A(G169), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n327), .B(new_n340), .C1(G179), .C2(new_n335), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n295), .A2(G77), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G20), .A2(G77), .ZN(new_n343));
  XNOR2_X1  g0143(.A(KEYINPUT15), .B(G87), .ZN(new_n344));
  OAI221_X1 g0144(.A(new_n343), .B1(new_n324), .B2(new_n305), .C1(new_n303), .C2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n342), .B1(new_n345), .B2(new_n299), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n300), .A2(G77), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G274), .ZN(new_n349));
  AOI211_X1 g0149(.A(G1), .B(new_n349), .C1(new_n248), .C2(new_n252), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n261), .A2(G33), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n351), .A2(new_n352), .A3(G232), .A4(new_n330), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n351), .A2(new_n352), .A3(G238), .A4(G1698), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n353), .B(new_n354), .C1(new_n263), .C2(new_n213), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n350), .B1(new_n267), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n272), .A2(G244), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n348), .B(KEYINPUT68), .C1(new_n358), .C2(G169), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT68), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n346), .A2(new_n347), .ZN(new_n361));
  AOI21_X1  g0161(.A(G169), .B1(new_n356), .B2(new_n357), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G179), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n358), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n359), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n321), .A2(new_n338), .A3(new_n341), .A4(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G159), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n305), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G58), .A2(G68), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n370), .B(KEYINPUT76), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n204), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n369), .B1(new_n372), .B2(G20), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT75), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n251), .ZN(new_n375));
  NAND2_X1  g0175(.A1(KEYINPUT75), .A2(G33), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(KEYINPUT3), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(G20), .B1(new_n377), .B2(new_n351), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT7), .ZN(new_n379));
  OAI21_X1  g0179(.A(G68), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI211_X1 g0180(.A(KEYINPUT7), .B(G20), .C1(new_n377), .C2(new_n351), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n373), .B(KEYINPUT16), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT77), .ZN(new_n383));
  AND2_X1   g0183(.A1(KEYINPUT75), .A2(G33), .ZN(new_n384));
  NOR2_X1   g0184(.A1(KEYINPUT75), .A2(G33), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n260), .B1(new_n386), .B2(KEYINPUT3), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT7), .B1(new_n387), .B2(G20), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n378), .A2(new_n379), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(G68), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT77), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT16), .A4(new_n373), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT16), .ZN(new_n393));
  INV_X1    g0193(.A(new_n373), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n351), .A2(new_n352), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT7), .B1(new_n395), .B2(new_n227), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT3), .B1(new_n375), .B2(new_n376), .ZN(new_n398));
  OAI211_X1 g0198(.A(KEYINPUT7), .B(new_n227), .C1(new_n398), .C2(new_n262), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n203), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n393), .B1(new_n394), .B2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n383), .A2(new_n392), .A3(new_n299), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n295), .A2(new_n324), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n300), .B2(new_n324), .ZN(new_n404));
  OR2_X1    g0204(.A1(G223), .A2(G1698), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n334), .A2(G1698), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n377), .A2(new_n351), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G33), .A2(G87), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n268), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n257), .A2(G232), .A3(new_n258), .ZN(new_n410));
  NOR3_X1   g0210(.A1(new_n409), .A2(new_n350), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n314), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n411), .B2(G200), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n402), .A2(new_n404), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT17), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n402), .A2(new_n413), .A3(KEYINPUT17), .A4(new_n404), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT78), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n416), .A2(KEYINPUT78), .A3(new_n417), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR4_X1   g0222(.A1(new_n409), .A2(new_n410), .A3(new_n350), .A4(new_n364), .ZN(new_n423));
  INV_X1    g0223(.A(new_n411), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n423), .B1(new_n424), .B2(G169), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n402), .B2(new_n404), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT18), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n358), .A2(G190), .ZN(new_n428));
  INV_X1    g0228(.A(G200), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n428), .B(new_n361), .C1(new_n429), .C2(new_n358), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n422), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n367), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  AOI211_X1 g0233(.A(new_n299), .B(new_n294), .C1(new_n247), .C2(G33), .ZN(new_n434));
  INV_X1    g0234(.A(new_n344), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT82), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n377), .A2(new_n227), .A3(G68), .A4(new_n351), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT19), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n439), .A2(KEYINPUT81), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(KEYINPUT81), .ZN(new_n441));
  INV_X1    g0241(.A(G97), .ZN(new_n442));
  OAI22_X1  g0242(.A1(new_n440), .A2(new_n441), .B1(new_n303), .B2(new_n442), .ZN(new_n443));
  XNOR2_X1  g0243(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n227), .B1(new_n251), .B2(new_n442), .ZN(new_n445));
  NOR2_X1   g0245(.A1(G97), .A2(G107), .ZN(new_n446));
  INV_X1    g0246(.A(G87), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n444), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n438), .A2(new_n443), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n299), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n435), .A2(new_n295), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n437), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  AOI211_X1 g0254(.A(KEYINPUT82), .B(new_n452), .C1(new_n450), .C2(new_n299), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n436), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G45), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n257), .B(G250), .C1(G1), .C2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n247), .A2(G45), .A3(G274), .ZN(new_n459));
  INV_X1    g0259(.A(G116), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n386), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(G238), .A2(G1698), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n462), .B1(new_n212), .B2(G1698), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n461), .B1(new_n387), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n458), .B(new_n459), .C1(new_n464), .C2(new_n268), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n364), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n339), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n456), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n305), .A2(new_n211), .ZN(new_n470));
  XOR2_X1   g0270(.A(new_n470), .B(KEYINPUT79), .Z(new_n471));
  NAND3_X1  g0271(.A1(new_n213), .A2(KEYINPUT6), .A3(G97), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n442), .A2(new_n213), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(new_n446), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n472), .B1(new_n474), .B2(KEYINPUT6), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G20), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n261), .B1(new_n384), .B2(new_n385), .ZN(new_n477));
  AOI21_X1  g0277(.A(G20), .B1(new_n477), .B2(new_n352), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n396), .B1(new_n478), .B2(KEYINPUT7), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n471), .B(new_n476), .C1(new_n479), .C2(new_n213), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n480), .A2(new_n299), .B1(new_n442), .B2(new_n294), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n434), .A2(G97), .ZN(new_n482));
  OR2_X1    g0282(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n483), .A2(new_n484), .A3(new_n247), .A4(G45), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(new_n349), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n257), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n486), .B1(new_n488), .B2(G257), .ZN(new_n489));
  INV_X1    g0289(.A(G250), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n395), .A2(new_n490), .A3(new_n330), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n377), .A2(G244), .A3(new_n330), .A4(new_n351), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G283), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT80), .ZN(new_n496));
  XNOR2_X1  g0296(.A(new_n495), .B(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n492), .A2(new_n212), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n498), .A2(new_n330), .A3(new_n351), .A4(new_n352), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n489), .B1(new_n501), .B2(new_n268), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n481), .A2(new_n482), .B1(new_n502), .B2(new_n339), .ZN(new_n503));
  INV_X1    g0303(.A(new_n486), .ZN(new_n504));
  INV_X1    g0304(.A(G257), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n504), .B1(new_n505), .B2(new_n487), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n494), .A2(new_n497), .A3(new_n499), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n507), .B2(new_n267), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n364), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n502), .A2(G200), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n508), .A2(G190), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n511), .A2(new_n512), .A3(new_n481), .A4(new_n482), .ZN(new_n513));
  INV_X1    g0313(.A(new_n299), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n449), .A2(new_n443), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n514), .B1(new_n515), .B2(new_n438), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT82), .B1(new_n516), .B2(new_n452), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n451), .A2(new_n437), .A3(new_n453), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n466), .A2(G190), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n465), .A2(G200), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n434), .A2(G87), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n519), .A2(new_n520), .A3(new_n521), .A4(new_n523), .ZN(new_n524));
  AND4_X1   g0324(.A1(new_n469), .A2(new_n510), .A3(new_n513), .A4(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n447), .A2(G20), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n377), .A2(new_n351), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT83), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT83), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n377), .A2(new_n529), .A3(new_n351), .A4(new_n526), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(KEYINPUT22), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT22), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n263), .A2(new_n532), .A3(new_n526), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n461), .A2(new_n227), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT84), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT84), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n461), .A2(new_n537), .A3(new_n227), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n227), .A2(G107), .ZN(new_n540));
  XNOR2_X1  g0340(.A(new_n540), .B(KEYINPUT23), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n534), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT85), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT85), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n534), .A2(new_n544), .A3(new_n539), .A4(new_n541), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(KEYINPUT24), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT24), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n542), .A2(KEYINPUT85), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n299), .A3(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n487), .A2(new_n214), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n490), .A2(new_n330), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n505), .A2(G1698), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n377), .A2(new_n351), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(G294), .B1(new_n384), .B2(new_n385), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n268), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n550), .A2(new_n555), .A3(new_n486), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G190), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT25), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n295), .B2(G107), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n294), .A2(KEYINPUT25), .A3(new_n213), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n434), .A2(G107), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n550), .A2(new_n555), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n504), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G200), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n549), .A2(new_n557), .A3(new_n561), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n525), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(KEYINPUT86), .A3(G169), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT86), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n556), .B2(new_n339), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n556), .A2(G179), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n567), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n549), .B2(new_n561), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n505), .A2(new_n330), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n214), .A2(G1698), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n387), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n395), .A2(G303), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n578), .A2(new_n267), .B1(G270), .B2(new_n488), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n504), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n514), .B1(G20), .B2(new_n460), .ZN(new_n581));
  AOI21_X1  g0381(.A(G20), .B1(new_n251), .B2(G97), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n497), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT20), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n581), .A2(new_n583), .A3(KEYINPUT20), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n295), .A2(G116), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n434), .A2(G116), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n580), .A2(new_n592), .A3(G169), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n579), .A2(G190), .A3(new_n504), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n578), .A2(new_n267), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n488), .A2(G270), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n598), .A2(new_n504), .A3(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n596), .B(new_n597), .C1(new_n600), .C2(new_n429), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n580), .A2(new_n592), .A3(KEYINPUT21), .A4(G169), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n600), .A2(G179), .A3(new_n592), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n595), .A2(new_n601), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  NOR4_X1   g0404(.A1(new_n433), .A2(new_n566), .A3(new_n573), .A4(new_n604), .ZN(G372));
  INV_X1    g0405(.A(new_n320), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n313), .B1(new_n606), .B2(new_n366), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n607), .A2(new_n422), .ZN(new_n608));
  INV_X1    g0408(.A(new_n427), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n338), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n341), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT87), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n549), .A2(new_n561), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n614), .B2(new_n571), .ZN(new_n615));
  AOI211_X1 g0415(.A(KEYINPUT87), .B(new_n572), .C1(new_n549), .C2(new_n561), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n595), .A2(new_n603), .A3(new_n602), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n566), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n469), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n503), .A2(new_n469), .A3(new_n524), .A4(new_n509), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n621), .B1(new_n622), .B2(KEYINPUT26), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT89), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n481), .A2(new_n482), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n502), .A2(new_n339), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n625), .A2(new_n626), .A3(new_n509), .ZN(new_n627));
  XOR2_X1   g0427(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n628));
  NAND4_X1  g0428(.A1(new_n627), .A2(new_n469), .A3(new_n524), .A4(new_n628), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n623), .A2(new_n624), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n624), .B1(new_n623), .B2(new_n629), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n432), .B1(new_n620), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n612), .A2(new_n633), .ZN(G369));
  NOR2_X1   g0434(.A1(new_n293), .A2(G20), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n247), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(G213), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n639), .B(KEYINPUT90), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(G343), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n592), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n643), .B(KEYINPUT91), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n618), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n604), .B2(new_n644), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G330), .ZN(new_n647));
  XOR2_X1   g0447(.A(new_n647), .B(KEYINPUT92), .Z(new_n648));
  INV_X1    g0448(.A(new_n573), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n649), .A2(new_n565), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n614), .A2(new_n642), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n649), .B2(new_n641), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n641), .B1(new_n615), .B2(new_n616), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n619), .A2(new_n642), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n654), .A2(new_n655), .A3(new_n657), .ZN(G399));
  INV_X1    g0458(.A(new_n208), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(G41), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G1), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n446), .A2(new_n447), .A3(new_n460), .ZN(new_n663));
  OAI22_X1  g0463(.A1(new_n662), .A2(new_n663), .B1(new_n229), .B2(new_n661), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n664), .B(KEYINPUT28), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n641), .B1(new_n620), .B2(new_n632), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(KEYINPUT29), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT29), .ZN(new_n668));
  INV_X1    g0468(.A(new_n622), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(new_n628), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT26), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n621), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n524), .B1(new_n573), .B2(new_n618), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n510), .A2(new_n513), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n565), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n670), .B(new_n672), .C1(new_n673), .C2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n668), .B1(new_n676), .B2(new_n641), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n667), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G330), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT30), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n600), .A2(new_n466), .A3(G179), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n508), .A2(new_n562), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AND4_X1   g0483(.A1(G179), .A2(new_n466), .A3(new_n579), .A4(new_n504), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n684), .A2(KEYINPUT30), .A3(new_n508), .A4(new_n562), .ZN(new_n685));
  AOI21_X1  g0485(.A(G179), .B1(new_n579), .B2(new_n504), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n686), .A2(new_n465), .A3(new_n502), .A4(new_n563), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n683), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n688), .A2(KEYINPUT31), .A3(new_n642), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT31), .B1(new_n688), .B2(new_n642), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n604), .B1(new_n614), .B2(new_n571), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n692), .A2(new_n525), .A3(new_n565), .A4(new_n641), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n679), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n678), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n665), .B1(new_n697), .B2(G1), .ZN(G364));
  INV_X1    g0498(.A(new_n648), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n662), .B1(G45), .B2(new_n635), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n699), .B(new_n701), .C1(G330), .C2(new_n646), .ZN(new_n702));
  INV_X1    g0502(.A(new_n646), .ZN(new_n703));
  NOR2_X1   g0503(.A1(G13), .A2(G33), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G20), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n263), .A2(G355), .A3(new_n208), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n245), .A2(new_n457), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n387), .A2(new_n659), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n229), .B2(new_n249), .ZN(new_n711));
  OAI221_X1 g0511(.A(new_n708), .B1(G116), .B2(new_n208), .C1(new_n709), .C2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n226), .B1(G20), .B2(new_n339), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n706), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n429), .A2(G179), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(G20), .A3(G190), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n447), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n227), .A2(new_n364), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(G190), .A3(G200), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n718), .B1(G50), .B2(new_n721), .ZN(new_n722));
  XOR2_X1   g0522(.A(new_n719), .B(KEYINPUT93), .Z(new_n723));
  NOR2_X1   g0523(.A1(new_n314), .A2(G200), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n723), .A2(new_n314), .A3(new_n429), .ZN(new_n726));
  OAI221_X1 g0526(.A(new_n722), .B1(new_n725), .B2(new_n202), .C1(new_n211), .C2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(G179), .A2(G200), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(G20), .A3(new_n314), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n368), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT32), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n719), .A2(new_n314), .A3(G200), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n227), .B1(new_n728), .B2(G190), .ZN(new_n733));
  OAI221_X1 g0533(.A(new_n731), .B1(new_n203), .B2(new_n732), .C1(new_n442), .C2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n716), .A2(G20), .A3(new_n314), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n213), .ZN(new_n736));
  NOR4_X1   g0536(.A1(new_n727), .A2(new_n734), .A3(new_n395), .A4(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G311), .ZN(new_n738));
  INV_X1    g0538(.A(G322), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n726), .A2(new_n738), .B1(new_n725), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G283), .ZN(new_n741));
  INV_X1    g0541(.A(G329), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n735), .A2(new_n741), .B1(new_n742), .B2(new_n729), .ZN(new_n743));
  XOR2_X1   g0543(.A(new_n743), .B(KEYINPUT94), .Z(new_n744));
  INV_X1    g0544(.A(new_n732), .ZN(new_n745));
  INV_X1    g0545(.A(G317), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(KEYINPUT33), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n746), .A2(KEYINPUT33), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n721), .A2(G326), .ZN(new_n750));
  INV_X1    g0550(.A(G294), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n749), .B(new_n750), .C1(new_n751), .C2(new_n733), .ZN(new_n752));
  INV_X1    g0552(.A(G303), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n395), .B1(new_n717), .B2(new_n753), .ZN(new_n754));
  NOR4_X1   g0554(.A1(new_n740), .A2(new_n744), .A3(new_n752), .A4(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n713), .B1(new_n737), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n707), .A2(new_n700), .A3(new_n715), .A4(new_n756), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n702), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(G396));
  INV_X1    g0559(.A(KEYINPUT96), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n366), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n359), .A2(new_n363), .A3(KEYINPUT96), .A4(new_n365), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n642), .A2(new_n348), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n763), .A2(new_n430), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(KEYINPUT97), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n366), .A2(new_n764), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT97), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n763), .A2(new_n768), .A3(new_n430), .A4(new_n764), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n666), .B(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(new_n695), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n701), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n770), .A2(new_n705), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n735), .A2(new_n447), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n732), .A2(KEYINPUT95), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n732), .A2(KEYINPUT95), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n725), .A2(new_n751), .B1(new_n778), .B2(new_n741), .ZN(new_n779));
  INV_X1    g0579(.A(new_n726), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n775), .B(new_n779), .C1(G116), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n729), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G311), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n263), .B1(new_n721), .B2(G303), .ZN(new_n784));
  INV_X1    g0584(.A(new_n717), .ZN(new_n785));
  INV_X1    g0585(.A(new_n733), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n785), .A2(G107), .B1(new_n786), .B2(G97), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n781), .A2(new_n783), .A3(new_n784), .A4(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G143), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n726), .A2(new_n368), .B1(new_n725), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G137), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n791), .B1(new_n792), .B2(new_n720), .C1(new_n323), .C2(new_n732), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT34), .ZN(new_n794));
  INV_X1    g0594(.A(new_n735), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n785), .A2(G50), .B1(new_n795), .B2(G68), .ZN(new_n796));
  INV_X1    g0596(.A(new_n387), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(G132), .B2(new_n782), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n794), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n733), .A2(new_n202), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n788), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n713), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n713), .A2(new_n704), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n211), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n774), .A2(new_n700), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n773), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(G384));
  NAND3_X1  g0607(.A1(new_n420), .A2(new_n427), .A3(new_n421), .ZN(new_n808));
  INV_X1    g0608(.A(new_n640), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n373), .B1(new_n380), .B2(new_n381), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT101), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n390), .A2(KEYINPUT101), .A3(new_n373), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n812), .A2(new_n393), .A3(new_n813), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n814), .A2(new_n299), .A3(new_n383), .A4(new_n392), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n809), .B1(new_n815), .B2(new_n404), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n808), .A2(new_n816), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n815), .A2(new_n404), .B1(new_n425), .B2(new_n809), .ZN(new_n818));
  INV_X1    g0618(.A(new_n414), .ZN(new_n819));
  OAI21_X1  g0619(.A(KEYINPUT37), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT102), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n402), .A2(new_n404), .ZN(new_n823));
  INV_X1    g0623(.A(new_n425), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n640), .ZN(new_n826));
  XOR2_X1   g0626(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n825), .A2(new_n826), .A3(new_n414), .A4(new_n828), .ZN(new_n829));
  OAI211_X1 g0629(.A(KEYINPUT102), .B(KEYINPUT37), .C1(new_n818), .C2(new_n819), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n822), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  AND3_X1   g0631(.A1(new_n817), .A2(new_n831), .A3(KEYINPUT38), .ZN(new_n832));
  AOI21_X1  g0632(.A(KEYINPUT38), .B1(new_n817), .B2(new_n831), .ZN(new_n833));
  OAI21_X1  g0633(.A(KEYINPUT104), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n817), .A2(new_n831), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT38), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT104), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n817), .A2(new_n831), .A3(KEYINPUT38), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n691), .A2(new_n693), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n642), .A2(new_n312), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n313), .A2(new_n320), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n290), .A2(new_n312), .A3(new_n642), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND3_X1   g0645(.A1(new_n841), .A2(new_n770), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n834), .A2(new_n840), .A3(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT40), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n418), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n826), .B1(new_n427), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT107), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n829), .B(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT106), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n825), .A2(new_n854), .A3(new_n414), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n826), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n854), .B1(new_n825), .B2(new_n414), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n827), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n851), .B1(new_n853), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n839), .B1(new_n859), .B2(KEYINPUT38), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n860), .A2(KEYINPUT40), .A3(new_n846), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n849), .A2(G330), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n432), .A2(new_n694), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n861), .B1(new_n847), .B2(new_n848), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n866), .A2(new_n432), .A3(new_n841), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT108), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n667), .A2(new_n677), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n611), .B1(new_n870), .B2(new_n432), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n869), .B(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n845), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n641), .B(new_n770), .C1(new_n620), .C2(new_n632), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n763), .A2(new_n642), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n873), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(new_n834), .A3(new_n840), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT39), .B1(new_n832), .B2(new_n833), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT39), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n839), .B(new_n880), .C1(new_n859), .C2(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n290), .A2(new_n312), .A3(new_n641), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT105), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n609), .A2(new_n809), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n878), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n872), .B(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n247), .B2(new_n635), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n371), .A2(new_n230), .A3(G77), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n892), .B(KEYINPUT100), .Z(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n203), .B2(new_n201), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(G1), .A3(new_n293), .ZN(new_n895));
  OAI211_X1 g0695(.A(G116), .B(new_n228), .C1(new_n475), .C2(KEYINPUT35), .ZN(new_n896));
  XOR2_X1   g0696(.A(new_n896), .B(KEYINPUT98), .Z(new_n897));
  NAND2_X1  g0697(.A1(new_n475), .A2(KEYINPUT35), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g0699(.A(KEYINPUT99), .B(KEYINPUT36), .Z(new_n900));
  XNOR2_X1  g0700(.A(new_n899), .B(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n891), .A2(new_n895), .A3(new_n901), .ZN(G367));
  NAND2_X1  g0702(.A1(new_n625), .A2(new_n642), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n674), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n657), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT42), .Z(new_n906));
  NAND3_X1  g0706(.A1(new_n674), .A2(new_n573), .A3(new_n903), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n642), .B1(new_n907), .B2(new_n510), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT43), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n469), .A2(new_n524), .ZN(new_n910));
  INV_X1    g0710(.A(new_n519), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n642), .B1(new_n911), .B2(new_n522), .ZN(new_n912));
  MUX2_X1   g0712(.A(new_n469), .B(new_n910), .S(new_n912), .Z(new_n913));
  OAI22_X1  g0713(.A1(new_n906), .A2(new_n908), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n909), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n914), .B(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n904), .B1(new_n510), .B2(new_n641), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n654), .A2(new_n918), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n916), .B(new_n919), .Z(new_n920));
  XNOR2_X1  g0720(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n660), .B(new_n921), .Z(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n657), .A2(new_n655), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n924), .A2(new_n918), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT45), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n918), .ZN(new_n927));
  XOR2_X1   g0727(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n928));
  XNOR2_X1  g0728(.A(new_n927), .B(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT111), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n932), .A2(new_n654), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n657), .B1(new_n653), .B2(new_n656), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n648), .B(new_n934), .Z(new_n935));
  NOR2_X1   g0735(.A1(new_n935), .A2(new_n696), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n932), .A2(new_n654), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n933), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n923), .B1(new_n938), .B2(new_n697), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n247), .B1(new_n635), .B2(G45), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n920), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n733), .A2(new_n203), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n778), .A2(new_n368), .B1(new_n789), .B2(new_n720), .ZN(new_n944));
  INV_X1    g0744(.A(new_n725), .ZN(new_n945));
  AOI211_X1 g0745(.A(new_n943), .B(new_n944), .C1(G150), .C2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n201), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n263), .B1(new_n211), .B2(new_n735), .C1(new_n726), .C2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n717), .A2(new_n202), .B1(new_n792), .B2(new_n729), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT112), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n946), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n785), .A2(G116), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT46), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n953), .A2(new_n954), .B1(new_n746), .B2(new_n729), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n797), .B1(new_n725), .B2(new_n753), .C1(new_n741), .C2(new_n726), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n955), .B(new_n956), .C1(G97), .C2(new_n795), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n953), .A2(new_n954), .B1(G107), .B2(new_n786), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n957), .B(new_n958), .C1(new_n751), .C2(new_n778), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n720), .A2(new_n738), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n952), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT113), .Z(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT47), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n713), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n913), .A2(new_n706), .ZN(new_n965));
  INV_X1    g0765(.A(new_n710), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n714), .B1(new_n208), .B2(new_n344), .C1(new_n966), .C2(new_n238), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n964), .A2(new_n700), .A3(new_n965), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n942), .A2(new_n968), .ZN(G387));
  AND2_X1   g0769(.A1(new_n935), .A2(new_n696), .ZN(new_n970));
  OR3_X1    g0770(.A1(new_n970), .A2(new_n936), .A3(new_n661), .ZN(new_n971));
  INV_X1    g0771(.A(new_n778), .ZN(new_n972));
  AOI22_X1  g0772(.A1(G317), .A2(new_n945), .B1(new_n972), .B2(G311), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n973), .B1(new_n753), .B2(new_n726), .C1(new_n739), .C2(new_n720), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT48), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n975), .B1(new_n741), .B2(new_n733), .C1(new_n751), .C2(new_n717), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT49), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n387), .B1(new_n976), .B2(new_n977), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n782), .A2(G326), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G116), .B2(new_n795), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n785), .A2(G77), .B1(new_n795), .B2(G97), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n725), .B2(new_n306), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n720), .A2(new_n368), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n732), .A2(new_n324), .ZN(new_n986));
  NOR4_X1   g0786(.A1(new_n984), .A2(new_n797), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n786), .A2(new_n435), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(new_n323), .C2(new_n729), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G68), .B2(new_n780), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n713), .B1(new_n982), .B2(new_n990), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n652), .B(new_n706), .C1(new_n649), .C2(new_n641), .ZN(new_n992));
  INV_X1    g0792(.A(new_n324), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n306), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n663), .B1(new_n994), .B2(KEYINPUT50), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n995), .B(new_n457), .C1(KEYINPUT50), .C2(new_n994), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(G68), .B2(G77), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n710), .B1(new_n235), .B2(new_n248), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n263), .A2(new_n663), .A3(new_n208), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n208), .A2(G107), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n714), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n991), .A2(new_n700), .A3(new_n992), .A4(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT114), .Z(new_n1004));
  OAI211_X1 g0804(.A(new_n971), .B(new_n1004), .C1(new_n940), .C2(new_n935), .ZN(G393));
  XNOR2_X1  g0805(.A(new_n930), .B(new_n654), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n938), .B(new_n660), .C1(new_n936), .C2(new_n1006), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n714), .B1(new_n442), .B2(new_n208), .C1(new_n966), .C2(new_n242), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n725), .A2(new_n738), .B1(new_n746), .B2(new_n720), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n736), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n780), .A2(G294), .B1(new_n972), .B2(G303), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n717), .A2(new_n741), .B1(new_n733), .B2(new_n460), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n263), .B(new_n1014), .C1(G322), .C2(new_n782), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n725), .A2(new_n368), .B1(new_n323), .B2(new_n720), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT51), .Z(new_n1018));
  AOI211_X1 g0818(.A(new_n797), .B(new_n1018), .C1(new_n993), .C2(new_n780), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n733), .A2(new_n211), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1020), .B(new_n775), .C1(G68), .C2(new_n785), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1019), .B(new_n1021), .C1(new_n947), .C2(new_n778), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n729), .A2(new_n789), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1016), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n713), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n918), .A2(new_n706), .ZN(new_n1026));
  AND3_X1   g0826(.A1(new_n1025), .A2(new_n1026), .A3(new_n700), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n1006), .A2(new_n941), .B1(new_n1008), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1007), .A2(new_n1028), .ZN(G390));
  NAND2_X1  g0829(.A1(new_n694), .A2(new_n770), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT116), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n845), .B1(new_n1031), .B2(new_n770), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n676), .A2(new_n770), .A3(new_n641), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1036), .A2(new_n876), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1030), .A2(new_n873), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n694), .A2(new_n770), .A3(new_n845), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n874), .A2(new_n876), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n1035), .A2(new_n1037), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n612), .B(new_n864), .C1(new_n678), .C2(new_n433), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n879), .B(new_n881), .C1(new_n877), .C2(new_n885), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n884), .B(new_n860), .C1(new_n1037), .C2(new_n873), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1039), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n885), .B1(new_n1041), .B2(new_n845), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1039), .B(new_n1047), .C1(new_n1049), .C2(new_n882), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1045), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1039), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1044), .A2(new_n1055), .A3(new_n1050), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1052), .A2(new_n660), .A3(new_n1056), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT117), .Z(new_n1058));
  NAND3_X1  g0858(.A1(new_n879), .A2(new_n704), .A3(new_n881), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n803), .A2(new_n324), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n726), .A2(new_n442), .B1(new_n778), .B2(new_n213), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G116), .B2(new_n945), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n395), .B1(new_n733), .B2(new_n211), .C1(new_n720), .C2(new_n741), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n718), .B(new_n1064), .C1(G294), .C2(new_n782), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1063), .B(new_n1065), .C1(new_n203), .C2(new_n735), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(KEYINPUT54), .B(G143), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT118), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n780), .A2(new_n1068), .B1(G128), .B2(new_n721), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n778), .A2(new_n792), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G132), .B2(new_n945), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n263), .B1(new_n947), .B2(new_n735), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT119), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n786), .A2(G159), .B1(new_n782), .B2(G125), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1069), .A2(new_n1071), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n785), .A2(G150), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT53), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1066), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n701), .B(new_n1061), .C1(new_n713), .C2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1051), .A2(new_n1048), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1079), .B1(new_n1080), .B2(new_n941), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1058), .A2(new_n1081), .ZN(G378));
  INV_X1    g0882(.A(KEYINPUT122), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT121), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n834), .A2(new_n840), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1085), .A2(new_n877), .B1(new_n609), .B2(new_n809), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1084), .B1(new_n1086), .B2(new_n886), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n338), .A2(new_n341), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n327), .A2(new_n640), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1088), .B(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1090), .B(new_n1092), .ZN(new_n1093));
  AND4_X1   g0893(.A1(G330), .A2(new_n849), .A3(new_n1093), .A4(new_n862), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1093), .B1(new_n866), .B2(G330), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1087), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1093), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n863), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n888), .A2(KEYINPUT121), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n866), .A2(G330), .A3(new_n1093), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1096), .A2(new_n1101), .A3(new_n941), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n701), .B1(new_n1093), .B2(new_n704), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n721), .A2(G125), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n780), .A2(G137), .B1(G132), .B2(new_n745), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1068), .A2(new_n785), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT120), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1105), .B(new_n1107), .C1(new_n323), .C2(new_n733), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1104), .B(new_n1108), .C1(G128), .C2(new_n945), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT59), .ZN(new_n1110));
  AOI21_X1  g0910(.A(G33), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(G41), .B1(new_n782), .B2(G124), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1111), .B(new_n1112), .C1(new_n368), .C2(new_n735), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1114));
  AOI21_X1  g0914(.A(G41), .B1(new_n384), .B2(KEYINPUT3), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1113), .A2(new_n1114), .B1(G50), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n797), .B1(new_n460), .B2(new_n720), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n945), .A2(G107), .B1(G97), .B2(new_n745), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n741), .B2(new_n729), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1117), .B(new_n1119), .C1(new_n435), .C2(new_n780), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n735), .A2(new_n202), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n943), .B(new_n1121), .C1(G77), .C2(new_n785), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1120), .A2(new_n252), .A3(new_n1122), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT58), .Z(new_n1124));
  OAI21_X1  g0924(.A(new_n713), .B1(new_n1116), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n803), .A2(new_n947), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1103), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1102), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n888), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1098), .A2(new_n889), .A3(new_n1100), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT57), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1043), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1132), .B1(new_n1056), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n661), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1096), .A2(new_n1101), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1043), .B1(new_n1080), .B2(new_n1044), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1132), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1083), .B(new_n1128), .C1(new_n1135), .C2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1056), .A2(new_n1133), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1140), .A2(KEYINPUT57), .A3(new_n1130), .A4(new_n1129), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1138), .A2(new_n660), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1128), .ZN(new_n1143));
  AOI21_X1  g0943(.A(KEYINPUT122), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1139), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(G375));
  NAND2_X1  g0946(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1045), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1148), .A2(new_n923), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT123), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n873), .A2(new_n704), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1121), .B1(new_n780), .B2(G150), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n721), .A2(G132), .B1(new_n786), .B2(G50), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1152), .A2(new_n387), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n972), .A2(new_n1068), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1155), .B1(new_n792), .B2(new_n725), .C1(new_n368), .C2(new_n717), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1154), .B(new_n1156), .C1(G128), .C2(new_n782), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n780), .A2(G107), .B1(new_n972), .B2(G116), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n741), .B2(new_n725), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n729), .A2(new_n753), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n988), .B(new_n395), .C1(new_n751), .C2(new_n720), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n735), .A2(new_n211), .B1(new_n717), .B2(new_n442), .ZN(new_n1162));
  NOR4_X1   g0962(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n713), .B1(new_n1157), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n803), .A2(new_n203), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1151), .A2(new_n700), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n1042), .B2(new_n940), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1150), .A2(new_n1168), .ZN(G381));
  AND2_X1   g0969(.A1(new_n1057), .A2(new_n1081), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1145), .A2(new_n1170), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1171), .A2(G384), .A3(G381), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n942), .A2(new_n968), .A3(new_n1028), .A4(new_n1007), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1173), .A2(G396), .A3(G393), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(G407));
  OAI211_X1 g0975(.A(G407), .B(G213), .C1(G343), .C2(new_n1171), .ZN(G409));
  NAND2_X1  g0976(.A1(G387), .A2(G390), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n1173), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(G393), .B(new_n758), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1178), .B(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1128), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1131), .A2(new_n941), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n1127), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT124), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1140), .A2(new_n922), .A3(new_n1101), .A4(new_n1096), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1182), .A2(KEYINPUT124), .A3(new_n1127), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(G378), .A2(new_n1181), .B1(new_n1188), .B2(new_n1170), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1148), .A2(KEYINPUT60), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1147), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1191), .B(new_n660), .C1(KEYINPUT60), .C2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n1168), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n806), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(G384), .A3(new_n1168), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(G213), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1199), .A2(G343), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1190), .A2(new_n1198), .A3(new_n1201), .ZN(new_n1202));
  XOR2_X1   g1002(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n1203));
  NOR2_X1   g1003(.A1(new_n1189), .A2(new_n1200), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1200), .A2(G2897), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1197), .B(new_n1206), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n1202), .A2(new_n1203), .B1(new_n1204), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT61), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1189), .A2(new_n1197), .A3(new_n1200), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT125), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(KEYINPUT62), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1209), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1180), .B1(new_n1208), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(KEYINPUT63), .B1(new_n1204), .B2(new_n1207), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n1202), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1180), .B1(new_n1210), .B2(KEYINPUT63), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n1209), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1214), .A2(new_n1218), .ZN(G405));
  OAI21_X1  g1019(.A(new_n1170), .B1(new_n1139), .B2(new_n1144), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(KEYINPUT126), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(G378), .A2(new_n1181), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT126), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1223), .B(new_n1170), .C1(new_n1139), .C2(new_n1144), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1221), .A2(new_n1222), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n1197), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1179), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1178), .B(new_n1227), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1221), .A2(new_n1198), .A3(new_n1222), .A4(new_n1224), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1226), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(KEYINPUT127), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1226), .A2(new_n1229), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n1180), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT127), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1226), .A2(new_n1234), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1231), .A2(new_n1233), .A3(new_n1235), .ZN(G402));
endmodule


