//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  INV_X1    g000(.A(KEYINPUT26), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n206));
  AND3_X1   g005(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n205), .B(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT68), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT68), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n209), .A2(new_n213), .A3(new_n210), .ZN(new_n214));
  INV_X1    g013(.A(G183gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT27), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT27), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G183gat), .ZN(new_n218));
  INV_X1    g017(.A(G190gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT28), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(new_n222), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT27), .B(G183gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(KEYINPUT28), .A3(new_n219), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n226), .A3(KEYINPUT67), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n212), .A2(new_n214), .A3(new_n223), .A4(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT25), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(new_n203), .A3(new_n204), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(new_n208), .B2(new_n207), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n210), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n215), .A2(new_n219), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n229), .B1(new_n234), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n208), .ZN(new_n241));
  NAND3_X1  g040(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n241), .A2(new_n242), .B1(new_n231), .B2(new_n232), .ZN(new_n243));
  AND3_X1   g042(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n245));
  NOR3_X1   g044(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT24), .ZN(new_n246));
  OR3_X1    g045(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n237), .A3(new_n248), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n243), .B(KEYINPUT25), .C1(new_n246), .C2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n240), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n228), .A2(new_n251), .ZN(new_n252));
  AND2_X1   g051(.A1(G226gat), .A2(G233gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT29), .B1(new_n228), .B2(new_n251), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n254), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(G211gat), .A2(G218gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(G211gat), .A2(G218gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G197gat), .B(G204gat), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n260), .B(new_n261), .C1(KEYINPUT22), .C2(new_n257), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(KEYINPUT22), .B2(new_n257), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n259), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n256), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G8gat), .B(G36gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(G64gat), .B(G92gat), .ZN(new_n268));
  XOR2_X1   g067(.A(new_n267), .B(new_n268), .Z(new_n269));
  INV_X1    g068(.A(new_n265), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n254), .B(new_n270), .C1(new_n253), .C2(new_n255), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n266), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT74), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT74), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n266), .A2(new_n274), .A3(new_n269), .A4(new_n271), .ZN(new_n275));
  XOR2_X1   g074(.A(KEYINPUT75), .B(KEYINPUT30), .Z(new_n276));
  NAND3_X1  g075(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n269), .B1(new_n266), .B2(new_n271), .ZN(new_n278));
  INV_X1    g077(.A(new_n272), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n278), .B1(new_n279), .B2(KEYINPUT30), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(G113gat), .B(G120gat), .Z(new_n282));
  INV_X1    g081(.A(KEYINPUT1), .ZN(new_n283));
  INV_X1    g082(.A(G134gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G127gat), .ZN(new_n285));
  INV_X1    g084(.A(G127gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G134gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n282), .B(new_n283), .C1(KEYINPUT70), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(KEYINPUT69), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G113gat), .B(G120gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT70), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT1), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n285), .A2(new_n287), .A3(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G141gat), .B(G148gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G155gat), .ZN(new_n301));
  INV_X1    g100(.A(G162gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(KEYINPUT2), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n300), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n304), .B(new_n303), .C1(new_n299), .C2(KEYINPUT2), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT3), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n308), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT3), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n298), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G225gat), .A2(G233gat), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n289), .B(new_n290), .C1(new_n294), .C2(new_n296), .ZN(new_n316));
  INV_X1    g115(.A(new_n311), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT76), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT76), .B1(new_n316), .B2(new_n317), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT4), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT5), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n316), .A2(new_n317), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT4), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n315), .A2(new_n320), .A3(new_n321), .A4(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n316), .A2(new_n317), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n318), .A2(new_n319), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT5), .B1(new_n327), .B2(new_n314), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n318), .A2(new_n319), .A3(KEYINPUT4), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT4), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n313), .A2(new_n314), .A3(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n325), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G1gat), .B(G29gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(KEYINPUT0), .ZN(new_n335));
  XNOR2_X1  g134(.A(G57gat), .B(G85gat), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n335), .B(new_n336), .Z(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n333), .A2(KEYINPUT6), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n333), .A2(new_n338), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT6), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n337), .B(new_n325), .C1(new_n328), .C2(new_n332), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n281), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT71), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n228), .A2(new_n298), .A3(new_n251), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n298), .B1(new_n228), .B2(new_n251), .ZN(new_n349));
  INV_X1    g148(.A(G227gat), .ZN(new_n350));
  INV_X1    g149(.A(G233gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NOR3_X1   g152(.A1(new_n348), .A2(new_n349), .A3(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n347), .B1(new_n354), .B2(KEYINPUT33), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n252), .A2(new_n316), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n228), .A2(new_n298), .A3(new_n251), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(new_n352), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT33), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(KEYINPUT71), .A3(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G15gat), .B(G43gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(G71gat), .B(G99gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n363), .B1(new_n358), .B2(KEYINPUT32), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n355), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT34), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n356), .A2(new_n357), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n366), .B1(new_n367), .B2(new_n353), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n366), .B(new_n353), .C1(new_n348), .C2(new_n349), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n358), .B(KEYINPUT32), .C1(new_n359), .C2(new_n363), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n365), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n371), .B1(new_n365), .B2(new_n372), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT31), .B(G50gat), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT29), .B1(new_n262), .B2(new_n264), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n311), .B1(new_n377), .B2(KEYINPUT3), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT78), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT78), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n380), .B(new_n311), .C1(new_n377), .C2(KEYINPUT3), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT29), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n310), .A2(new_n382), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n383), .A2(new_n265), .B1(G228gat), .B2(G233gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n379), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G228gat), .A2(G233gat), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT79), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n310), .A2(KEYINPUT79), .A3(new_n382), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n265), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n387), .B1(new_n391), .B2(new_n378), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n376), .B1(new_n386), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n376), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n391), .A2(new_n378), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n385), .B(new_n394), .C1(new_n395), .C2(new_n387), .ZN(new_n396));
  XNOR2_X1  g195(.A(G78gat), .B(G106gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT77), .ZN(new_n398));
  INV_X1    g197(.A(G22gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n393), .A2(new_n396), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n400), .B1(new_n393), .B2(new_n396), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n375), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT35), .B1(new_n346), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n364), .A2(new_n360), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT71), .B1(new_n358), .B2(new_n359), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n372), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n371), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n365), .A2(new_n371), .A3(new_n372), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n413), .A2(new_n403), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT35), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n414), .A2(new_n415), .A3(new_n345), .A4(new_n281), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n406), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n343), .A2(new_n342), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT76), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n322), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT76), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n298), .A2(new_n311), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n314), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n321), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n425), .B1(new_n329), .B2(new_n331), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n337), .B1(new_n426), .B2(new_n325), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n418), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(new_n339), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n277), .A2(new_n280), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n403), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT73), .ZN(new_n432));
  XOR2_X1   g231(.A(KEYINPUT72), .B(KEYINPUT36), .Z(new_n433));
  OAI211_X1 g232(.A(new_n432), .B(new_n433), .C1(new_n373), .C2(new_n374), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n411), .A2(KEYINPUT36), .A3(new_n412), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n432), .B1(new_n413), .B2(new_n433), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n431), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT39), .B1(new_n423), .B2(new_n424), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n320), .A2(new_n313), .A3(new_n324), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n440), .B1(new_n442), .B2(new_n314), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT39), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n444), .A3(new_n424), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n443), .A2(KEYINPUT40), .A3(new_n337), .A4(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT40), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n337), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n439), .B1(new_n424), .B2(new_n441), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n446), .A2(new_n450), .A3(new_n341), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT81), .B1(new_n281), .B2(new_n451), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n450), .A2(new_n341), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT81), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n453), .A2(new_n430), .A3(new_n454), .A4(new_n446), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n273), .A2(new_n275), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n428), .A2(new_n339), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n266), .A2(new_n271), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n269), .B1(new_n459), .B2(KEYINPUT37), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT38), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT37), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n266), .A2(new_n462), .A3(new_n271), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n460), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n461), .B1(new_n460), .B2(new_n463), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n403), .B1(new_n458), .B2(new_n466), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n438), .A2(KEYINPUT80), .B1(new_n456), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT80), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n431), .B(new_n469), .C1(new_n436), .C2(new_n437), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n417), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT96), .ZN(new_n473));
  OR2_X1    g272(.A1(G71gat), .A2(G78gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(G71gat), .A2(G78gat), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(KEYINPUT87), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT87), .ZN(new_n477));
  AND2_X1   g276(.A1(G71gat), .A2(G78gat), .ZN(new_n478));
  NOR2_X1   g277(.A1(G71gat), .A2(G78gat), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n478), .A2(KEYINPUT9), .ZN(new_n481));
  XNOR2_X1  g280(.A(G57gat), .B(G64gat), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n476), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT88), .ZN(new_n484));
  AND2_X1   g283(.A1(KEYINPUT89), .A2(G64gat), .ZN(new_n485));
  NOR2_X1   g284(.A1(KEYINPUT89), .A2(G64gat), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n484), .B(G57gat), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT9), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n475), .B1(new_n474), .B2(new_n488), .ZN(new_n489));
  OR2_X1    g288(.A1(KEYINPUT89), .A2(G64gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n484), .A2(G57gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(KEYINPUT89), .A2(G64gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n487), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n483), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT90), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT21), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n483), .A2(new_n494), .A3(KEYINPUT90), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G127gat), .B(G155gat), .ZN(new_n501));
  XOR2_X1   g300(.A(new_n500), .B(new_n501), .Z(new_n502));
  AND3_X1   g301(.A1(new_n483), .A2(new_n494), .A3(KEYINPUT90), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT90), .B1(new_n483), .B2(new_n494), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT91), .ZN(new_n505));
  NOR3_X1   g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT91), .B1(new_n497), .B2(new_n499), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT21), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n399), .A2(G15gat), .ZN(new_n509));
  INV_X1    g308(.A(G15gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(G22gat), .ZN(new_n511));
  INV_X1    g310(.A(G1gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT16), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n509), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G8gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n514), .B(new_n515), .C1(G1gat), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT85), .ZN(new_n518));
  AOI21_X1  g317(.A(G1gat), .B1(new_n509), .B2(new_n511), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT85), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n520), .A2(new_n521), .A3(new_n515), .A4(new_n514), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT83), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n515), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n514), .B(KEYINPUT83), .C1(G1gat), .C2(new_n516), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n525), .A2(new_n526), .A3(KEYINPUT84), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT84), .B1(new_n525), .B2(new_n526), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n523), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n508), .A2(new_n530), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n502), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n502), .A2(new_n531), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n535));
  NAND2_X1  g334(.A1(G231gat), .A2(G233gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G183gat), .B(G211gat), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n537), .B(new_n538), .Z(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n534), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n532), .A2(new_n533), .A3(new_n539), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G190gat), .B(G218gat), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G29gat), .ZN(new_n547));
  INV_X1    g346(.A(G36gat), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT14), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT14), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(G29gat), .B2(G36gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(G29gat), .A2(G36gat), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT15), .ZN(new_n554));
  INV_X1    g353(.A(G43gat), .ZN(new_n555));
  INV_X1    g354(.A(G50gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G43gat), .A2(G50gat), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n553), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n558), .ZN(new_n561));
  NOR2_X1   g360(.A1(G43gat), .A2(G50gat), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT15), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n557), .A2(new_n554), .A3(new_n558), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n560), .B(KEYINPUT82), .C1(new_n565), .C2(new_n553), .ZN(new_n566));
  INV_X1    g365(.A(new_n553), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT82), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n567), .A2(new_n568), .A3(new_n563), .A4(new_n564), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT17), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT17), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n566), .A2(new_n572), .A3(new_n569), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT8), .ZN(new_n574));
  NAND2_X1  g373(.A1(G99gat), .A2(G106gat), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n574), .B1(new_n575), .B2(KEYINPUT93), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT93), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n577), .A2(G99gat), .A3(G106gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(G92gat), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n580), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n581));
  INV_X1    g380(.A(G92gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n579), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n575), .ZN(new_n586));
  NOR2_X1   g385(.A1(G99gat), .A2(G106gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT7), .ZN(new_n590));
  INV_X1    g389(.A(G85gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(G92gat), .A3(new_n593), .ZN(new_n594));
  AOI22_X1  g393(.A1(new_n594), .A2(new_n583), .B1(new_n576), .B2(new_n578), .ZN(new_n595));
  INV_X1    g394(.A(new_n588), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n589), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n571), .A2(new_n573), .A3(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n566), .A2(new_n569), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n589), .A2(new_n597), .ZN(new_n601));
  NAND2_X1  g400(.A1(G232gat), .A2(G233gat), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI22_X1  g402(.A1(new_n600), .A2(new_n601), .B1(KEYINPUT41), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n546), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n603), .A2(KEYINPUT41), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT92), .ZN(new_n608));
  XNOR2_X1  g407(.A(G134gat), .B(G162gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  NAND3_X1  g409(.A1(new_n599), .A2(new_n604), .A3(new_n546), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n606), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT94), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n611), .B1(new_n605), .B2(new_n614), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n599), .A2(new_n604), .A3(KEYINPUT94), .A4(new_n546), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n610), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n613), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI211_X1 g418(.A(KEYINPUT95), .B(new_n610), .C1(new_n615), .C2(new_n616), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n612), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n473), .B1(new_n544), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n612), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n617), .A2(new_n618), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT95), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n617), .A2(new_n613), .A3(new_n618), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n627), .A2(KEYINPUT96), .A3(new_n543), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n622), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G113gat), .B(G141gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G197gat), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT11), .B(G169gat), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  NAND2_X1  g433(.A1(new_n525), .A2(new_n526), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT84), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n525), .A2(new_n526), .A3(KEYINPUT84), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n571), .A2(new_n639), .A3(new_n523), .A4(new_n573), .ZN(new_n640));
  NAND2_X1  g439(.A1(G229gat), .A2(G233gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n529), .A2(new_n600), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(KEYINPUT86), .A2(KEYINPUT18), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n641), .B(KEYINPUT13), .Z(new_n646));
  NOR2_X1   g445(.A1(new_n529), .A2(new_n600), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n570), .B1(new_n639), .B2(new_n523), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n644), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n640), .A2(new_n641), .A3(new_n642), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n634), .B1(new_n645), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n643), .A2(new_n644), .ZN(new_n654));
  INV_X1    g453(.A(new_n634), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n654), .A2(new_n655), .A3(new_n649), .A4(new_n651), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G120gat), .B(G148gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(G176gat), .B(G204gat), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n659), .B(new_n660), .Z(new_n661));
  NAND2_X1  g460(.A1(G230gat), .A2(G233gat), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n598), .A2(new_n497), .A3(new_n499), .ZN(new_n663));
  INV_X1    g462(.A(new_n495), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT97), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n665), .B1(new_n586), .B2(new_n587), .ZN(new_n666));
  INV_X1    g465(.A(G99gat), .ZN(new_n667));
  INV_X1    g466(.A(G106gat), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n669), .A2(KEYINPUT97), .A3(new_n575), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT98), .B1(new_n595), .B2(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n666), .A2(new_n670), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT98), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n585), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n664), .A2(new_n672), .A3(new_n675), .A4(new_n597), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT10), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n663), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n589), .A2(KEYINPUT10), .A3(new_n597), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n505), .B1(new_n503), .B2(new_n504), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n497), .A2(KEYINPUT91), .A3(new_n499), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n662), .B1(new_n678), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n663), .A2(new_n676), .ZN(new_n684));
  INV_X1    g483(.A(new_n662), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n661), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n683), .A2(new_n686), .A3(new_n661), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n629), .A2(new_n658), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n472), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n345), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(new_n512), .ZN(G1324gat));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n695));
  INV_X1    g494(.A(new_n692), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n430), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT99), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT16), .B(G8gat), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n695), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(G8gat), .ZN(new_n702));
  OR3_X1    g501(.A1(new_n697), .A2(new_n695), .A3(new_n700), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(G1325gat));
  NOR2_X1   g503(.A1(new_n436), .A2(new_n437), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G15gat), .B1(new_n692), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n375), .A2(new_n510), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n707), .B1(new_n692), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT100), .ZN(G1326gat));
  NOR2_X1   g509(.A1(new_n692), .A2(new_n404), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT43), .B(G22gat), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  NOR2_X1   g512(.A1(new_n658), .A2(new_n690), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n544), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n471), .A2(new_n627), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n716), .A2(new_n547), .A3(new_n429), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT45), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT44), .B1(new_n471), .B2(new_n627), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n406), .A2(new_n416), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n456), .A2(new_n467), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n720), .B1(new_n721), .B2(new_n438), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n722), .A2(new_n723), .A3(new_n621), .ZN(new_n724));
  AOI211_X1 g523(.A(KEYINPUT101), .B(new_n715), .C1(new_n719), .C2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT101), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n438), .A2(KEYINPUT80), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n456), .A2(new_n467), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n727), .A2(new_n470), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n627), .B1(new_n729), .B2(new_n720), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n724), .B1(new_n730), .B2(new_n723), .ZN(new_n731));
  INV_X1    g530(.A(new_n715), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n726), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n725), .A2(new_n733), .A3(new_n345), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n718), .B1(new_n734), .B2(new_n547), .ZN(G1328gat));
  NOR2_X1   g534(.A1(new_n725), .A2(new_n733), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n548), .B1(new_n736), .B2(new_n430), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT102), .ZN(new_n738));
  AOI21_X1  g537(.A(G36gat), .B1(new_n738), .B2(KEYINPUT46), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n716), .A2(new_n430), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n738), .A2(KEYINPUT46), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT103), .B1(new_n737), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n725), .A2(new_n733), .A3(new_n281), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n742), .B(new_n745), .C1(new_n746), .C2(new_n548), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n747), .ZN(G1329gat));
  INV_X1    g547(.A(new_n716), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n749), .A2(G43gat), .A3(new_n413), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n731), .A2(new_n732), .ZN(new_n752));
  OAI21_X1  g551(.A(G43gat), .B1(new_n752), .B2(new_n706), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n751), .A2(KEYINPUT47), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n736), .A2(new_n705), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n750), .B1(new_n755), .B2(G43gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n756), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g556(.A(G50gat), .B1(new_n752), .B2(new_n404), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n716), .A2(KEYINPUT105), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n716), .A2(KEYINPUT105), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(new_n556), .A3(new_n403), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n758), .B(KEYINPUT48), .C1(new_n759), .C2(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n759), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n736), .A2(new_n403), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n764), .B2(G50gat), .ZN(new_n765));
  XOR2_X1   g564(.A(KEYINPUT104), .B(KEYINPUT48), .Z(new_n766));
  OAI21_X1  g565(.A(new_n762), .B1(new_n765), .B2(new_n766), .ZN(G1331gat));
  INV_X1    g566(.A(new_n690), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n629), .A2(new_n657), .A3(new_n768), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n722), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n429), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n430), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n774));
  XOR2_X1   g573(.A(KEYINPUT49), .B(G64gat), .Z(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT106), .ZN(G1333gat));
  NAND2_X1  g576(.A1(new_n770), .A2(new_n705), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n413), .A2(G71gat), .ZN(new_n779));
  AOI22_X1  g578(.A1(new_n778), .A2(G71gat), .B1(new_n770), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g580(.A1(new_n770), .A2(new_n403), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g582(.A1(new_n543), .A2(new_n657), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n690), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n719), .B2(new_n724), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(G85gat), .B1(new_n787), .B2(new_n345), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n722), .A2(new_n621), .A3(new_n784), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT51), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n345), .A2(G85gat), .A3(new_n768), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT107), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n788), .B1(new_n790), .B2(new_n792), .ZN(G1336gat));
  AOI21_X1  g592(.A(new_n582), .B1(new_n786), .B2(new_n430), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n722), .A2(new_n621), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT108), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n796), .A3(new_n784), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n789), .A2(KEYINPUT108), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT109), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n795), .A2(KEYINPUT51), .A3(new_n784), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n797), .A2(KEYINPUT109), .A3(new_n798), .A4(new_n799), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n281), .A2(G92gat), .A3(new_n768), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n794), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808));
  INV_X1    g607(.A(new_n806), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n808), .B1(new_n790), .B2(new_n809), .ZN(new_n810));
  OAI22_X1  g609(.A1(new_n807), .A2(new_n808), .B1(new_n794), .B2(new_n810), .ZN(G1337gat));
  OAI21_X1  g610(.A(G99gat), .B1(new_n787), .B2(new_n706), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n375), .A2(new_n667), .A3(new_n690), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n812), .B1(new_n790), .B2(new_n813), .ZN(G1338gat));
  AOI21_X1  g613(.A(new_n668), .B1(new_n786), .B2(new_n403), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n404), .A2(G106gat), .A3(new_n768), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n815), .B1(new_n805), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818));
  INV_X1    g617(.A(new_n816), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n818), .B1(new_n790), .B2(new_n819), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n817), .A2(new_n818), .B1(new_n815), .B2(new_n820), .ZN(G1339gat));
  INV_X1    g620(.A(KEYINPUT111), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n647), .A2(new_n648), .A3(new_n646), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n641), .B1(new_n640), .B2(new_n642), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n633), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n689), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n656), .B(new_n825), .C1(new_n826), .C2(new_n687), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828));
  INV_X1    g627(.A(new_n679), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n506), .B2(new_n507), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n663), .A2(new_n676), .A3(new_n677), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(new_n831), .A3(new_n685), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n683), .A2(KEYINPUT54), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n661), .ZN(new_n834));
  XNOR2_X1  g633(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n834), .B1(new_n683), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n828), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n685), .B1(new_n830), .B2(new_n831), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n661), .B1(new_n839), .B2(new_n835), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n683), .A2(KEYINPUT54), .A3(new_n832), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(KEYINPUT55), .A3(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n657), .A2(new_n838), .A3(new_n689), .A4(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n621), .B1(new_n827), .B2(new_n843), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n656), .A2(new_n825), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n845), .A2(new_n838), .A3(new_n689), .A4(new_n842), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n627), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n822), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n843), .A2(new_n827), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n627), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n842), .A2(new_n689), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n621), .A2(new_n845), .A3(new_n838), .A4(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(KEYINPUT111), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n848), .A2(new_n853), .A3(new_n544), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n657), .A2(new_n690), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n622), .A2(new_n628), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n403), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n857), .A2(KEYINPUT112), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n375), .B1(new_n857), .B2(KEYINPUT112), .ZN(new_n859));
  OR4_X1    g658(.A1(new_n345), .A2(new_n858), .A3(new_n859), .A4(new_n430), .ZN(new_n860));
  OAI21_X1  g659(.A(G113gat), .B1(new_n860), .B2(new_n658), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n345), .B1(new_n854), .B2(new_n856), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n281), .A3(new_n414), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n658), .A2(G113gat), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n864), .B(KEYINPUT113), .Z(new_n865));
  OAI21_X1  g664(.A(new_n861), .B1(new_n863), .B2(new_n865), .ZN(G1340gat));
  OAI21_X1  g665(.A(G120gat), .B1(new_n860), .B2(new_n768), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n768), .A2(G120gat), .ZN(new_n868));
  XOR2_X1   g667(.A(new_n868), .B(KEYINPUT114), .Z(new_n869));
  OAI21_X1  g668(.A(new_n867), .B1(new_n863), .B2(new_n869), .ZN(G1341gat));
  OAI21_X1  g669(.A(G127gat), .B1(new_n860), .B2(new_n544), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n543), .A2(new_n286), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n871), .B1(new_n863), .B2(new_n872), .ZN(G1342gat));
  OAI21_X1  g672(.A(G134gat), .B1(new_n860), .B2(new_n627), .ZN(new_n874));
  INV_X1    g673(.A(new_n862), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n281), .A2(new_n621), .A3(new_n284), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n875), .A2(new_n405), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT56), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n874), .A2(new_n878), .ZN(G1343gat));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n845), .A2(new_n690), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n827), .A2(KEYINPUT115), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n840), .A2(new_n883), .A3(new_n841), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n883), .B1(new_n840), .B2(new_n841), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT55), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n657), .A2(new_n689), .A3(new_n842), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n881), .B(new_n882), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n627), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n543), .B1(new_n889), .B2(new_n852), .ZN(new_n890));
  INV_X1    g689(.A(new_n856), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n403), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(KEYINPUT57), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n854), .A2(new_n856), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n404), .A2(KEYINPUT57), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n705), .A2(new_n345), .A3(new_n430), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n893), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(G141gat), .B1(new_n898), .B2(new_n658), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n875), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n706), .A2(new_n403), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n902), .B1(new_n862), .B2(KEYINPUT119), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n658), .A2(G141gat), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n901), .A2(new_n903), .A3(new_n281), .A4(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT58), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n899), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n898), .A2(KEYINPUT117), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n893), .A2(new_n896), .A3(new_n909), .A4(new_n897), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n908), .A2(new_n657), .A3(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT118), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n911), .A2(new_n912), .A3(G141gat), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n911), .B2(G141gat), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n862), .A2(KEYINPUT119), .ZN(new_n915));
  AOI211_X1 g714(.A(new_n900), .B(new_n345), .C1(new_n854), .C2(new_n856), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n915), .A2(new_n916), .A3(new_n902), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n917), .A2(KEYINPUT120), .A3(new_n281), .A4(new_n904), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n905), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n913), .A2(new_n914), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n907), .B1(new_n922), .B2(new_n906), .ZN(G1344gat));
  AND2_X1   g722(.A1(new_n908), .A2(new_n910), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n690), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT121), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT59), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n925), .A2(new_n926), .A3(new_n927), .A4(G148gat), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n917), .A2(new_n281), .ZN(new_n929));
  INV_X1    g728(.A(G148gat), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n690), .A2(new_n930), .ZN(new_n931));
  AOI211_X1 g730(.A(KEYINPUT59), .B(new_n930), .C1(new_n924), .C2(new_n690), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n894), .A2(KEYINPUT57), .A3(new_n403), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT57), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n892), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n897), .A2(new_n690), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n930), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT121), .B1(new_n939), .B2(new_n927), .ZN(new_n940));
  OAI221_X1 g739(.A(new_n928), .B1(new_n929), .B2(new_n931), .C1(new_n932), .C2(new_n940), .ZN(G1345gat));
  INV_X1    g740(.A(new_n924), .ZN(new_n942));
  OAI21_X1  g741(.A(G155gat), .B1(new_n942), .B2(new_n544), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n543), .A2(new_n301), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n929), .B2(new_n944), .ZN(G1346gat));
  OAI21_X1  g744(.A(G162gat), .B1(new_n942), .B2(new_n627), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n917), .A2(new_n302), .A3(new_n281), .A4(new_n621), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1347gat));
  AOI21_X1  g747(.A(new_n429), .B1(new_n854), .B2(new_n856), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n430), .A3(new_n414), .ZN(new_n950));
  XOR2_X1   g749(.A(new_n950), .B(KEYINPUT122), .Z(new_n951));
  AOI21_X1  g750(.A(G169gat), .B1(new_n951), .B2(new_n657), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n429), .A2(new_n281), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n858), .A2(new_n859), .A3(new_n954), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n658), .A2(new_n203), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(G1348gat));
  NAND3_X1  g756(.A1(new_n951), .A2(new_n204), .A3(new_n690), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n955), .A2(new_n690), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n959), .B2(new_n204), .ZN(G1349gat));
  NAND2_X1  g759(.A1(new_n543), .A2(new_n225), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n950), .A2(new_n961), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n955), .A2(new_n543), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n963), .B2(new_n215), .ZN(new_n964));
  AND2_X1   g763(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n964), .B(new_n965), .ZN(G1350gat));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n219), .A3(new_n621), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n955), .A2(new_n621), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n969), .B2(G190gat), .ZN(new_n970));
  AOI211_X1 g769(.A(KEYINPUT61), .B(new_n219), .C1(new_n955), .C2(new_n621), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(G1351gat));
  INV_X1    g771(.A(new_n902), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n949), .A2(new_n430), .A3(new_n973), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n974), .A2(G197gat), .A3(new_n658), .ZN(new_n975));
  XOR2_X1   g774(.A(new_n975), .B(KEYINPUT124), .Z(new_n976));
  NOR2_X1   g775(.A1(new_n705), .A2(new_n954), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n936), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g777(.A(G197gat), .B1(new_n978), .B2(new_n658), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n976), .A2(new_n979), .ZN(G1352gat));
  NOR3_X1   g779(.A1(new_n974), .A2(G204gat), .A3(new_n768), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g782(.A(G204gat), .B1(new_n978), .B2(new_n768), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n981), .A2(new_n982), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  XOR2_X1   g785(.A(new_n986), .B(KEYINPUT125), .Z(G1353gat));
  NOR3_X1   g786(.A1(new_n974), .A2(G211gat), .A3(new_n544), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n936), .A2(new_n977), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(new_n543), .ZN(new_n990));
  AOI21_X1  g789(.A(KEYINPUT63), .B1(new_n990), .B2(G211gat), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OR2_X1    g792(.A1(new_n991), .A2(new_n992), .ZN(new_n994));
  AND3_X1   g793(.A1(new_n990), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n993), .B1(new_n994), .B2(new_n995), .ZN(G1354gat));
  OR2_X1    g795(.A1(new_n989), .A2(KEYINPUT127), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n989), .A2(KEYINPUT127), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n997), .A2(new_n621), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(G218gat), .ZN(new_n1000));
  OR2_X1    g799(.A1(new_n627), .A2(G218gat), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n1000), .B1(new_n974), .B2(new_n1001), .ZN(G1355gat));
endmodule


