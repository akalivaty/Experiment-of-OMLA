//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n917, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n202));
  OAI21_X1  g001(.A(new_n202), .B1(G169gat), .B2(G176gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  AND2_X1   g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n206), .B1(KEYINPUT23), .B2(new_n207), .ZN(new_n208));
  AND2_X1   g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT24), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT66), .B(G183gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n211), .B1(G190gat), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n209), .A2(KEYINPUT25), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n211), .B1(G183gat), .B2(G190gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT25), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n214), .A2(KEYINPUT67), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n214), .A2(KEYINPUT67), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT27), .B(G183gat), .ZN(new_n221));
  INV_X1    g020(.A(G190gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(KEYINPUT28), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n212), .A2(KEYINPUT27), .ZN(new_n224));
  OR2_X1    g023(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n225));
  AOI21_X1  g024(.A(G190gat), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n223), .B1(new_n226), .B2(KEYINPUT28), .ZN(new_n227));
  INV_X1    g026(.A(new_n207), .ZN(new_n228));
  OAI22_X1  g027(.A1(new_n228), .A2(KEYINPUT68), .B1(KEYINPUT26), .B2(new_n206), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n228), .A2(KEYINPUT68), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n229), .B1(KEYINPUT26), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n227), .A2(new_n210), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n220), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G120gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G113gat), .ZN(new_n235));
  INV_X1    g034(.A(G113gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G120gat), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT1), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G127gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(KEYINPUT69), .A2(G127gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n240), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(G134gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n233), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G227gat), .A2(G233gat), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n246), .B(KEYINPUT64), .Z(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT32), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT33), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G15gat), .B(G43gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT70), .ZN(new_n253));
  XNOR2_X1  g052(.A(G71gat), .B(G99gat), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n253), .B(new_n254), .Z(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n249), .A2(new_n251), .A3(new_n256), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n248), .B(KEYINPUT32), .C1(new_n250), .C2(new_n255), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n242), .B(G134gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n233), .B(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n247), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT72), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n245), .A2(new_n247), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT34), .ZN(new_n268));
  AOI22_X1  g067(.A1(new_n265), .A2(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT72), .B1(new_n267), .B2(new_n261), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n259), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n257), .A2(new_n269), .A3(new_n270), .A4(new_n258), .ZN(new_n273));
  NOR2_X1   g072(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  XOR2_X1   g074(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n277), .B1(new_n272), .B2(new_n273), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT29), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n233), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G226gat), .A2(G233gat), .ZN(new_n282));
  XOR2_X1   g081(.A(new_n282), .B(KEYINPUT74), .Z(new_n283));
  AOI22_X1  g082(.A1(new_n281), .A2(new_n282), .B1(new_n233), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G197gat), .B(G204gat), .ZN(new_n285));
  INV_X1    g084(.A(G211gat), .ZN(new_n286));
  INV_X1    g085(.A(G218gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n285), .B1(KEYINPUT22), .B2(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(G211gat), .B(G218gat), .Z(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT75), .ZN(new_n293));
  INV_X1    g092(.A(new_n233), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n293), .B1(new_n294), .B2(new_n282), .ZN(new_n295));
  INV_X1    g094(.A(new_n283), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n233), .A2(KEYINPUT75), .A3(G226gat), .A4(G233gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n295), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT76), .ZN(new_n300));
  INV_X1    g099(.A(new_n291), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n300), .B1(new_n299), .B2(new_n301), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n292), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G8gat), .B(G36gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(G64gat), .B(G92gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n307), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n292), .B(new_n309), .C1(new_n302), .C2(new_n303), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(KEYINPUT30), .A3(new_n310), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n310), .A2(KEYINPUT30), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT77), .ZN(new_n313));
  INV_X1    g112(.A(G141gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n313), .B1(new_n314), .B2(G148gat), .ZN(new_n315));
  INV_X1    g114(.A(G148gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(KEYINPUT77), .A3(G141gat), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n315), .B(new_n317), .C1(G141gat), .C2(new_n316), .ZN(new_n318));
  OR2_X1    g117(.A1(new_n318), .A2(KEYINPUT78), .ZN(new_n319));
  NAND2_X1  g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320));
  OR3_X1    g119(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n318), .A2(KEYINPUT78), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  OR2_X1    g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(G141gat), .B(G148gat), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n320), .B(new_n324), .C1(new_n325), .C2(KEYINPUT2), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n262), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(KEYINPUT4), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(KEYINPUT4), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n329), .B1(KEYINPUT80), .B2(new_n330), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n330), .A2(KEYINPUT80), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT79), .B1(new_n327), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n323), .A2(new_n326), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT79), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT3), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n327), .A2(new_n335), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n336), .A2(new_n244), .A3(new_n339), .A4(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n333), .A2(new_n334), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT5), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n244), .A2(new_n337), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n334), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n343), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n330), .ZN(new_n349));
  OR2_X1    g148(.A1(new_n349), .A2(new_n329), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n346), .A2(KEYINPUT5), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n350), .A2(new_n341), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G1gat), .B(G29gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT0), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(KEYINPUT81), .ZN(new_n357));
  XOR2_X1   g156(.A(G57gat), .B(G85gat), .Z(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT6), .B1(new_n354), .B2(new_n360), .ZN(new_n361));
  NOR3_X1   g160(.A1(new_n354), .A2(KEYINPUT82), .A3(new_n360), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT82), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n352), .B1(new_n342), .B2(new_n347), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n363), .B1(new_n364), .B2(new_n359), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n361), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n354), .A2(KEYINPUT6), .A3(new_n360), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n311), .A2(new_n312), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n340), .A2(new_n280), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n335), .B1(new_n301), .B2(KEYINPUT29), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n369), .A2(new_n301), .B1(new_n337), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G228gat), .A2(G233gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G22gat), .ZN(new_n374));
  OR2_X1    g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n374), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G78gat), .B(G106gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT31), .B(G50gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT83), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n380), .B1(new_n376), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n375), .B(new_n376), .C1(new_n381), .C2(new_n380), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n279), .B1(new_n368), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT37), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n387), .B(new_n292), .C1(new_n302), .C2(new_n303), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n299), .A2(new_n291), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n387), .B1(new_n284), .B2(new_n301), .ZN(new_n390));
  AOI211_X1 g189(.A(KEYINPUT38), .B(new_n309), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n392), .A2(new_n310), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n359), .B(KEYINPUT84), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT6), .B1(new_n354), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n395), .B1(new_n362), .B2(new_n365), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n393), .A2(KEYINPUT86), .A3(new_n367), .A4(new_n396), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n396), .A2(new_n367), .A3(new_n392), .A4(new_n310), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT86), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n304), .A2(KEYINPUT37), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n388), .A2(new_n307), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT38), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n397), .A2(new_n400), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n385), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n334), .B1(new_n350), .B2(new_n341), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT39), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n394), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT39), .B1(new_n345), .B2(new_n346), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n410), .B(KEYINPUT85), .Z(new_n411));
  OAI211_X1 g210(.A(new_n408), .B(new_n409), .C1(new_n411), .C2(new_n406), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT40), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n412), .A2(new_n413), .ZN(new_n415));
  AOI211_X1 g214(.A(new_n414), .B(new_n415), .C1(new_n354), .C2(new_n394), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n310), .A2(KEYINPUT30), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n310), .A2(KEYINPUT30), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n417), .B1(new_n418), .B2(new_n308), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n405), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n386), .B1(new_n404), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT35), .ZN(new_n422));
  AND4_X1   g221(.A1(new_n422), .A2(new_n272), .A3(new_n273), .A4(new_n385), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n311), .A2(new_n312), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n396), .A2(new_n367), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n272), .A2(new_n273), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(new_n405), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n422), .B1(new_n368), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT87), .B1(new_n421), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n400), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n403), .B1(new_n398), .B2(new_n399), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n420), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n428), .A2(new_n276), .ZN(new_n436));
  INV_X1    g235(.A(new_n274), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n436), .B1(new_n428), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n368), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n438), .B1(new_n439), .B2(new_n405), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT87), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n368), .A2(new_n429), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT35), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n426), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G113gat), .B(G141gat), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT11), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(G169gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(G197gat), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n450), .A2(G197gat), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT12), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n453), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT12), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n456), .A3(new_n451), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT92), .ZN(new_n460));
  INV_X1    g259(.A(G1gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT16), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n374), .A2(G15gat), .ZN(new_n463));
  INV_X1    g262(.A(G15gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G22gat), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(G8gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G15gat), .B(G22gat), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n469), .A2(G1gat), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n460), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n463), .A2(new_n465), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n461), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n473), .A2(KEYINPUT92), .A3(new_n467), .A4(new_n466), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n466), .A2(KEYINPUT91), .B1(new_n472), .B2(new_n461), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT91), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n469), .A2(new_n477), .A3(new_n462), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n467), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(G43gat), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n481), .A2(G50gat), .ZN(new_n482));
  INV_X1    g281(.A(G50gat), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n483), .A2(G43gat), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT88), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(G43gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n481), .A2(G50gat), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT88), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n485), .A2(KEYINPUT15), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT14), .ZN(new_n491));
  INV_X1    g290(.A(G29gat), .ZN(new_n492));
  INV_X1    g291(.A(G36gat), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AND3_X1   g295(.A1(KEYINPUT90), .A2(G29gat), .A3(G36gat), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT90), .B1(G29gat), .B2(G36gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT15), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT89), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n502), .B1(new_n483), .B2(G43gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n486), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n487), .A2(new_n502), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n500), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT17), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n496), .B1(new_n492), .B2(new_n493), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n509), .A2(KEYINPUT15), .A3(new_n485), .A4(new_n489), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n508), .B1(new_n507), .B2(new_n510), .ZN(new_n512));
  OAI211_X1 g311(.A(KEYINPUT93), .B(new_n480), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G229gat), .A2(G233gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n466), .A2(KEYINPUT91), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n515), .A2(new_n478), .A3(new_n473), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G8gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(new_n471), .A3(new_n474), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n507), .A2(new_n510), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT17), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n507), .A2(new_n510), .A3(new_n508), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT93), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n523), .B1(new_n518), .B2(new_n519), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n513), .B(new_n514), .C1(new_n522), .C2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT18), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n514), .B(KEYINPUT13), .Z(new_n529));
  AND2_X1   g328(.A1(new_n507), .A2(new_n510), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n480), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n518), .A2(new_n519), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(new_n525), .B2(new_n526), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n459), .B1(new_n528), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n480), .B1(new_n511), .B2(new_n512), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(new_n531), .B2(new_n523), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n537), .A2(KEYINPUT18), .A3(new_n514), .A4(new_n513), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n527), .A2(new_n538), .A3(new_n458), .A4(new_n533), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n432), .A2(new_n446), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT94), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT94), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n432), .A2(new_n446), .A3(new_n543), .A4(new_n540), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G183gat), .B(G211gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT95), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G57gat), .B(G64gat), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G71gat), .ZN(new_n551));
  INV_X1    g350(.A(G78gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G71gat), .A2(G78gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n550), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n554), .B(new_n553), .C1(new_n549), .C2(new_n556), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n560), .A2(KEYINPUT21), .ZN(new_n561));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n561), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G127gat), .B(G155gat), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n561), .B(new_n562), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n565), .ZN(new_n569));
  XOR2_X1   g368(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n567), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n571), .B1(new_n567), .B2(new_n569), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n518), .B1(KEYINPUT21), .B2(new_n560), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n575), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n567), .A2(new_n569), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n570), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n577), .B1(new_n579), .B2(new_n572), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n548), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n575), .B1(new_n573), .B2(new_n574), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(new_n577), .A3(new_n572), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n582), .A2(new_n583), .A3(new_n547), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT100), .ZN(new_n586));
  XOR2_X1   g385(.A(G99gat), .B(G106gat), .Z(new_n587));
  NAND2_X1  g386(.A1(G99gat), .A2(G106gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT8), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT99), .ZN(new_n590));
  OR2_X1    g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n590), .B1(new_n589), .B2(new_n591), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(KEYINPUT97), .A2(KEYINPUT98), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n595), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT7), .ZN(new_n597));
  NAND2_X1  g396(.A1(G85gat), .A2(G92gat), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n597), .B1(new_n598), .B2(KEYINPUT98), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(KEYINPUT97), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n596), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n587), .B1(new_n594), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT8), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n603), .B1(G99gat), .B2(G106gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(G85gat), .A2(G92gat), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT99), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n589), .A2(new_n591), .A3(new_n590), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n587), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n596), .A2(new_n599), .A3(new_n600), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n602), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n612), .B1(new_n511), .B2(new_n512), .ZN(new_n613));
  AND3_X1   g412(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n609), .B1(new_n608), .B2(new_n610), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n614), .B1(new_n617), .B2(new_n519), .ZN(new_n618));
  XNOR2_X1  g417(.A(G190gat), .B(G218gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n613), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n620), .B1(new_n613), .B2(new_n618), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT96), .ZN(new_n624));
  XOR2_X1   g423(.A(G134gat), .B(G162gat), .Z(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  OR4_X1    g425(.A1(new_n586), .A2(new_n621), .A3(new_n622), .A4(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n586), .B1(new_n621), .B2(new_n622), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n618), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n619), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n613), .A2(new_n618), .A3(new_n620), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n631), .A3(KEYINPUT100), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n628), .A2(new_n632), .A3(new_n626), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n585), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n558), .A2(new_n559), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n636), .B1(new_n615), .B2(new_n616), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT10), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n602), .A2(new_n560), .A3(new_n611), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n617), .A2(KEYINPUT10), .A3(new_n560), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(G230gat), .A2(G233gat), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n643), .B1(new_n637), .B2(new_n639), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n644), .A2(new_n646), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n643), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n640), .B2(new_n641), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n649), .B1(new_n653), .B2(new_n645), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n545), .A2(new_n635), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n366), .A2(new_n367), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(G1gat), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n657), .A2(new_n461), .A3(new_n659), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(G1324gat));
  NAND2_X1  g462(.A1(new_n467), .A2(KEYINPUT42), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n664), .B1(new_n657), .B2(new_n419), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n657), .A2(new_n419), .ZN(new_n666));
  NOR2_X1   g465(.A1(KEYINPUT102), .A2(KEYINPUT42), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT101), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT16), .B(G8gat), .Z(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n665), .B1(new_n666), .B2(new_n670), .ZN(G1325gat));
  INV_X1    g470(.A(new_n428), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n657), .A2(new_n464), .A3(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n657), .A2(new_n438), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n673), .B1(new_n674), .B2(new_n464), .ZN(G1326gat));
  XNOR2_X1  g474(.A(KEYINPUT43), .B(G22gat), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n657), .A2(new_n405), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n676), .B1(new_n657), .B2(new_n405), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(G1327gat));
  INV_X1    g478(.A(KEYINPUT45), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n585), .A2(new_n634), .A3(new_n656), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT103), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n658), .A2(G29gat), .ZN(new_n684));
  AND4_X1   g483(.A1(new_n681), .A2(new_n545), .A3(new_n683), .A4(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n683), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n686), .B1(new_n542), .B2(new_n544), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n681), .B1(new_n687), .B2(new_n684), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n680), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n545), .A2(new_n683), .A3(new_n684), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT104), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n687), .A2(new_n681), .A3(new_n684), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(KEYINPUT45), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT105), .B1(new_n427), .B2(new_n430), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n444), .A2(new_n695), .A3(new_n426), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n441), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n634), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n432), .A2(new_n446), .A3(KEYINPUT44), .A4(new_n634), .ZN(new_n701));
  INV_X1    g500(.A(new_n585), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n535), .A2(new_n539), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n702), .A2(new_n703), .A3(new_n655), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n700), .A2(new_n659), .A3(new_n701), .A4(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n492), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(new_n706), .B2(new_n705), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n689), .A2(new_n693), .A3(new_n708), .ZN(G1328gat));
  NAND2_X1  g508(.A1(new_n419), .A2(new_n493), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n687), .A2(KEYINPUT46), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT46), .B1(new_n687), .B2(new_n711), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n700), .A2(new_n701), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n714), .A2(new_n419), .A3(new_n704), .ZN(new_n715));
  OAI22_X1  g514(.A1(new_n712), .A2(new_n713), .B1(new_n715), .B2(new_n493), .ZN(G1329gat));
  INV_X1    g515(.A(KEYINPUT47), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n279), .A2(new_n481), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n714), .A2(new_n704), .A3(new_n718), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n687), .A2(new_n672), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n717), .B(new_n719), .C1(new_n720), .C2(G43gat), .ZN(new_n721));
  INV_X1    g520(.A(new_n719), .ZN(new_n722));
  AOI21_X1  g521(.A(G43gat), .B1(new_n687), .B2(new_n672), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT47), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n724), .ZN(G1330gat));
  NAND3_X1  g524(.A1(new_n545), .A2(new_n405), .A3(new_n683), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n483), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n385), .A2(new_n483), .ZN(new_n728));
  AND4_X1   g527(.A1(new_n700), .A2(new_n701), .A3(new_n704), .A4(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT48), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT48), .ZN(new_n732));
  AOI211_X1 g531(.A(new_n732), .B(new_n729), .C1(new_n726), .C2(new_n483), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n731), .A2(new_n733), .ZN(G1331gat));
  NAND2_X1  g533(.A1(new_n635), .A2(new_n703), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n656), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT107), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n697), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n659), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n419), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  AND2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n745), .B1(new_n743), .B2(new_n742), .ZN(G1333gat));
  OAI21_X1  g545(.A(new_n551), .B1(new_n738), .B2(new_n428), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n438), .A2(G71gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n738), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g549(.A1(new_n738), .A2(new_n385), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(new_n552), .ZN(G1335gat));
  NOR3_X1   g551(.A1(new_n702), .A2(new_n540), .A3(new_n656), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n714), .A2(new_n659), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT108), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G85gat), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n754), .A2(KEYINPUT108), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n697), .A2(new_n703), .A3(new_n585), .A4(new_n634), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(KEYINPUT109), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n758), .B2(new_n759), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n761), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(G85gat), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n659), .A2(new_n765), .A3(new_n655), .ZN(new_n766));
  OAI22_X1  g565(.A1(new_n756), .A2(new_n757), .B1(new_n764), .B2(new_n766), .ZN(G1336gat));
  OR3_X1    g566(.A1(new_n424), .A2(G92gat), .A3(new_n656), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n700), .A2(new_n419), .A3(new_n701), .A4(new_n753), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G92gat), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n759), .A2(KEYINPUT111), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n758), .B(new_n774), .Z(new_n775));
  XOR2_X1   g574(.A(new_n768), .B(KEYINPUT110), .Z(new_n776));
  AOI22_X1  g575(.A1(new_n775), .A2(new_n776), .B1(new_n770), .B2(G92gat), .ZN(new_n777));
  OAI22_X1  g576(.A1(new_n769), .A2(new_n773), .B1(new_n777), .B2(new_n772), .ZN(G1337gat));
  NAND3_X1  g577(.A1(new_n714), .A2(new_n438), .A3(new_n753), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G99gat), .ZN(new_n780));
  OR3_X1    g579(.A1(new_n428), .A2(G99gat), .A3(new_n656), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n764), .B2(new_n781), .ZN(G1338gat));
  NOR3_X1   g581(.A1(new_n385), .A2(G106gat), .A3(new_n656), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n764), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n700), .A2(new_n405), .A3(new_n701), .A4(new_n753), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G106gat), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n775), .A2(new_n783), .B1(new_n786), .B2(G106gat), .ZN(new_n790));
  OAI22_X1  g589(.A1(new_n785), .A2(new_n789), .B1(new_n790), .B2(new_n788), .ZN(G1339gat));
  NAND3_X1  g590(.A1(new_n635), .A2(new_n703), .A3(new_n656), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n640), .A2(new_n641), .A3(new_n652), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n644), .A2(KEYINPUT54), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n650), .B1(new_n653), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n794), .A2(KEYINPUT55), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n651), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT55), .B1(new_n794), .B2(new_n796), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n514), .B1(new_n537), .B2(new_n513), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n531), .A2(new_n532), .A3(new_n529), .ZN(new_n802));
  OAI22_X1  g601(.A1(new_n801), .A2(new_n802), .B1(new_n452), .B2(new_n453), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n800), .A2(new_n634), .A3(new_n539), .A4(new_n803), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n539), .A2(new_n803), .A3(new_n655), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n805), .B1(new_n800), .B2(new_n540), .ZN(new_n806));
  OAI211_X1 g605(.A(KEYINPUT112), .B(new_n804), .C1(new_n806), .C2(new_n634), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n585), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n539), .A2(new_n803), .A3(new_n655), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n796), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(new_n651), .A3(new_n797), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n809), .B1(new_n703), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n634), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT112), .B1(new_n816), .B2(new_n804), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n792), .B1(new_n808), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT113), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n820), .B(new_n792), .C1(new_n808), .C2(new_n817), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n659), .ZN(new_n823));
  NOR4_X1   g622(.A1(new_n823), .A2(new_n419), .A3(new_n428), .A4(new_n405), .ZN(new_n824));
  AOI21_X1  g623(.A(G113gat), .B1(new_n824), .B2(new_n540), .ZN(new_n825));
  XOR2_X1   g624(.A(new_n824), .B(KEYINPUT114), .Z(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n703), .A2(new_n236), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(G1340gat));
  AOI21_X1  g628(.A(G120gat), .B1(new_n824), .B2(new_n655), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n656), .A2(new_n234), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n830), .B1(new_n827), .B2(new_n831), .ZN(G1341gat));
  OAI21_X1  g631(.A(G127gat), .B1(new_n826), .B2(new_n585), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n824), .A2(new_n239), .A3(new_n702), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(G1342gat));
  OAI21_X1  g634(.A(G134gat), .B1(new_n826), .B2(new_n815), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n823), .A2(new_n428), .A3(new_n405), .ZN(new_n837));
  XOR2_X1   g636(.A(KEYINPUT69), .B(G134gat), .Z(new_n838));
  NAND4_X1  g637(.A1(new_n837), .A2(new_n424), .A3(new_n634), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT56), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT115), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n836), .B(new_n841), .C1(KEYINPUT56), .C2(new_n839), .ZN(G1343gat));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n438), .A2(new_n658), .A3(new_n419), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n819), .A2(new_n405), .A3(new_n821), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n810), .B(KEYINPUT117), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(KEYINPUT55), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n540), .A2(new_n651), .A3(new_n797), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n809), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n815), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n702), .B1(new_n853), .B2(new_n804), .ZN(new_n854));
  INV_X1    g653(.A(new_n792), .ZN(new_n855));
  OAI211_X1 g654(.A(KEYINPUT57), .B(new_n405), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n848), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n846), .B1(new_n845), .B2(new_n847), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n844), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n843), .B1(new_n859), .B2(new_n703), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n847), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT116), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n848), .A3(new_n856), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n863), .A2(KEYINPUT120), .A3(new_n540), .A4(new_n844), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n860), .A2(G141gat), .A3(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n823), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n822), .A2(KEYINPUT119), .A3(new_n659), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n438), .A2(new_n385), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n867), .A2(new_n424), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n703), .A2(G141gat), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT58), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n865), .A2(new_n873), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n870), .A2(G141gat), .A3(new_n703), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n859), .A2(KEYINPUT118), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n863), .A2(new_n877), .A3(new_n844), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n540), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n875), .B1(new_n879), .B2(G141gat), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT58), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n874), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g683(.A(KEYINPUT121), .B(new_n874), .C1(new_n880), .C2(new_n881), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1344gat));
  NAND4_X1  g685(.A1(new_n819), .A2(KEYINPUT57), .A3(new_n405), .A4(new_n821), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n887), .B(new_n888), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n792), .A2(KEYINPUT123), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n792), .A2(KEYINPUT123), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n854), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n847), .B1(new_n892), .B2(new_n385), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(new_n656), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n895), .A2(new_n844), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT59), .B1(new_n896), .B2(new_n316), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n316), .A2(KEYINPUT59), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n876), .A2(new_n878), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(new_n656), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n871), .A2(new_n316), .A3(new_n655), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1345gat));
  INV_X1    g702(.A(G155gat), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n899), .A2(new_n904), .A3(new_n585), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n870), .A2(new_n585), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n906), .A2(KEYINPUT124), .ZN(new_n907));
  AOI21_X1  g706(.A(G155gat), .B1(new_n906), .B2(KEYINPUT124), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(G1346gat));
  OAI21_X1  g708(.A(G162gat), .B1(new_n899), .B2(new_n815), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n419), .A2(G162gat), .A3(new_n815), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n867), .A2(new_n868), .A3(new_n869), .A4(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1347gat));
  AND4_X1   g712(.A1(new_n658), .A2(new_n822), .A3(new_n419), .A4(new_n429), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n540), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n655), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g717(.A1(new_n914), .A2(new_n702), .ZN(new_n919));
  MUX2_X1   g718(.A(new_n221), .B(new_n212), .S(new_n919), .Z(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g720(.A1(new_n914), .A2(new_n634), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(G190gat), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT61), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n924), .B1(G190gat), .B2(new_n922), .ZN(G1351gat));
  NOR3_X1   g724(.A1(new_n438), .A2(new_n659), .A3(new_n424), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n927), .A2(new_n845), .ZN(new_n928));
  AOI21_X1  g727(.A(G197gat), .B1(new_n928), .B2(new_n540), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n927), .B1(new_n889), .B2(new_n893), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n540), .A2(G197gat), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(G1352gat));
  XNOR2_X1  g731(.A(KEYINPUT125), .B(G204gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n928), .A2(new_n655), .A3(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT126), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n894), .A2(new_n656), .A3(new_n927), .ZN(new_n939));
  OAI221_X1 g738(.A(new_n938), .B1(new_n936), .B2(new_n935), .C1(new_n939), .C2(new_n933), .ZN(G1353gat));
  NAND3_X1  g739(.A1(new_n928), .A2(new_n286), .A3(new_n702), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n286), .B1(new_n930), .B2(new_n702), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n942), .A2(KEYINPUT63), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(KEYINPUT63), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g746(.A(KEYINPUT127), .B(new_n941), .C1(new_n943), .C2(new_n944), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1354gat));
  NAND3_X1  g748(.A1(new_n928), .A2(new_n287), .A3(new_n634), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n930), .A2(new_n634), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(new_n951), .B2(new_n287), .ZN(G1355gat));
endmodule


