//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n968, new_n969;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n202));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203));
  OR3_X1    g002(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n204), .B(new_n205), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G183gat), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(new_n209), .B2(KEYINPUT27), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT27), .B(G183gat), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n210), .B(new_n214), .C1(new_n215), .C2(new_n213), .ZN(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n215), .A2(KEYINPUT28), .A3(new_n210), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n208), .B(new_n212), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(new_n206), .A3(new_n207), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n222), .A2(new_n223), .B1(G169gat), .B2(G176gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(new_n209), .B2(new_n210), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(G183gat), .B2(G190gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n224), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT25), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n229), .B(new_n225), .C1(G183gat), .C2(G190gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(KEYINPUT25), .A3(new_n224), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT65), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n234), .A2(new_n237), .A3(new_n224), .A4(KEYINPUT25), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n233), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n203), .B1(new_n220), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n239), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n240), .B1(new_n244), .B2(new_n203), .ZN(new_n245));
  INV_X1    g044(.A(G218gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT22), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT73), .B(G218gat), .ZN(new_n248));
  INV_X1    g047(.A(G211gat), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G197gat), .B(G204gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n246), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n250), .A2(new_n251), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G211gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n257), .A2(G218gat), .A3(new_n252), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n202), .B1(new_n245), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n203), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n241), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n242), .B1(new_n220), .B2(new_n239), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n262), .B1(new_n263), .B2(new_n261), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n264), .A2(KEYINPUT75), .A3(new_n258), .A4(new_n255), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT29), .B1(new_n220), .B2(new_n239), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n262), .B(new_n259), .C1(new_n266), .C2(new_n261), .ZN(new_n267));
  XNOR2_X1  g066(.A(G8gat), .B(G36gat), .ZN(new_n268));
  INV_X1    g067(.A(G64gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G92gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n260), .A2(new_n265), .A3(new_n267), .A4(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT30), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n265), .A3(new_n267), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n272), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT76), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n274), .B(new_n279), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n276), .B(new_n278), .C1(new_n280), .C2(KEYINPUT30), .ZN(new_n281));
  XOR2_X1   g080(.A(G141gat), .B(G148gat), .Z(new_n282));
  XOR2_X1   g081(.A(KEYINPUT78), .B(KEYINPUT2), .Z(new_n283));
  AOI22_X1  g082(.A1(new_n282), .A2(new_n283), .B1(G155gat), .B2(G162gat), .ZN(new_n284));
  OR2_X1    g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n285), .B(KEYINPUT77), .ZN(new_n286));
  NAND2_X1  g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(new_n285), .B2(KEYINPUT2), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n284), .A2(new_n286), .B1(new_n288), .B2(new_n282), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT3), .ZN(new_n291));
  XOR2_X1   g090(.A(KEYINPUT68), .B(G134gat), .Z(new_n292));
  INV_X1    g091(.A(G127gat), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(G127gat), .A2(G134gat), .ZN(new_n295));
  XOR2_X1   g094(.A(G113gat), .B(G120gat), .Z(new_n296));
  INV_X1    g095(.A(KEYINPUT1), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G127gat), .B(G134gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n296), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT69), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n301), .A2(new_n302), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n299), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT79), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT3), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n289), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n307), .B1(new_n289), .B2(new_n308), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n291), .B(new_n306), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT4), .B1(new_n306), .B2(new_n290), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n301), .A2(new_n302), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(new_n303), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT4), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n315), .A2(new_n316), .A3(new_n289), .A4(new_n299), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G225gat), .A2(G233gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n320), .B(KEYINPUT80), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  OR2_X1    g121(.A1(new_n322), .A2(KEYINPUT39), .ZN(new_n323));
  XNOR2_X1  g122(.A(G1gat), .B(G29gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(KEYINPUT0), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n325), .B(G57gat), .ZN(new_n326));
  INV_X1    g125(.A(G85gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n314), .A2(new_n303), .B1(new_n294), .B2(new_n298), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n289), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n306), .A2(new_n290), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT39), .B1(new_n332), .B2(new_n321), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(KEYINPUT86), .ZN(new_n334));
  INV_X1    g133(.A(new_n322), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n323), .B(new_n328), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(KEYINPUT40), .ZN(new_n337));
  INV_X1    g136(.A(new_n319), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n321), .A2(KEYINPUT5), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT82), .B1(new_n332), .B2(new_n321), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT82), .ZN(new_n342));
  INV_X1    g141(.A(new_n321), .ZN(new_n343));
  AOI211_X1 g142(.A(new_n342), .B(new_n343), .C1(new_n330), .C2(new_n331), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT5), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT81), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n317), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n329), .A2(KEYINPUT81), .A3(new_n316), .A4(new_n289), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n348), .A3(new_n313), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n349), .A2(new_n312), .A3(new_n343), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n340), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT87), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n328), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n349), .A2(new_n312), .A3(new_n343), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n355), .B(KEYINPUT5), .C1(new_n341), .C2(new_n344), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n356), .A2(KEYINPUT87), .A3(new_n340), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n353), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n281), .A2(new_n337), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G22gat), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT29), .ZN(new_n361));
  NOR3_X1   g160(.A1(new_n253), .A2(new_n246), .A3(new_n254), .ZN(new_n362));
  AOI21_X1  g161(.A(G218gat), .B1(new_n257), .B2(new_n252), .ZN(new_n363));
  OAI211_X1 g162(.A(KEYINPUT83), .B(new_n361), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n308), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT83), .B1(new_n259), .B2(new_n361), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n290), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n289), .A2(new_n308), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT79), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n242), .B1(new_n369), .B2(new_n309), .ZN(new_n370));
  OR2_X1    g169(.A1(new_n370), .A2(new_n259), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n367), .A2(G228gat), .A3(new_n371), .A4(G233gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(G228gat), .A2(G233gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n370), .A2(new_n259), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n259), .A2(new_n243), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n289), .B1(new_n375), .B2(new_n308), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n373), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n360), .B1(new_n372), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n372), .A2(new_n360), .A3(new_n377), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(KEYINPUT84), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n380), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT84), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XOR2_X1   g183(.A(G78gat), .B(G106gat), .Z(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(KEYINPUT31), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n386), .B(G50gat), .Z(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n381), .A2(new_n384), .A3(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n382), .A2(new_n378), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT85), .B1(new_n390), .B2(new_n387), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n392));
  NOR4_X1   g191(.A1(new_n382), .A2(new_n378), .A3(new_n392), .A4(new_n388), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n389), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT6), .ZN(new_n395));
  AOI211_X1 g194(.A(new_n395), .B(new_n328), .C1(new_n356), .C2(new_n340), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n356), .A2(new_n328), .A3(new_n340), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n397), .A2(new_n395), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n396), .B1(new_n358), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n274), .B(KEYINPUT76), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n277), .A2(KEYINPUT37), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n272), .B1(new_n277), .B2(KEYINPUT37), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT38), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n264), .A2(new_n259), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n262), .B1(new_n266), .B2(new_n261), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n404), .B(KEYINPUT37), .C1(new_n405), .C2(new_n259), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT38), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n399), .A2(new_n400), .A3(new_n403), .A4(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n359), .A2(new_n394), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT88), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n241), .B(new_n306), .ZN(new_n413));
  NAND2_X1  g212(.A1(G227gat), .A2(G233gat), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT32), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT33), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G15gat), .B(G43gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT70), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(G71gat), .ZN(new_n422));
  INV_X1    g221(.A(G99gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n417), .A2(new_n419), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(KEYINPUT33), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n416), .A2(KEYINPUT32), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n425), .A2(KEYINPUT71), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT71), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n417), .A2(new_n419), .A3(new_n429), .A4(new_n424), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  OAI22_X1  g230(.A1(new_n413), .A2(new_n415), .B1(KEYINPUT72), .B2(KEYINPUT34), .ZN(new_n432));
  NAND2_X1  g231(.A1(KEYINPUT72), .A2(KEYINPUT34), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n428), .A2(new_n430), .A3(new_n434), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(KEYINPUT36), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n437), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT36), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n390), .A2(KEYINPUT85), .A3(new_n387), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n379), .A2(new_n380), .A3(new_n387), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n392), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n378), .A2(new_n383), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n387), .B1(new_n445), .B2(new_n380), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n442), .A2(new_n444), .B1(new_n446), .B2(new_n384), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n400), .A2(new_n275), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n351), .A2(new_n354), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n449), .A2(new_n395), .A3(new_n397), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n351), .A2(KEYINPUT6), .A3(new_n354), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n448), .A2(new_n452), .A3(new_n276), .A4(new_n278), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n438), .A2(new_n441), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT88), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n359), .A2(new_n394), .A3(new_n410), .A4(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n412), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n444), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n439), .B1(new_n458), .B2(new_n389), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n281), .A2(new_n399), .A3(KEYINPUT35), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n447), .A2(new_n453), .A3(new_n439), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT35), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n457), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G15gat), .B(G22gat), .ZN(new_n466));
  INV_X1    g265(.A(G1gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT16), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n466), .A2(G1gat), .ZN(new_n471));
  OAI21_X1  g270(.A(G8gat), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(G8gat), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n469), .B(new_n473), .C1(G1gat), .C2(new_n466), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT17), .ZN(new_n476));
  XNOR2_X1  g275(.A(G43gat), .B(G50gat), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT15), .ZN(new_n479));
  NOR2_X1   g278(.A1(G29gat), .A2(G36gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(G29gat), .A2(G36gat), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n480), .B1(KEYINPUT14), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(G29gat), .ZN(new_n483));
  INV_X1    g282(.A(G36gat), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT14), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n479), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n481), .A2(KEYINPUT14), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n483), .A2(new_n484), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n480), .A2(KEYINPUT14), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(KEYINPUT15), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n478), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n491), .A2(new_n478), .ZN(new_n493));
  OAI211_X1 g292(.A(KEYINPUT90), .B(new_n476), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NOR3_X1   g293(.A1(new_n482), .A2(new_n479), .A3(new_n485), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT15), .B1(new_n489), .B2(new_n490), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n477), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n491), .A2(new_n478), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n476), .A2(KEYINPUT90), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n476), .A2(KEYINPUT90), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n475), .B1(new_n494), .B2(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n472), .A2(new_n474), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n497), .A2(new_n498), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(G229gat), .A2(G233gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT91), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n502), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT18), .B1(new_n509), .B2(KEYINPUT92), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n501), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(new_n503), .ZN(new_n512));
  INV_X1    g311(.A(new_n504), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n475), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n512), .A2(new_n514), .A3(new_n507), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT92), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT18), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n507), .B(KEYINPUT13), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n504), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n520), .B1(new_n522), .B2(new_n505), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n510), .A2(new_n518), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n525));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  XOR2_X1   g326(.A(G169gat), .B(G197gat), .Z(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT12), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n510), .A2(new_n518), .A3(new_n530), .A4(new_n523), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(KEYINPUT93), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT93), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n524), .A2(new_n535), .A3(new_n531), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G71gat), .A2(G78gat), .ZN(new_n538));
  INV_X1    g337(.A(G71gat), .ZN(new_n539));
  INV_X1    g338(.A(G78gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G57gat), .A2(G64gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT9), .ZN(new_n543));
  NOR2_X1   g342(.A1(G57gat), .A2(G64gat), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n538), .B(new_n541), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT94), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT9), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n538), .B1(new_n541), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(KEYINPUT95), .A2(G57gat), .A3(G64gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT95), .ZN(new_n551));
  INV_X1    g350(.A(G57gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n269), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n549), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n269), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n555), .A2(KEYINPUT9), .A3(new_n542), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n556), .A2(KEYINPUT94), .A3(new_n538), .A4(new_n541), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n547), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G85gat), .A2(G92gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT7), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT7), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(G85gat), .A3(G92gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G99gat), .A2(G106gat), .ZN(new_n564));
  AOI22_X1  g363(.A1(KEYINPUT8), .A2(new_n564), .B1(new_n327), .B2(new_n271), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n564), .ZN(new_n567));
  NOR2_X1   g366(.A1(G99gat), .A2(G106gat), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n567), .A2(new_n568), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n563), .A2(new_n570), .A3(new_n565), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n558), .A2(new_n572), .A3(KEYINPUT10), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n563), .A2(new_n570), .A3(new_n565), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n570), .B1(new_n563), .B2(new_n565), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n566), .A2(KEYINPUT100), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n558), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n577), .A2(new_n547), .A3(new_n554), .A4(new_n557), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n572), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT10), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT101), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT101), .ZN(new_n584));
  AOI211_X1 g383(.A(new_n584), .B(KEYINPUT10), .C1(new_n578), .C2(new_n580), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n573), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G230gat), .A2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT102), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n578), .A2(new_n588), .A3(new_n580), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G120gat), .B(G148gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(new_n207), .ZN(new_n594));
  INV_X1    g393(.A(G204gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n596), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n590), .A2(new_n591), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n537), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n547), .A2(new_n554), .A3(new_n557), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT21), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(G127gat), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n503), .B1(new_n603), .B2(new_n602), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n608));
  XNOR2_X1  g407(.A(G183gat), .B(G211gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n607), .B(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(KEYINPUT96), .B(G155gat), .Z(new_n612));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n611), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n511), .A2(new_n576), .ZN(new_n617));
  NAND2_X1  g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n618), .B(KEYINPUT97), .Z(new_n619));
  INV_X1    g418(.A(KEYINPUT41), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n504), .A2(new_n576), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n617), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(G190gat), .B(G218gat), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT98), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n619), .A2(new_n620), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G134gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G162gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(KEYINPUT99), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n625), .A2(new_n627), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n572), .B1(new_n494), .B2(new_n501), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n635), .A2(new_n621), .A3(new_n623), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n626), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT98), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n639), .B1(new_n636), .B2(new_n626), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT99), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(new_n641), .A3(new_n631), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n633), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n638), .B1(new_n633), .B2(new_n642), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n616), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n465), .A2(new_n601), .A3(new_n646), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n647), .A2(KEYINPUT103), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(KEYINPUT103), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n452), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT104), .B(G1gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1324gat));
  NAND2_X1  g453(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n655));
  INV_X1    g454(.A(new_n649), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n647), .A2(KEYINPUT103), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n281), .B(new_n655), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n659));
  INV_X1    g458(.A(new_n281), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n660), .B1(new_n648), .B2(new_n649), .ZN(new_n661));
  OAI22_X1  g460(.A1(new_n658), .A2(new_n659), .B1(new_n661), .B2(new_n473), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT42), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT42), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n664), .B1(new_n658), .B2(new_n659), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(G1325gat));
  NAND2_X1  g465(.A1(new_n441), .A2(new_n438), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n667), .B1(new_n648), .B2(new_n649), .ZN(new_n668));
  INV_X1    g467(.A(G15gat), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI211_X1 g469(.A(G15gat), .B(new_n439), .C1(new_n648), .C2(new_n649), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT105), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n439), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n650), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n674), .B(new_n675), .C1(new_n669), .C2(new_n668), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n672), .A2(new_n676), .ZN(G1326gat));
  NAND2_X1  g476(.A1(new_n650), .A2(new_n447), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT43), .B(G22gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  NAND2_X1  g479(.A1(new_n465), .A2(new_n645), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n601), .A2(new_n616), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n683), .A2(new_n483), .A3(new_n651), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT45), .ZN(new_n685));
  INV_X1    g484(.A(new_n645), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(KEYINPUT44), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n457), .A2(new_n688), .A3(new_n464), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n457), .B2(new_n464), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n687), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n681), .A2(KEYINPUT44), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n682), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G29gat), .B1(new_n694), .B2(new_n452), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n685), .A2(new_n695), .ZN(G1328gat));
  NAND3_X1  g495(.A1(new_n683), .A2(new_n484), .A3(new_n281), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT46), .Z(new_n698));
  OAI21_X1  g497(.A(G36gat), .B1(new_n694), .B2(new_n660), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(G1329gat));
  INV_X1    g499(.A(G43gat), .ZN(new_n701));
  INV_X1    g500(.A(new_n667), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n693), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT47), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n686), .B1(new_n457), .B2(new_n464), .ZN(new_n705));
  INV_X1    g504(.A(new_n682), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n705), .A2(new_n701), .A3(new_n673), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT107), .ZN(new_n708));
  OR3_X1    g507(.A1(new_n703), .A2(new_n704), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n704), .B1(new_n703), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(G1330gat));
  INV_X1    g510(.A(new_n687), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n465), .A2(KEYINPUT106), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n457), .A2(new_n688), .A3(new_n464), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n705), .A2(new_n716), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n447), .B(new_n706), .C1(new_n715), .C2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n718), .A2(new_n719), .A3(G50gat), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT48), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n394), .A2(G50gat), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT108), .B1(new_n722), .B2(KEYINPUT109), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n683), .B(new_n723), .C1(KEYINPUT109), .C2(new_n722), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n720), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n721), .B1(new_n720), .B2(new_n724), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(G1331gat));
  INV_X1    g526(.A(new_n600), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(new_n713), .B2(new_n714), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n534), .A2(new_n536), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n730), .A2(new_n616), .A3(new_n645), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n452), .B(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(KEYINPUT111), .B(G57gat), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1332gat));
  XOR2_X1   g537(.A(new_n281), .B(KEYINPUT112), .Z(new_n739));
  NOR2_X1   g538(.A1(new_n732), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  AND2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(new_n740), .B2(new_n741), .ZN(G1333gat));
  OAI21_X1  g543(.A(G71gat), .B1(new_n732), .B2(new_n667), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n729), .A2(new_n539), .A3(new_n673), .A4(new_n731), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1334gat));
  NOR2_X1   g548(.A1(new_n732), .A2(new_n394), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(new_n540), .ZN(G1335gat));
  INV_X1    g550(.A(new_n616), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n730), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n465), .A2(new_n645), .A3(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n705), .A2(KEYINPUT51), .A3(new_n753), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n758), .A2(new_n327), .A3(new_n651), .A4(new_n600), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n753), .A2(new_n600), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n760), .B1(new_n691), .B2(new_n692), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n761), .A2(new_n651), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n759), .B1(new_n762), .B2(new_n327), .ZN(G1336gat));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n281), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n739), .B1(new_n756), .B2(new_n757), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n728), .A2(G92gat), .ZN(new_n766));
  AOI22_X1  g565(.A1(new_n764), .A2(G92gat), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  INV_X1    g567(.A(new_n739), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n271), .B1(new_n761), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n765), .A2(new_n766), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n768), .ZN(new_n772));
  OAI22_X1  g571(.A1(new_n767), .A2(new_n768), .B1(new_n770), .B2(new_n772), .ZN(G1337gat));
  NAND4_X1  g572(.A1(new_n758), .A2(new_n423), .A3(new_n600), .A4(new_n673), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n761), .A2(new_n702), .ZN(new_n775));
  OAI211_X1 g574(.A(KEYINPUT113), .B(new_n774), .C1(new_n775), .C2(new_n423), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777));
  INV_X1    g576(.A(new_n774), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n423), .B1(new_n761), .B2(new_n702), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n776), .A2(new_n780), .ZN(G1338gat));
  INV_X1    g580(.A(new_n760), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n447), .B(new_n782), .C1(new_n715), .C2(new_n717), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G106gat), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(G106gat), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n758), .A2(new_n787), .A3(new_n600), .A4(new_n447), .ZN(new_n788));
  AOI211_X1 g587(.A(new_n394), .B(new_n760), .C1(new_n691), .C2(new_n692), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n789), .B2(new_n787), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n786), .A2(new_n790), .A3(KEYINPUT53), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n784), .B(new_n788), .C1(new_n785), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(G1339gat));
  AND2_X1   g593(.A1(new_n731), .A2(new_n728), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n508), .B1(new_n502), .B2(new_n505), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n514), .A2(new_n521), .A3(new_n519), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n529), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT115), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n798), .A2(new_n801), .A3(new_n529), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n533), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n600), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n588), .B(new_n573), .C1(new_n583), .C2(new_n585), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT54), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n576), .B1(new_n558), .B2(new_n577), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n579), .A2(new_n572), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n582), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n584), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n581), .A2(KEYINPUT101), .A3(new_n582), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n588), .B1(new_n813), .B2(new_n573), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n807), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n586), .A2(new_n816), .A3(new_n589), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n596), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n805), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n590), .A2(KEYINPUT54), .A3(new_n806), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n820), .A2(KEYINPUT55), .A3(new_n596), .A4(new_n817), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n819), .A2(new_n599), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n804), .B1(new_n822), .B2(new_n537), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n686), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n634), .A2(new_n637), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n628), .A2(KEYINPUT99), .A3(new_n632), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n641), .B1(new_n640), .B2(new_n631), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n633), .A2(new_n638), .A3(new_n642), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n803), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT116), .B1(new_n822), .B2(new_n830), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n819), .A2(new_n599), .A3(new_n821), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n533), .A2(new_n800), .A3(new_n802), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n643), .A2(new_n644), .A3(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n832), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n824), .A2(new_n831), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n795), .B1(new_n837), .B2(new_n616), .ZN(new_n838));
  INV_X1    g637(.A(new_n459), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n841), .A2(new_n452), .A3(new_n769), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G113gat), .B1(new_n843), .B2(new_n537), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n838), .A2(new_n839), .A3(new_n735), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n845), .A2(new_n739), .ZN(new_n846));
  INV_X1    g645(.A(G113gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n847), .A3(new_n730), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n844), .A2(new_n848), .ZN(G1340gat));
  OAI21_X1  g648(.A(G120gat), .B1(new_n843), .B2(new_n728), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n728), .A2(G120gat), .ZN(new_n851));
  XOR2_X1   g650(.A(new_n851), .B(KEYINPUT117), .Z(new_n852));
  NAND2_X1  g651(.A1(new_n846), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n853), .ZN(G1341gat));
  NAND3_X1  g653(.A1(new_n842), .A2(G127gat), .A3(new_n752), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT118), .ZN(new_n856));
  AOI21_X1  g655(.A(G127gat), .B1(new_n846), .B2(new_n752), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(G1342gat));
  NOR2_X1   g657(.A1(new_n281), .A2(new_n686), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n845), .A2(new_n292), .A3(new_n859), .ZN(new_n860));
  XOR2_X1   g659(.A(new_n860), .B(KEYINPUT56), .Z(new_n861));
  OAI21_X1  g660(.A(G134gat), .B1(new_n843), .B2(new_n686), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1343gat));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n739), .A2(new_n651), .A3(new_n667), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n832), .A2(new_n730), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n645), .B1(new_n867), .B2(new_n804), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n836), .A2(new_n831), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n616), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n731), .A2(new_n728), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT57), .B1(new_n872), .B2(new_n447), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  AOI211_X1 g673(.A(new_n874), .B(new_n394), .C1(new_n870), .C2(new_n871), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n866), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n874), .B1(new_n838), .B2(new_n394), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n872), .A2(KEYINPUT57), .A3(new_n447), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(KEYINPUT119), .A3(new_n866), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n537), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(G141gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n864), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n838), .A2(new_n735), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT121), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n702), .A2(new_n394), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n889), .A2(new_n884), .A3(new_n730), .A4(new_n739), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT119), .B1(new_n881), .B2(new_n866), .ZN(new_n891));
  AOI211_X1 g690(.A(new_n877), .B(new_n865), .C1(new_n879), .C2(new_n880), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n730), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(KEYINPUT120), .A3(G141gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n885), .A2(new_n890), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT58), .ZN(new_n896));
  OAI21_X1  g695(.A(G141gat), .B1(new_n876), .B2(new_n537), .ZN(new_n897));
  XOR2_X1   g696(.A(KEYINPUT122), .B(KEYINPUT58), .Z(new_n898));
  NAND3_X1  g697(.A1(new_n890), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n896), .A2(new_n899), .ZN(G1344gat));
  INV_X1    g699(.A(G148gat), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n878), .A2(new_n882), .ZN(new_n902));
  AOI211_X1 g701(.A(KEYINPUT59), .B(new_n901), .C1(new_n902), .C2(new_n600), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n824), .B1(new_n822), .B2(new_n830), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n795), .B1(new_n904), .B2(new_n616), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n874), .B1(new_n905), .B2(new_n394), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n880), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n600), .ZN(new_n908));
  OAI21_X1  g707(.A(G148gat), .B1(new_n908), .B2(new_n865), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n909), .A2(KEYINPUT59), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n887), .A2(new_n739), .A3(new_n888), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n600), .A2(new_n901), .ZN(new_n912));
  OAI22_X1  g711(.A1(new_n903), .A2(new_n910), .B1(new_n911), .B2(new_n912), .ZN(G1345gat));
  NAND4_X1  g712(.A1(new_n889), .A2(KEYINPUT123), .A3(new_n752), .A4(new_n739), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n915), .B1(new_n911), .B2(new_n616), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n752), .ZN(new_n918));
  MUX2_X1   g717(.A(new_n917), .B(new_n918), .S(G155gat), .Z(G1346gat));
  INV_X1    g718(.A(G162gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n889), .A2(new_n920), .A3(new_n859), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n686), .B1(new_n878), .B2(new_n882), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n920), .ZN(G1347gat));
  NOR2_X1   g722(.A1(new_n739), .A2(new_n651), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n840), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n206), .A3(new_n730), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n840), .A2(new_n281), .A3(new_n735), .ZN(new_n927));
  OAI21_X1  g726(.A(G169gat), .B1(new_n927), .B2(new_n537), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(G1348gat));
  NAND3_X1  g728(.A1(new_n925), .A2(new_n207), .A3(new_n600), .ZN(new_n930));
  OAI21_X1  g729(.A(G176gat), .B1(new_n927), .B2(new_n728), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT124), .ZN(G1349gat));
  NAND3_X1  g732(.A1(new_n925), .A2(new_n752), .A3(new_n215), .ZN(new_n934));
  OAI21_X1  g733(.A(G183gat), .B1(new_n927), .B2(new_n616), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT60), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n934), .B(new_n935), .C1(KEYINPUT125), .C2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(KEYINPUT125), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n937), .B(new_n938), .ZN(G1350gat));
  OAI21_X1  g738(.A(G190gat), .B1(new_n927), .B2(new_n686), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT61), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n925), .A2(new_n210), .A3(new_n645), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1351gat));
  NOR3_X1   g742(.A1(new_n838), .A2(new_n394), .A3(new_n702), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n924), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n945), .A2(KEYINPUT126), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n945), .A2(KEYINPUT126), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(G197gat), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n730), .A2(new_n949), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n702), .A2(new_n660), .A3(new_n734), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n952), .B1(new_n880), .B2(new_n906), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n953), .A2(new_n730), .ZN(new_n954));
  OAI22_X1  g753(.A1(new_n948), .A2(new_n950), .B1(new_n949), .B2(new_n954), .ZN(G1352gat));
  NAND3_X1  g754(.A1(new_n944), .A2(new_n595), .A3(new_n924), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n957));
  OAI22_X1  g756(.A1(new_n956), .A2(new_n728), .B1(new_n957), .B2(KEYINPUT62), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT62), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(KEYINPUT127), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(G204gat), .B1(new_n908), .B2(new_n952), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n957), .B(KEYINPUT62), .C1(new_n956), .C2(new_n728), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(G1353gat));
  AOI21_X1  g762(.A(new_n249), .B1(new_n953), .B2(new_n752), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT63), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n752), .A2(new_n249), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n965), .B1(new_n948), .B2(new_n966), .ZN(G1354gat));
  OAI21_X1  g766(.A(new_n645), .B1(new_n946), .B2(new_n947), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n686), .A2(new_n248), .ZN(new_n969));
  AOI22_X1  g768(.A1(new_n968), .A2(new_n246), .B1(new_n953), .B2(new_n969), .ZN(G1355gat));
endmodule


