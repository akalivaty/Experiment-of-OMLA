//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0' ..
//Module:
 module locked_locked_c1908( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110,
    G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146,
    G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478,
    G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  , KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64);
input KEYINPUT64;
input KEYINPUT65;
input KEYINPUT66;
input KEYINPUT67;
input KEYINPUT68;
input KEYINPUT69;
input KEYINPUT70;
input KEYINPUT71;
input KEYINPUT72;
input KEYINPUT73;
input KEYINPUT74;
input KEYINPUT75;
input KEYINPUT76;
input KEYINPUT77;
input KEYINPUT78;
input KEYINPUT79;
input KEYINPUT80;
input KEYINPUT81;
input KEYINPUT82;
input KEYINPUT83;
input KEYINPUT84;
input KEYINPUT85;
input KEYINPUT86;
input KEYINPUT87;
input KEYINPUT88;
input KEYINPUT89;
input KEYINPUT90;
input KEYINPUT91;
input KEYINPUT92;
input KEYINPUT93;
input KEYINPUT94;
input KEYINPUT95;
input KEYINPUT96;
input KEYINPUT97;
input KEYINPUT98;
input KEYINPUT99;
input KEYINPUT100;
input KEYINPUT101;
input KEYINPUT102;
input KEYINPUT103;
input KEYINPUT104;
input KEYINPUT105;
input KEYINPUT106;
input KEYINPUT107;
input KEYINPUT108;
input KEYINPUT109;
input KEYINPUT110;
input KEYINPUT111;
input KEYINPUT112;
input KEYINPUT113;
input KEYINPUT114;
input KEYINPUT115;
input KEYINPUT116;
input KEYINPUT117;
input KEYINPUT118;
input KEYINPUT119;
input KEYINPUT120;
input KEYINPUT121;
input KEYINPUT122;
input KEYINPUT123;
input KEYINPUT124;
input KEYINPUT125;
input KEYINPUT126;
input KEYINPUT127;
//Header:
   input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104,
    G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140,
    G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472,
    G475, G478, G898, G900, G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n123, new_n124, new_n125, new_n126, new_n127, new_n128, new_n129,
    new_n130, new_n131, new_n132, new_n133, new_n134, new_n135, new_n136,
    new_n137, new_n138, new_n139, new_n140, new_n141, new_n142, new_n143,
    new_n144, new_n145, new_n146, new_n147, new_n148, new_n149, new_n150,
    new_n151, new_n152, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n190, new_n191, new_n192,
    new_n193, new_n194, new_n195, new_n196, new_n197, new_n198, new_n199,
    new_n200, new_n201, new_n202, new_n203, new_n204, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n260, new_n261, new_n262,
    new_n263, new_n264, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n322, new_n323, new_n324, new_n325,
    new_n326, new_n327, new_n328, new_n329, new_n330, new_n331, new_n332,
    new_n333, new_n334, new_n335, new_n336, new_n337, new_n338, new_n339,
    new_n340, new_n341, new_n342, new_n343, new_n344, new_n345, new_n346,
    new_n347, new_n348, new_n349, new_n350, new_n351, new_n352, new_n353,
    new_n354, new_n355, new_n356, new_n357, new_n358, new_n359, new_n360,
    new_n361, new_n362, new_n363, new_n364, new_n365, new_n366, new_n367,
    new_n368, new_n369, new_n370, new_n371, new_n372, new_n373, new_n374,
    new_n375, new_n376, new_n377, new_n378, new_n379, new_n380, new_n381,
    new_n382, new_n383, new_n384, new_n385, new_n386, new_n387, new_n388,
    new_n389, new_n390, new_n391, new_n392, new_n393, new_n394, new_n395,
    new_n396, new_n397, new_n398, new_n399, new_n400, new_n401, new_n402,
    new_n403, new_n404, new_n405, new_n406, new_n407, new_n408, new_n409,
    new_n410, new_n411, new_n412, new_n413, new_n414, new_n415, new_n416,
    new_n417, new_n418, new_n419, new_n420, new_n421, new_n422, new_n423,
    new_n424, new_n425, new_n426, new_n427, new_n428, new_n429, new_n430,
    new_n431, new_n432, new_n433, new_n434, new_n435, new_n436, new_n437,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n472, new_n473, new_n474, new_n475,
    new_n476, new_n477, new_n478, new_n479, new_n481, new_n482, new_n483,
    new_n484, new_n485, new_n486, new_n487, new_n489, new_n490, new_n491,
    new_n492, new_n493, new_n494, new_n495, new_n496, new_n497, new_n498,
    new_n499, new_n500, new_n501, new_n502, new_n504, new_n505, new_n506,
    new_n508, new_n509, new_n510, new_n511, new_n512, new_n513, new_n515,
    new_n517, new_n518, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755;
wire RLL_wire_A_64;
wire RLL_wire_A_65;
wire RLL_wire_A_66;
wire RLL_wire_A_67;
wire RLL_wire_A_68;
wire RLL_wire_A_69;
wire RLL_wire_A_70;
wire RLL_wire_A_71;
wire RLL_wire_A_72;
wire RLL_wire_A_73;
wire RLL_wire_A_74;
wire RLL_wire_A_75;
wire RLL_wire_A_76;
wire RLL_wire_A_77;
wire RLL_wire_A_78;
wire RLL_wire_A_79;
wire RLL_wire_A_80;
wire RLL_wire_A_81;
wire RLL_wire_A_82;
wire RLL_wire_A_83;
wire RLL_wire_A_84;
wire RLL_wire_A_85;
wire RLL_wire_A_86;
wire RLL_wire_A_87;
wire RLL_wire_A_88;
wire RLL_wire_A_89;
wire RLL_wire_A_90;
wire RLL_wire_A_91;
wire RLL_wire_A_92;
wire RLL_wire_A_93;
wire RLL_wire_A_94;
wire RLL_wire_A_95;
wire RLL_wire_A_96;
wire RLL_wire_A_97;
wire RLL_wire_A_98;
wire RLL_wire_A_99;
wire RLL_wire_A_100;
wire RLL_wire_A_101;
wire RLL_wire_A_102;
wire RLL_wire_A_103;
wire RLL_wire_A_104;
wire RLL_wire_A_105;
wire RLL_wire_A_106;
wire RLL_wire_A_107;
wire RLL_wire_A_108;
wire RLL_wire_A_109;
wire RLL_wire_A_110;
wire RLL_wire_A_111;
wire RLL_wire_A_112;
wire RLL_wire_A_113;
wire RLL_wire_A_114;
wire RLL_wire_A_115;
wire RLL_wire_A_116;
wire RLL_wire_A_117;
wire RLL_wire_A_118;
wire RLL_wire_A_119;
wire RLL_wire_A_120;
wire RLL_wire_A_121;
wire RLL_wire_A_122;
wire RLL_wire_A_123;
wire RLL_wire_A_124;
wire RLL_wire_A_125;
wire RLL_wire_A_126;
wire RLL_wire_A_127;

//Body:
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n123));
  OR2_X1    g001(.A1(KEYINPUT0), .A2(G128), .ZN(new_n124));
  NAND2_X1  g002(.A1(KEYINPUT0), .A2(G128), .ZN(new_n125));
  INV_X1    g003(.A(G143), .ZN(new_n126));
  NOR2_X1   g004(.A1(new_n126), .A2(G146), .ZN(new_n127));
  INV_X1    g005(.A(G146), .ZN(new_n128));
  NOR2_X1   g006(.A1(new_n128), .A2(G143), .ZN(new_n129));
  OAI211_X1 g007(.A(new_n124), .B(new_n125), .C1(new_n127), .C2(new_n129), .ZN(RLL_wire_A_64));
  XNOR2_X1 RLL_XNOR_64 (.A(RLL_wire_A_64), .B(KEYINPUT64), .ZN(new_n130) );
  NAND2_X1  g008(.A1(new_n128), .A2(G143), .ZN(new_n131));
  NAND2_X1  g009(.A1(new_n126), .A2(G146), .ZN(new_n132));
  NAND4_X1  g010(.A1(new_n131), .A2(new_n132), .A3(KEYINPUT0), .A4(G128), .ZN(new_n133));
  NAND2_X1  g011(.A1(new_n130), .A2(new_n133), .ZN(RLL_wire_A_65));
  XNOR2_X1 RLL_XNOR_65 (.A(RLL_wire_A_65), .B(KEYINPUT65), .ZN(new_n134) );
  INV_X1    g012(.A(KEYINPUT11), .ZN(new_n135));
  INV_X1    g013(.A(G134), .ZN(new_n136));
  OAI21_X1  g014(.A(new_n135), .B1(new_n136), .B2(G137), .ZN(new_n137));
  INV_X1    g015(.A(G137), .ZN(new_n138));
  NAND3_X1  g016(.A1(new_n138), .A2(KEYINPUT11), .A3(G134), .ZN(new_n139));
  INV_X1    g017(.A(G131), .ZN(new_n140));
  NAND2_X1  g018(.A1(new_n136), .A2(G137), .ZN(new_n141));
  NAND4_X1  g019(.A1(new_n137), .A2(new_n139), .A3(new_n140), .A4(new_n141), .ZN(new_n142));
  NAND3_X1  g020(.A1(new_n137), .A2(new_n139), .A3(new_n141), .ZN(new_n143));
  NAND2_X1  g021(.A1(new_n143), .A2(G131), .ZN(new_n144));
  AOI21_X1  g022(.A(new_n134), .B1(new_n142), .B2(new_n144), .ZN(new_n145));
  NOR2_X1   g023(.A1(new_n136), .A2(G137), .ZN(RLL_wire_A_66));
  XOR2_X1 RLL_XOR_66 (.A(RLL_wire_A_66), .B(KEYINPUT66), .Z(new_n146) );
  NOR2_X1   g024(.A1(new_n138), .A2(G134), .ZN(RLL_wire_A_67));
  XNOR2_X1 RLL_XNOR_67 (.A(RLL_wire_A_67), .B(KEYINPUT67), .ZN(new_n147) );
  OAI21_X1  g025(.A(G131), .B1(new_n146), .B2(new_n147), .ZN(new_n148));
  NAND2_X1  g026(.A1(new_n142), .A2(new_n148), .ZN(new_n149));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n150));
  NAND4_X1  g028(.A1(new_n131), .A2(new_n132), .A3(new_n150), .A4(G128), .ZN(new_n151));
  AOI21_X1  g029(.A(new_n150), .B1(G143), .B2(new_n128), .ZN(RLL_wire_A_68));
  XNOR2_X1 RLL_XNOR_68 (.A(RLL_wire_A_68), .B(KEYINPUT68), .ZN(new_n152) );
  INV_X1    g030(.A(G128), .ZN(new_n153));
  OAI22_X1  g031(.A1(new_n152), .A2(new_n153), .B1(new_n127), .B2(new_n129), .ZN(new_n154));
  AOI21_X1  g032(.A(new_n149), .B1(new_n151), .B2(new_n154), .ZN(new_n155));
  OAI21_X1  g033(.A(new_n123), .B1(new_n145), .B2(new_n155), .ZN(new_n156));
  OR2_X1    g034(.A1(KEYINPUT2), .A2(G113), .ZN(new_n157));
  NAND2_X1  g035(.A1(KEYINPUT2), .A2(G113), .ZN(new_n158));
  NAND2_X1  g036(.A1(new_n157), .A2(new_n158), .ZN(new_n159));
  INV_X1    g037(.A(G119), .ZN(new_n160));
  NAND2_X1  g038(.A1(new_n160), .A2(G116), .ZN(new_n161));
  INV_X1    g039(.A(G116), .ZN(new_n162));
  NAND2_X1  g040(.A1(new_n162), .A2(G119), .ZN(RLL_wire_A_69));
  XOR2_X1 RLL_XOR_69 (.A(RLL_wire_A_69), .B(KEYINPUT69), .Z(new_n163) );
  NAND2_X1  g041(.A1(new_n161), .A2(new_n163), .ZN(new_n164));
  NAND2_X1  g042(.A1(new_n159), .A2(new_n164), .ZN(new_n165));
  NAND4_X1  g043(.A1(new_n157), .A2(new_n161), .A3(new_n163), .A4(new_n158), .ZN(new_n166));
  NAND2_X1  g044(.A1(new_n165), .A2(new_n166), .ZN(new_n167));
  AND2_X1   g045(.A1(new_n130), .A2(new_n133), .ZN(new_n168));
  NAND2_X1  g046(.A1(new_n144), .A2(new_n142), .ZN(new_n169));
  NAND2_X1  g047(.A1(new_n168), .A2(new_n169), .ZN(new_n170));
  AND2_X1   g048(.A1(new_n142), .A2(new_n148), .ZN(new_n171));
  NAND2_X1  g049(.A1(new_n154), .A2(new_n151), .ZN(new_n172));
  NAND2_X1  g050(.A1(new_n171), .A2(new_n172), .ZN(new_n173));
  NAND3_X1  g051(.A1(new_n170), .A2(KEYINPUT30), .A3(new_n173), .ZN(new_n174));
  NAND3_X1  g052(.A1(new_n156), .A2(new_n167), .A3(new_n174), .ZN(new_n175));
  INV_X1    g053(.A(new_n167), .ZN(new_n176));
  NAND3_X1  g054(.A1(new_n170), .A2(new_n176), .A3(new_n173), .ZN(new_n177));
  INV_X1    g055(.A(G237), .ZN(new_n178));
  INV_X1    g056(.A(G953), .ZN(new_n179));
  NAND3_X1  g057(.A1(new_n178), .A2(new_n179), .A3(G210), .ZN(new_n180));
  XNOR2_X1  g058(.A(new_n180), .B(KEYINPUT27), .ZN(RLL_wire_A_70));
  XNOR2_X1 RLL_XNOR_70 (.A(RLL_wire_A_70), .B(KEYINPUT70), .ZN(new_n181) );
  XNOR2_X1  g059(.A(KEYINPUT26), .B(G101), .ZN(new_n182));
  XNOR2_X1  g060(.A(new_n181), .B(new_n182), .ZN(new_n183));
  AND2_X1   g061(.A1(new_n177), .A2(new_n183), .ZN(new_n184));
  NAND2_X1  g062(.A1(new_n175), .A2(new_n184), .ZN(new_n185));
  NAND2_X1  g063(.A1(new_n185), .A2(KEYINPUT31), .ZN(new_n186));
  INV_X1    g064(.A(KEYINPUT31), .ZN(new_n187));
  NAND3_X1  g065(.A1(new_n175), .A2(new_n184), .A3(new_n187), .ZN(RLL_wire_A_71));
  XNOR2_X1 RLL_XNOR_71 (.A(RLL_wire_A_71), .B(KEYINPUT71), .ZN(new_n188) );
  INV_X1    g066(.A(new_n183), .ZN(new_n189));
  INV_X1    g067(.A(KEYINPUT28), .ZN(new_n190));
  OAI21_X1  g068(.A(new_n167), .B1(new_n145), .B2(new_n155), .ZN(new_n191));
  AOI21_X1  g069(.A(new_n190), .B1(new_n191), .B2(new_n177), .ZN(new_n192));
  AOI22_X1  g070(.A1(new_n169), .A2(new_n168), .B1(new_n171), .B2(new_n172), .ZN(new_n193));
  AOI21_X1  g071(.A(KEYINPUT28), .B1(new_n193), .B2(new_n176), .ZN(new_n194));
  OAI21_X1  g072(.A(new_n189), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  NAND3_X1  g073(.A1(new_n186), .A2(new_n188), .A3(new_n195), .ZN(new_n196));
  NOR2_X1   g074(.A1(G472), .A2(G902), .ZN(new_n197));
  NAND2_X1  g075(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g076(.A(KEYINPUT32), .ZN(new_n199));
  NAND2_X1  g077(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NOR3_X1   g078(.A1(new_n192), .A2(new_n189), .A3(new_n194), .ZN(new_n201));
  AOI21_X1  g079(.A(new_n183), .B1(new_n175), .B2(new_n177), .ZN(new_n202));
  NOR3_X1   g080(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT29), .ZN(new_n203));
  INV_X1    g081(.A(new_n177), .ZN(new_n204));
  AOI21_X1  g082(.A(new_n176), .B1(new_n170), .B2(new_n173), .ZN(new_n205));
  OAI21_X1  g083(.A(KEYINPUT28), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g084(.A(new_n194), .ZN(new_n207));
  NAND4_X1  g085(.A1(new_n206), .A2(KEYINPUT29), .A3(new_n183), .A4(new_n207), .ZN(new_n208));
  INV_X1    g086(.A(G902), .ZN(new_n209));
  NAND2_X1  g087(.A1(new_n208), .A2(new_n209), .ZN(RLL_wire_A_72));
  XNOR2_X1 RLL_XNOR_72 (.A(RLL_wire_A_72), .B(KEYINPUT72), .ZN(new_n210) );
  OAI21_X1  g088(.A(G472), .B1(new_n203), .B2(new_n210), .ZN(new_n211));
  NAND3_X1  g089(.A1(new_n196), .A2(KEYINPUT32), .A3(new_n197), .ZN(new_n212));
  NAND3_X1  g090(.A1(new_n200), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g091(.A(G217), .ZN(new_n214));
  AOI21_X1  g092(.A(new_n214), .B1(G234), .B2(new_n209), .ZN(new_n215));
  INV_X1    g093(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g094(.A1(new_n153), .A2(G119), .ZN(RLL_wire_A_73));
  XNOR2_X1 RLL_XNOR_73 (.A(RLL_wire_A_73), .B(KEYINPUT73), .ZN(new_n217) );
  NAND2_X1  g095(.A1(new_n160), .A2(G128), .ZN(new_n218));
  NAND2_X1  g096(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g097(.A(KEYINPUT24), .B(G110), .ZN(new_n220));
  OR2_X1    g098(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g099(.A1(new_n153), .A2(KEYINPUT23), .A3(G119), .ZN(new_n222));
  INV_X1    g100(.A(KEYINPUT23), .ZN(new_n223));
  AOI21_X1  g101(.A(new_n223), .B1(new_n160), .B2(G128), .ZN(RLL_wire_A_74));
  XOR2_X1 RLL_XOR_74 (.A(RLL_wire_A_74), .B(KEYINPUT74), .Z(new_n224) );
  NOR2_X1   g102(.A1(new_n160), .A2(G128), .ZN(new_n225));
  OAI21_X1  g103(.A(new_n222), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g104(.A1(new_n226), .A2(G110), .ZN(RLL_wire_A_75));
  XOR2_X1 RLL_XOR_75 (.A(RLL_wire_A_75), .B(KEYINPUT75), .Z(new_n227) );
  INV_X1    g105(.A(G140), .ZN(new_n228));
  NAND2_X1  g106(.A1(new_n228), .A2(G125), .ZN(new_n229));
  INV_X1    g107(.A(G125), .ZN(new_n230));
  NAND2_X1  g108(.A1(new_n230), .A2(G140), .ZN(new_n231));
  NAND3_X1  g109(.A1(new_n229), .A2(new_n231), .A3(KEYINPUT16), .ZN(new_n232));
  OR3_X1    g110(.A1(new_n230), .A2(KEYINPUT16), .A3(G140), .ZN(new_n233));
  AND3_X1   g111(.A1(new_n232), .A2(G146), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g112(.A(G146), .B1(new_n232), .B2(new_n233), .ZN(RLL_wire_A_76));
  XOR2_X1 RLL_XOR_76 (.A(RLL_wire_A_76), .B(KEYINPUT76), .Z(new_n235) );
  OAI211_X1 g113(.A(new_n221), .B(new_n227), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  INV_X1    g114(.A(G110), .ZN(new_n237));
  OAI211_X1 g115(.A(new_n237), .B(new_n222), .C1(new_n224), .C2(new_n225), .ZN(new_n238));
  NAND2_X1  g116(.A1(new_n219), .A2(new_n220), .ZN(new_n239));
  NAND2_X1  g117(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g118(.A1(new_n232), .A2(new_n233), .A3(G146), .ZN(RLL_wire_A_77));
  XNOR2_X1 RLL_XNOR_77 (.A(RLL_wire_A_77), .B(KEYINPUT77), .ZN(new_n241) );
  XNOR2_X1  g119(.A(G125), .B(G140), .ZN(new_n242));
  NAND2_X1  g120(.A1(new_n242), .A2(new_n128), .ZN(new_n243));
  NAND3_X1  g121(.A1(new_n240), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g122(.A1(new_n236), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g123(.A(KEYINPUT22), .B(G137), .ZN(new_n246));
  NAND3_X1  g124(.A1(new_n179), .A2(G221), .A3(G234), .ZN(new_n247));
  XNOR2_X1  g125(.A(new_n246), .B(new_n247), .ZN(RLL_wire_A_78));
  XNOR2_X1 RLL_XNOR_78 (.A(RLL_wire_A_78), .B(KEYINPUT78), .ZN(new_n248) );
  INV_X1    g126(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g127(.A1(new_n245), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g128(.A1(new_n236), .A2(new_n244), .A3(new_n248), .ZN(new_n251));
  NAND3_X1  g129(.A1(new_n250), .A2(new_n209), .A3(new_n251), .ZN(new_n252));
  INV_X1    g130(.A(KEYINPUT25), .ZN(new_n253));
  NAND2_X1  g131(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g132(.A1(new_n250), .A2(KEYINPUT25), .A3(new_n209), .A4(new_n251), .ZN(new_n255));
  AOI21_X1  g133(.A(new_n216), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g134(.A1(new_n250), .A2(new_n251), .ZN(new_n257));
  NOR2_X1   g135(.A1(new_n215), .A2(G902), .ZN(new_n258));
  INV_X1    g136(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g137(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g138(.A1(new_n256), .A2(new_n260), .ZN(RLL_wire_A_79));
  XOR2_X1 RLL_XOR_79 (.A(RLL_wire_A_79), .B(KEYINPUT79), .Z(new_n261) );
  NAND2_X1  g139(.A1(new_n213), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g140(.A(KEYINPUT9), .B(G234), .ZN(new_n263));
  OAI21_X1  g141(.A(G221), .B1(new_n263), .B2(G902), .ZN(RLL_wire_A_80));
  XOR2_X1 RLL_XOR_80 (.A(RLL_wire_A_80), .B(KEYINPUT80), .Z(new_n264) );
  INV_X1    g142(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g143(.A(G110), .B(G140), .ZN(new_n266));
  AND2_X1   g144(.A1(new_n179), .A2(G227), .ZN(new_n267));
  XOR2_X1   g145(.A(new_n266), .B(new_n267), .Z(new_n268));
  INV_X1    g146(.A(new_n268), .ZN(new_n269));
  INV_X1    g147(.A(G104), .ZN(new_n270));
  OAI21_X1  g148(.A(KEYINPUT3), .B1(new_n270), .B2(G107), .ZN(RLL_wire_A_81));
  XNOR2_X1 RLL_XNOR_81 (.A(RLL_wire_A_81), .B(KEYINPUT81), .ZN(new_n271) );
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n272));
  INV_X1    g150(.A(G107), .ZN(new_n273));
  NAND3_X1  g151(.A1(new_n272), .A2(new_n273), .A3(G104), .ZN(new_n274));
  NAND2_X1  g152(.A1(new_n270), .A2(G107), .ZN(new_n275));
  NAND3_X1  g153(.A1(new_n271), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g154(.A1(new_n276), .A2(G101), .ZN(new_n277));
  INV_X1    g155(.A(G101), .ZN(new_n278));
  NAND4_X1  g156(.A1(new_n271), .A2(new_n274), .A3(new_n278), .A4(new_n275), .ZN(new_n279));
  NAND3_X1  g157(.A1(new_n277), .A2(KEYINPUT4), .A3(new_n279), .ZN(new_n280));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n281));
  NAND3_X1  g159(.A1(new_n276), .A2(new_n281), .A3(G101), .ZN(new_n282));
  NAND3_X1  g160(.A1(new_n280), .A2(new_n168), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g161(.A1(new_n270), .A2(G107), .ZN(RLL_wire_A_82));
  XNOR2_X1 RLL_XNOR_82 (.A(RLL_wire_A_82), .B(KEYINPUT82), .ZN(new_n284) );
  NOR2_X1   g162(.A1(new_n273), .A2(G104), .ZN(new_n285));
  OAI21_X1  g163(.A(G101), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g164(.A(new_n151), .ZN(new_n287));
  OAI21_X1  g165(.A(KEYINPUT1), .B1(new_n126), .B2(G146), .ZN(new_n288));
  AOI22_X1  g166(.A1(new_n288), .A2(G128), .B1(new_n131), .B2(new_n132), .ZN(new_n289));
  OAI211_X1 g167(.A(new_n279), .B(new_n286), .C1(new_n287), .C2(new_n289), .ZN(new_n290));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n291));
  NAND2_X1  g169(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g170(.A1(new_n279), .A2(new_n286), .ZN(new_n293));
  INV_X1    g171(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g172(.A1(new_n294), .A2(new_n172), .A3(KEYINPUT10), .ZN(new_n295));
  INV_X1    g173(.A(new_n169), .ZN(new_n296));
  NAND4_X1  g174(.A1(new_n283), .A2(new_n292), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  INV_X1    g175(.A(KEYINPUT12), .ZN(RLL_wire_A_83));
  XOR2_X1 RLL_XOR_83 (.A(RLL_wire_A_83), .B(KEYINPUT83), .Z(new_n298) );
  NAND3_X1  g176(.A1(new_n293), .A2(new_n151), .A3(new_n154), .ZN(new_n299));
  AOI221_X4 g177(.A(new_n298), .B1(new_n142), .B2(new_n144), .C1(new_n299), .C2(new_n290), .ZN(new_n300));
  NAND2_X1  g178(.A1(new_n299), .A2(new_n290), .ZN(new_n301));
  AOI21_X1  g179(.A(KEYINPUT12), .B1(new_n301), .B2(new_n169), .ZN(new_n302));
  OAI21_X1  g180(.A(new_n297), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g181(.A1(new_n297), .A2(new_n268), .ZN(new_n304));
  NAND3_X1  g182(.A1(new_n283), .A2(new_n292), .A3(new_n295), .ZN(new_n305));
  NAND2_X1  g183(.A1(new_n305), .A2(new_n169), .ZN(new_n306));
  AOI22_X1  g184(.A1(new_n269), .A2(new_n303), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g185(.A(G469), .B1(new_n307), .B2(G902), .ZN(new_n308));
  INV_X1    g186(.A(G469), .ZN(new_n309));
  NOR2_X1   g187(.A1(new_n300), .A2(new_n302), .ZN(new_n310));
  NAND2_X1  g188(.A1(new_n297), .A2(new_n268), .ZN(new_n311));
  NOR2_X1   g189(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g190(.A(new_n268), .B1(new_n306), .B2(new_n297), .ZN(new_n313));
  OAI211_X1 g191(.A(new_n309), .B(new_n209), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  AOI21_X1  g192(.A(new_n265), .B1(new_n308), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g193(.A(G214), .B1(G237), .B2(G902), .ZN(new_n316));
  INV_X1    g194(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g195(.A1(new_n280), .A2(new_n167), .A3(new_n282), .ZN(new_n318));
  INV_X1    g196(.A(KEYINPUT5), .ZN(new_n319));
  NAND3_X1  g197(.A1(new_n319), .A2(new_n160), .A3(G116), .ZN(new_n320));
  OAI211_X1 g198(.A(G113), .B(new_n320), .C1(new_n164), .C2(new_n319), .ZN(new_n321));
  NAND3_X1  g199(.A1(new_n294), .A2(new_n166), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g200(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g201(.A(G110), .B(G122), .ZN(RLL_wire_A_84));
  XOR2_X1 RLL_XOR_84 (.A(RLL_wire_A_84), .B(KEYINPUT84), .Z(new_n324) );
  INV_X1    g202(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g203(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g204(.A1(new_n318), .A2(new_n322), .A3(new_n324), .ZN(new_n327));
  NAND3_X1  g205(.A1(new_n326), .A2(KEYINPUT6), .A3(new_n327), .ZN(new_n328));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n329));
  NAND3_X1  g207(.A1(new_n323), .A2(new_n329), .A3(new_n325), .ZN(new_n330));
  AOI21_X1  g208(.A(new_n230), .B1(new_n130), .B2(new_n133), .ZN(new_n331));
  INV_X1    g209(.A(new_n331), .ZN(new_n332));
  NAND3_X1  g210(.A1(new_n154), .A2(new_n230), .A3(new_n151), .ZN(new_n333));
  NAND2_X1  g211(.A1(new_n332), .A2(new_n333), .ZN(RLL_wire_A_85));
  XOR2_X1 RLL_XOR_85 (.A(RLL_wire_A_85), .B(KEYINPUT85), .Z(new_n334) );
  INV_X1    g212(.A(G224), .ZN(new_n335));
  NOR2_X1   g213(.A1(new_n335), .A2(G953), .ZN(new_n336));
  XNOR2_X1  g214(.A(new_n334), .B(new_n336), .ZN(new_n337));
  NAND3_X1  g215(.A1(new_n328), .A2(new_n330), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g216(.A(new_n324), .B(KEYINPUT8), .ZN(new_n339));
  AND3_X1   g217(.A1(new_n161), .A2(new_n163), .A3(KEYINPUT5), .ZN(new_n340));
  NAND2_X1  g218(.A1(new_n320), .A2(G113), .ZN(new_n341));
  OAI21_X1  g219(.A(new_n166), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g220(.A1(new_n342), .A2(new_n293), .ZN(new_n343));
  AOI22_X1  g221(.A1(new_n321), .A2(new_n166), .B1(new_n279), .B2(new_n286), .ZN(new_n344));
  OAI21_X1  g222(.A(new_n339), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g223(.A(new_n333), .ZN(new_n346));
  INV_X1    g224(.A(KEYINPUT7), .ZN(new_n347));
  OAI22_X1  g225(.A1(new_n346), .A2(new_n331), .B1(new_n347), .B2(new_n336), .ZN(new_n348));
  INV_X1    g226(.A(new_n336), .ZN(RLL_wire_A_86));
  XNOR2_X1 RLL_XNOR_86 (.A(RLL_wire_A_86), .B(KEYINPUT86), .ZN(new_n349) );
  NAND4_X1  g227(.A1(new_n332), .A2(KEYINPUT7), .A3(new_n349), .A4(new_n333), .ZN(new_n350));
  AND3_X1   g228(.A1(new_n345), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g229(.A(G902), .B1(new_n351), .B2(new_n327), .ZN(new_n352));
  NAND2_X1  g230(.A1(new_n338), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g231(.A(G210), .B1(G237), .B2(G902), .ZN(new_n354));
  INV_X1    g232(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g233(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g234(.A1(new_n338), .A2(new_n352), .A3(new_n354), .ZN(new_n357));
  AOI21_X1  g235(.A(new_n317), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g236(.A(KEYINPUT20), .ZN(new_n359));
  NAND3_X1  g237(.A1(new_n178), .A2(new_n179), .A3(G214), .ZN(new_n360));
  NAND2_X1  g238(.A1(new_n360), .A2(new_n126), .ZN(RLL_wire_A_87));
  XOR2_X1 RLL_XOR_87 (.A(RLL_wire_A_87), .B(KEYINPUT87), .Z(new_n361) );
  NAND4_X1  g239(.A1(new_n178), .A2(new_n179), .A3(G143), .A4(G214), .ZN(new_n362));
  NAND2_X1  g240(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g241(.A1(new_n363), .A2(KEYINPUT18), .A3(G131), .ZN(new_n364));
  NAND2_X1  g242(.A1(new_n229), .A2(new_n231), .ZN(new_n365));
  NAND2_X1  g243(.A1(new_n365), .A2(G146), .ZN(new_n366));
  NAND2_X1  g244(.A1(new_n366), .A2(new_n243), .ZN(new_n367));
  NAND2_X1  g245(.A1(KEYINPUT18), .A2(G131), .ZN(new_n368));
  NAND3_X1  g246(.A1(new_n361), .A2(new_n362), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g247(.A1(new_n364), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  AND3_X1   g248(.A1(new_n361), .A2(new_n140), .A3(new_n362), .ZN(new_n371));
  AOI21_X1  g249(.A(new_n140), .B1(new_n361), .B2(new_n362), .ZN(new_n372));
  NOR2_X1   g250(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g251(.A1(new_n365), .A2(KEYINPUT19), .ZN(RLL_wire_A_88));
  XNOR2_X1 RLL_XNOR_88 (.A(RLL_wire_A_88), .B(KEYINPUT88), .ZN(new_n374) );
  INV_X1    g252(.A(KEYINPUT19), .ZN(RLL_wire_A_89));
  XNOR2_X1 RLL_XNOR_89 (.A(RLL_wire_A_89), .B(KEYINPUT89), .ZN(new_n375) );
  NAND2_X1  g253(.A1(new_n242), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g254(.A1(new_n374), .A2(new_n376), .A3(new_n128), .ZN(new_n377));
  NAND2_X1  g255(.A1(new_n377), .A2(new_n241), .ZN(new_n378));
  OAI21_X1  g256(.A(new_n370), .B1(new_n373), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g257(.A(G113), .B(G122), .ZN(new_n380));
  XNOR2_X1  g258(.A(new_n380), .B(G104), .ZN(new_n381));
  NAND2_X1  g259(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g260(.A(new_n381), .ZN(new_n383));
  NOR2_X1   g261(.A1(new_n234), .A2(new_n235), .ZN(new_n384));
  NAND2_X1  g262(.A1(new_n372), .A2(KEYINPUT17), .ZN(new_n385));
  NAND2_X1  g263(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR3_X1   g264(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT17), .ZN(new_n387));
  OAI211_X1 g265(.A(new_n383), .B(new_n370), .C1(new_n386), .C2(new_n387), .ZN(RLL_wire_A_90));
  XNOR2_X1 RLL_XNOR_90 (.A(RLL_wire_A_90), .B(KEYINPUT90), .ZN(new_n388) );
  NAND2_X1  g266(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g267(.A1(G475), .A2(G902), .ZN(new_n390));
  AOI21_X1  g268(.A(new_n359), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g269(.A(new_n390), .ZN(new_n392));
  AOI211_X1 g270(.A(KEYINPUT20), .B(new_n392), .C1(new_n382), .C2(new_n388), .ZN(new_n393));
  INV_X1    g271(.A(G475), .ZN(new_n394));
  OAI21_X1  g272(.A(new_n370), .B1(new_n386), .B2(new_n387), .ZN(new_n395));
  NAND2_X1  g273(.A1(new_n395), .A2(new_n381), .ZN(new_n396));
  AOI21_X1  g274(.A(G902), .B1(new_n396), .B2(new_n388), .ZN(new_n397));
  OAI22_X1  g275(.A1(new_n391), .A2(new_n393), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  INV_X1    g276(.A(G122), .ZN(new_n399));
  NAND2_X1  g277(.A1(new_n399), .A2(G116), .ZN(new_n400));
  NAND2_X1  g278(.A1(new_n162), .A2(G122), .ZN(new_n401));
  AND2_X1   g279(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g280(.A(new_n402), .B(new_n273), .ZN(new_n403));
  NAND2_X1  g281(.A1(new_n126), .A2(G128), .ZN(new_n404));
  INV_X1    g282(.A(KEYINPUT13), .ZN(new_n405));
  NAND2_X1  g283(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g284(.A1(new_n153), .A2(G143), .ZN(new_n407));
  NAND2_X1  g285(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g286(.A1(new_n404), .A2(new_n405), .ZN(new_n409));
  OAI21_X1  g287(.A(G134), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AND2_X1   g288(.A1(new_n404), .A2(new_n407), .ZN(new_n411));
  NAND2_X1  g289(.A1(new_n411), .A2(new_n136), .ZN(new_n412));
  NAND3_X1  g290(.A1(new_n403), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g291(.A(new_n411), .B(new_n136), .ZN(RLL_wire_A_91));
  XNOR2_X1 RLL_XNOR_91 (.A(RLL_wire_A_91), .B(KEYINPUT91), .ZN(new_n414) );
  NAND2_X1  g292(.A1(new_n402), .A2(new_n273), .ZN(new_n415));
  NAND2_X1  g293(.A1(new_n401), .A2(KEYINPUT14), .ZN(new_n416));
  NAND2_X1  g294(.A1(new_n416), .A2(new_n400), .ZN(new_n417));
  NOR2_X1   g295(.A1(new_n401), .A2(KEYINPUT14), .ZN(RLL_wire_A_92));
  XOR2_X1 RLL_XOR_92 (.A(RLL_wire_A_92), .B(KEYINPUT92), .Z(new_n418) );
  OAI21_X1  g296(.A(G107), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g297(.A1(new_n414), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  NOR3_X1   g298(.A1(new_n263), .A2(new_n214), .A3(G953), .ZN(new_n421));
  AND3_X1   g299(.A1(new_n413), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g300(.A(new_n421), .B1(new_n413), .B2(new_n420), .ZN(new_n423));
  OAI21_X1  g301(.A(new_n209), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g302(.A(KEYINPUT15), .ZN(new_n425));
  NAND3_X1  g303(.A1(new_n424), .A2(new_n425), .A3(G478), .ZN(new_n426));
  NAND2_X1  g304(.A1(new_n425), .A2(G478), .ZN(new_n427));
  OAI211_X1 g305(.A(new_n209), .B(new_n427), .C1(new_n422), .C2(new_n423), .ZN(new_n428));
  NAND2_X1  g306(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g307(.A(G952), .ZN(new_n430));
  AOI211_X1 g308(.A(G953), .B(new_n430), .C1(G234), .C2(G237), .ZN(new_n431));
  AOI211_X1 g309(.A(new_n209), .B(new_n179), .C1(G234), .C2(G237), .ZN(new_n432));
  XNOR2_X1  g310(.A(KEYINPUT21), .B(G898), .ZN(new_n433));
  AOI21_X1  g311(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NOR3_X1   g312(.A1(new_n398), .A2(new_n429), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g313(.A1(new_n315), .A2(new_n358), .A3(new_n435), .ZN(new_n436));
  NOR2_X1   g314(.A1(new_n262), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g315(.A(new_n437), .B(new_n278), .ZN(G3));
  NAND2_X1  g316(.A1(new_n196), .A2(new_n209), .ZN(RLL_wire_A_93));
  XOR2_X1 RLL_XOR_93 (.A(RLL_wire_A_93), .B(KEYINPUT93), .Z(new_n439) );
  NAND2_X1  g317(.A1(new_n439), .A2(G472), .ZN(new_n440));
  NAND4_X1  g318(.A1(new_n315), .A2(new_n198), .A3(new_n440), .A4(new_n261), .ZN(new_n441));
  INV_X1    g319(.A(new_n441), .ZN(RLL_wire_A_94));
  XOR2_X1 RLL_XOR_94 (.A(RLL_wire_A_94), .B(KEYINPUT94), .Z(new_n442) );
  AND3_X1   g320(.A1(new_n338), .A2(new_n352), .A3(new_n354), .ZN(new_n443));
  AOI21_X1  g321(.A(new_n354), .B1(new_n338), .B2(new_n352), .ZN(new_n444));
  OAI21_X1  g322(.A(new_n316), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g323(.A(KEYINPUT33), .ZN(new_n446));
  OAI21_X1  g324(.A(new_n446), .B1(new_n422), .B2(new_n423), .ZN(new_n447));
  NAND2_X1  g325(.A1(new_n413), .A2(new_n420), .ZN(new_n448));
  INV_X1    g326(.A(new_n421), .ZN(new_n449));
  NAND2_X1  g327(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g328(.A1(new_n413), .A2(new_n420), .A3(new_n421), .ZN(new_n451));
  NAND3_X1  g329(.A1(new_n450), .A2(KEYINPUT33), .A3(new_n451), .ZN(new_n452));
  NAND4_X1  g330(.A1(new_n447), .A2(new_n452), .A3(G478), .A4(new_n209), .ZN(new_n453));
  INV_X1    g331(.A(G478), .ZN(new_n454));
  NAND2_X1  g332(.A1(new_n424), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g333(.A1(new_n453), .A2(new_n455), .ZN(RLL_wire_A_95));
  XNOR2_X1 RLL_XNOR_95 (.A(RLL_wire_A_95), .B(KEYINPUT95), .ZN(new_n456) );
  NAND2_X1  g334(.A1(new_n398), .A2(new_n456), .ZN(new_n457));
  NOR3_X1   g335(.A1(new_n445), .A2(new_n457), .A3(new_n434), .ZN(new_n458));
  NAND2_X1  g336(.A1(new_n442), .A2(new_n458), .ZN(new_n459));
  XOR2_X1   g337(.A(KEYINPUT34), .B(G104), .Z(new_n460));
  XNOR2_X1  g338(.A(new_n459), .B(new_n460), .ZN(G6));
  INV_X1    g339(.A(new_n391), .ZN(new_n462));
  NAND3_X1  g340(.A1(new_n389), .A2(new_n359), .A3(new_n390), .ZN(new_n463));
  NAND2_X1  g341(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OR2_X1    g342(.A1(new_n397), .A2(new_n394), .ZN(new_n465));
  INV_X1    g343(.A(new_n434), .ZN(new_n466));
  NAND4_X1  g344(.A1(new_n464), .A2(new_n429), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  NOR2_X1   g345(.A1(new_n445), .A2(new_n467), .ZN(RLL_wire_A_96));
  XNOR2_X1 RLL_XNOR_96 (.A(RLL_wire_A_96), .B(KEYINPUT96), .ZN(new_n468) );
  NAND2_X1  g346(.A1(new_n442), .A2(new_n468), .ZN(new_n469));
  XOR2_X1   g347(.A(KEYINPUT35), .B(G107), .Z(new_n470));
  XNOR2_X1  g348(.A(new_n469), .B(new_n470), .ZN(G9));
  OR2_X1    g349(.A1(new_n249), .A2(KEYINPUT36), .ZN(new_n472));
  XNOR2_X1  g350(.A(new_n472), .B(new_n245), .ZN(new_n473));
  NOR2_X1   g351(.A1(new_n473), .A2(new_n259), .ZN(new_n474));
  NOR2_X1   g352(.A1(new_n256), .A2(new_n474), .ZN(new_n475));
  INV_X1    g353(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g354(.A1(new_n440), .A2(new_n198), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g355(.A1(new_n436), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g356(.A(KEYINPUT37), .B(G110), .ZN(new_n479));
  XNOR2_X1  g357(.A(new_n478), .B(new_n479), .ZN(G12));
  INV_X1    g358(.A(G900), .ZN(new_n481));
  NAND2_X1  g359(.A1(new_n432), .A2(new_n481), .ZN(new_n482));
  INV_X1    g360(.A(new_n431), .ZN(new_n483));
  NAND2_X1  g361(.A1(new_n482), .A2(new_n483), .ZN(RLL_wire_A_97));
  XOR2_X1 RLL_XOR_97 (.A(RLL_wire_A_97), .B(KEYINPUT97), .Z(new_n484) );
  NAND4_X1  g362(.A1(new_n464), .A2(new_n429), .A3(new_n465), .A4(new_n484), .ZN(new_n485));
  NOR2_X1   g363(.A1(new_n445), .A2(new_n485), .ZN(RLL_wire_A_98));
  XNOR2_X1 RLL_XNOR_98 (.A(RLL_wire_A_98), .B(KEYINPUT98), .ZN(new_n486) );
  NAND4_X1  g364(.A1(new_n486), .A2(new_n213), .A3(new_n315), .A4(new_n476), .ZN(new_n487));
  XNOR2_X1  g365(.A(new_n487), .B(G128), .ZN(G30));
  NAND2_X1  g366(.A1(new_n356), .A2(new_n357), .ZN(new_n489));
  INV_X1    g367(.A(KEYINPUT38), .ZN(RLL_wire_A_99));
  XNOR2_X1 RLL_XNOR_99 (.A(RLL_wire_A_99), .B(KEYINPUT99), .ZN(new_n490) );
  XNOR2_X1  g368(.A(new_n489), .B(new_n490), .ZN(new_n491));
  OAI21_X1  g369(.A(new_n189), .B1(new_n204), .B2(new_n205), .ZN(new_n492));
  AND2_X1   g370(.A1(new_n185), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g371(.A(G472), .B1(new_n493), .B2(G902), .ZN(new_n494));
  NAND3_X1  g372(.A1(new_n200), .A2(new_n212), .A3(new_n494), .ZN(new_n495));
  INV_X1    g373(.A(new_n495), .ZN(new_n496));
  NAND4_X1  g374(.A1(new_n475), .A2(new_n316), .A3(new_n398), .A4(new_n429), .ZN(new_n497));
  OR3_X1    g375(.A1(new_n491), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  XNOR2_X1  g376(.A(new_n484), .B(KEYINPUT39), .ZN(new_n499));
  NAND2_X1  g377(.A1(new_n315), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g378(.A(new_n500), .B(KEYINPUT40), .ZN(new_n501));
  NOR2_X1   g379(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g380(.A(new_n502), .B(new_n126), .ZN(G45));
  NAND3_X1  g381(.A1(new_n398), .A2(new_n456), .A3(new_n484), .ZN(new_n504));
  NOR2_X1   g382(.A1(new_n445), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g383(.A1(new_n505), .A2(new_n213), .A3(new_n315), .A4(new_n476), .ZN(new_n506));
  XNOR2_X1  g384(.A(new_n506), .B(G146), .ZN(G48));
  OAI21_X1  g385(.A(new_n209), .B1(new_n312), .B2(new_n313), .ZN(new_n508));
  NAND2_X1  g386(.A1(new_n508), .A2(G469), .ZN(new_n509));
  NAND3_X1  g387(.A1(new_n509), .A2(new_n264), .A3(new_n314), .ZN(new_n510));
  INV_X1    g388(.A(new_n510), .ZN(new_n511));
  NAND4_X1  g389(.A1(new_n458), .A2(new_n213), .A3(new_n261), .A4(new_n511), .ZN(new_n512));
  XNOR2_X1  g390(.A(KEYINPUT41), .B(G113), .ZN(new_n513));
  XNOR2_X1  g391(.A(new_n512), .B(new_n513), .ZN(G15));
  NAND4_X1  g392(.A1(new_n468), .A2(new_n213), .A3(new_n511), .A4(new_n261), .ZN(new_n515));
  XNOR2_X1  g393(.A(new_n515), .B(G116), .ZN(G18));
  NOR2_X1   g394(.A1(new_n510), .A2(new_n445), .ZN(new_n517));
  NAND4_X1  g395(.A1(new_n517), .A2(new_n213), .A3(new_n435), .A4(new_n476), .ZN(new_n518));
  XNOR2_X1  g396(.A(new_n518), .B(G119), .ZN(G21));
  INV_X1    g397(.A(new_n197), .ZN(new_n520));
  NAND2_X1  g398(.A1(new_n206), .A2(new_n207), .ZN(new_n521));
  AOI22_X1  g399(.A1(new_n521), .A2(new_n189), .B1(new_n185), .B2(KEYINPUT31), .ZN(RLL_wire_A_100));
  XNOR2_X1 RLL_XNOR_100 (.A(RLL_wire_A_100), .B(KEYINPUT100), .ZN(new_n522) );
  AOI21_X1  g400(.A(new_n520), .B1(new_n522), .B2(new_n188), .ZN(new_n523));
  INV_X1    g401(.A(G472), .ZN(new_n524));
  AOI21_X1  g402(.A(new_n524), .B1(new_n196), .B2(new_n209), .ZN(new_n525));
  OR2_X1    g403(.A1(new_n256), .A2(new_n260), .ZN(new_n526));
  NOR3_X1   g404(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g405(.A1(new_n398), .A2(new_n429), .ZN(new_n528));
  NOR2_X1   g406(.A1(new_n445), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g407(.A1(new_n527), .A2(new_n529), .A3(new_n466), .A4(new_n511), .ZN(RLL_wire_A_101));
  XNOR2_X1 RLL_XNOR_101 (.A(RLL_wire_A_101), .B(KEYINPUT101), .ZN(new_n530) );
  XNOR2_X1  g408(.A(new_n530), .B(G122), .ZN(G24));
  NOR3_X1   g409(.A1(new_n525), .A2(new_n523), .A3(new_n475), .ZN(new_n532));
  INV_X1    g410(.A(new_n504), .ZN(new_n533));
  NAND3_X1  g411(.A1(new_n517), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  XNOR2_X1  g412(.A(new_n534), .B(G125), .ZN(G27));
  NAND2_X1  g413(.A1(G469), .A2(G902), .ZN(new_n536));
  NAND2_X1  g414(.A1(new_n303), .A2(new_n269), .ZN(new_n537));
  NAND2_X1  g415(.A1(new_n304), .A2(new_n306), .ZN(new_n538));
  NAND3_X1  g416(.A1(new_n537), .A2(new_n538), .A3(G469), .ZN(new_n539));
  NAND3_X1  g417(.A1(new_n314), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g418(.A1(new_n540), .A2(new_n264), .ZN(RLL_wire_A_102));
  XOR2_X1 RLL_XOR_102 (.A(RLL_wire_A_102), .B(KEYINPUT102), .Z(new_n541) );
  NAND3_X1  g419(.A1(new_n356), .A2(new_n316), .A3(new_n357), .ZN(new_n542));
  NOR2_X1   g420(.A1(new_n541), .A2(new_n542), .ZN(RLL_wire_A_103));
  XOR2_X1 RLL_XOR_103 (.A(RLL_wire_A_103), .B(KEYINPUT103), .Z(new_n543) );
  NAND4_X1  g421(.A1(new_n543), .A2(new_n213), .A3(new_n261), .A4(new_n533), .ZN(new_n544));
  INV_X1    g422(.A(KEYINPUT42), .ZN(new_n545));
  NAND2_X1  g423(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AND3_X1   g424(.A1(new_n196), .A2(KEYINPUT32), .A3(new_n197), .ZN(new_n547));
  AOI21_X1  g425(.A(KEYINPUT32), .B1(new_n196), .B2(new_n197), .ZN(new_n548));
  NOR2_X1   g426(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g427(.A(new_n526), .B1(new_n549), .B2(new_n211), .ZN(RLL_wire_A_104));
  XNOR2_X1 RLL_XNOR_104 (.A(RLL_wire_A_104), .B(KEYINPUT104), .ZN(new_n550) );
  NAND4_X1  g428(.A1(new_n550), .A2(KEYINPUT42), .A3(new_n533), .A4(new_n543), .ZN(new_n551));
  NAND2_X1  g429(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g430(.A(new_n552), .B(G131), .ZN(G33));
  INV_X1    g431(.A(new_n485), .ZN(RLL_wire_A_105));
  XOR2_X1 RLL_XOR_105 (.A(RLL_wire_A_105), .B(KEYINPUT105), .Z(new_n554) );
  NAND4_X1  g432(.A1(new_n543), .A2(new_n213), .A3(new_n261), .A4(new_n554), .ZN(new_n555));
  XNOR2_X1  g433(.A(new_n555), .B(G134), .ZN(RLL_wire_A_106));
  XNOR2_X1 RLL_XNOR_106 (.A(RLL_wire_A_106), .B(KEYINPUT106), .ZN(G36) );
  OAI21_X1  g434(.A(G469), .B1(new_n307), .B2(KEYINPUT45), .ZN(new_n557));
  AND3_X1   g435(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT45), .ZN(new_n558));
  OR2_X1    g436(.A1(new_n557), .A2(new_n558), .ZN(RLL_wire_A_107));
  XOR2_X1 RLL_XOR_107 (.A(RLL_wire_A_107), .B(KEYINPUT107), .Z(new_n559) );
  NAND3_X1  g437(.A1(new_n559), .A2(KEYINPUT46), .A3(new_n536), .ZN(new_n560));
  NAND2_X1  g438(.A1(new_n560), .A2(new_n314), .ZN(new_n561));
  AOI21_X1  g439(.A(KEYINPUT46), .B1(new_n559), .B2(new_n536), .ZN(new_n562));
  OAI211_X1 g440(.A(new_n264), .B(new_n499), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  INV_X1    g441(.A(new_n563), .ZN(new_n564));
  INV_X1    g442(.A(KEYINPUT43), .ZN(new_n565));
  INV_X1    g443(.A(new_n456), .ZN(new_n566));
  OAI21_X1  g444(.A(new_n565), .B1(new_n566), .B2(new_n398), .ZN(new_n567));
  INV_X1    g445(.A(new_n398), .ZN(new_n568));
  NAND3_X1  g446(.A1(new_n568), .A2(KEYINPUT43), .A3(new_n456), .ZN(new_n569));
  NAND2_X1  g447(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g448(.A(new_n475), .B1(new_n440), .B2(new_n198), .ZN(new_n571));
  NAND3_X1  g449(.A1(new_n570), .A2(new_n571), .A3(KEYINPUT44), .ZN(new_n572));
  INV_X1    g450(.A(new_n542), .ZN(new_n573));
  NAND2_X1  g451(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g452(.A(KEYINPUT44), .B1(new_n570), .B2(new_n571), .ZN(new_n575));
  NOR2_X1   g453(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g454(.A1(new_n564), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g455(.A(new_n577), .B(G137), .ZN(RLL_wire_A_108));
  XOR2_X1 RLL_XOR_108 (.A(RLL_wire_A_108), .B(KEYINPUT108), .Z(G39) );
  OAI21_X1  g456(.A(new_n264), .B1(new_n561), .B2(new_n562), .ZN(new_n579));
  OR2_X1    g457(.A1(new_n579), .A2(KEYINPUT47), .ZN(new_n580));
  NAND2_X1  g458(.A1(new_n579), .A2(KEYINPUT47), .ZN(new_n581));
  NOR4_X1   g459(.A1(new_n213), .A2(new_n261), .A3(new_n504), .A4(new_n542), .ZN(new_n582));
  NAND3_X1  g460(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g461(.A(new_n583), .B(G140), .ZN(G42));
  NOR3_X1   g462(.A1(new_n526), .A2(new_n317), .A3(new_n265), .ZN(new_n585));
  NAND3_X1  g463(.A1(new_n585), .A2(new_n568), .A3(new_n456), .ZN(new_n586));
  NAND2_X1  g464(.A1(new_n509), .A2(new_n314), .ZN(new_n587));
  AOI21_X1  g465(.A(new_n586), .B1(KEYINPUT49), .B2(new_n587), .ZN(RLL_wire_A_109));
  XNOR2_X1 RLL_XNOR_109 (.A(RLL_wire_A_109), .B(KEYINPUT109), .ZN(new_n588) );
  OR2_X1    g466(.A1(new_n587), .A2(KEYINPUT49), .ZN(new_n589));
  NAND4_X1  g467(.A1(new_n588), .A2(new_n491), .A3(new_n496), .A4(new_n589), .ZN(RLL_wire_A_110));
  XOR2_X1 RLL_XOR_110 (.A(RLL_wire_A_110), .B(KEYINPUT110), .Z(new_n590) );
  AND4_X1   g468(.A1(new_n512), .A2(new_n530), .A3(new_n518), .A4(new_n515), .ZN(new_n591));
  AND2_X1   g469(.A1(new_n398), .A2(new_n456), .ZN(new_n592));
  NAND3_X1  g470(.A1(new_n358), .A2(new_n592), .A3(new_n466), .ZN(new_n593));
  OAI22_X1  g471(.A1(new_n262), .A2(new_n436), .B1(new_n441), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g472(.A1(new_n426), .A2(new_n428), .ZN(new_n595));
  NOR2_X1   g473(.A1(new_n595), .A2(new_n398), .ZN(new_n596));
  NAND3_X1  g474(.A1(new_n358), .A2(new_n466), .A3(new_n596), .ZN(new_n597));
  OAI22_X1  g475(.A1(new_n441), .A2(new_n597), .B1(new_n436), .B2(new_n477), .ZN(new_n598));
  NOR2_X1   g476(.A1(new_n594), .A2(new_n598), .ZN(RLL_wire_A_111));
  XOR2_X1 RLL_XOR_111 (.A(RLL_wire_A_111), .B(KEYINPUT111), .Z(new_n599) );
  NAND4_X1  g477(.A1(new_n595), .A2(new_n464), .A3(new_n465), .A4(new_n484), .ZN(new_n600));
  NOR2_X1   g478(.A1(new_n600), .A2(new_n542), .ZN(RLL_wire_A_112));
  XNOR2_X1 RLL_XNOR_112 (.A(RLL_wire_A_112), .B(KEYINPUT112), .ZN(new_n601) );
  NAND4_X1  g479(.A1(new_n601), .A2(new_n213), .A3(new_n315), .A4(new_n476), .ZN(new_n602));
  NAND3_X1  g480(.A1(new_n543), .A2(new_n532), .A3(new_n533), .ZN(new_n603));
  AND3_X1   g481(.A1(new_n555), .A2(new_n602), .A3(new_n603), .ZN(RLL_wire_A_113));
  XOR2_X1 RLL_XOR_113 (.A(RLL_wire_A_113), .B(KEYINPUT113), .Z(new_n604) );
  NAND4_X1  g482(.A1(new_n591), .A2(new_n552), .A3(new_n599), .A4(new_n604), .ZN(new_n605));
  INV_X1    g483(.A(new_n605), .ZN(new_n606));
  AND2_X1   g484(.A1(new_n487), .A2(new_n534), .ZN(new_n607));
  INV_X1    g485(.A(new_n484), .ZN(new_n608));
  NOR3_X1   g486(.A1(new_n256), .A2(new_n474), .A3(new_n608), .ZN(new_n609));
  AND3_X1   g487(.A1(new_n540), .A2(new_n609), .A3(new_n264), .ZN(new_n610));
  NAND3_X1  g488(.A1(new_n529), .A2(new_n495), .A3(new_n610), .ZN(new_n611));
  NAND4_X1  g489(.A1(new_n607), .A2(KEYINPUT52), .A3(new_n506), .A4(new_n611), .ZN(new_n612));
  NAND4_X1  g490(.A1(new_n487), .A2(new_n506), .A3(new_n534), .A4(new_n611), .ZN(new_n613));
  INV_X1    g491(.A(KEYINPUT52), .ZN(RLL_wire_A_114));
  XOR2_X1 RLL_XOR_114 (.A(RLL_wire_A_114), .B(KEYINPUT114), .Z(new_n614) );
  NAND2_X1  g492(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g493(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g494(.A(KEYINPUT53), .B1(new_n606), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g495(.A(new_n613), .B(KEYINPUT52), .ZN(new_n618));
  INV_X1    g496(.A(KEYINPUT53), .ZN(new_n619));
  NOR3_X1   g497(.A1(new_n618), .A2(new_n605), .A3(new_n619), .ZN(RLL_wire_A_115));
  XNOR2_X1 RLL_XNOR_115 (.A(RLL_wire_A_115), .B(KEYINPUT115), .ZN(new_n620) );
  OAI21_X1  g498(.A(KEYINPUT54), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g499(.A(new_n619), .B1(new_n618), .B2(new_n605), .ZN(new_n622));
  AND2_X1   g500(.A1(new_n599), .A2(new_n604), .ZN(new_n623));
  NAND4_X1  g501(.A1(new_n512), .A2(new_n530), .A3(new_n518), .A4(new_n515), .ZN(new_n624));
  AOI21_X1  g502(.A(new_n624), .B1(new_n546), .B2(new_n551), .ZN(new_n625));
  NAND4_X1  g503(.A1(new_n616), .A2(new_n623), .A3(KEYINPUT53), .A4(new_n625), .ZN(new_n626));
  INV_X1    g504(.A(KEYINPUT54), .ZN(new_n627));
  NAND3_X1  g505(.A1(new_n622), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g506(.A1(new_n621), .A2(new_n628), .ZN(new_n629));
  INV_X1    g507(.A(KEYINPUT51), .ZN(new_n630));
  AOI21_X1  g508(.A(new_n483), .B1(new_n567), .B2(new_n569), .ZN(new_n631));
  NAND3_X1  g509(.A1(new_n631), .A2(new_n527), .A3(new_n573), .ZN(new_n632));
  NAND2_X1  g510(.A1(new_n580), .A2(new_n581), .ZN(new_n633));
  INV_X1    g511(.A(new_n587), .ZN(new_n634));
  NAND2_X1  g512(.A1(new_n634), .A2(new_n265), .ZN(new_n635));
  AOI21_X1  g513(.A(new_n632), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g514(.A1(new_n510), .A2(new_n316), .ZN(new_n637));
  AND2_X1   g515(.A1(new_n491), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g516(.A1(new_n638), .A2(new_n527), .A3(new_n631), .ZN(new_n639));
  INV_X1    g517(.A(KEYINPUT50), .ZN(new_n640));
  NAND2_X1  g518(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g519(.A1(new_n638), .A2(KEYINPUT50), .A3(new_n527), .A4(new_n631), .ZN(new_n642));
  NAND2_X1  g520(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g521(.A1(new_n510), .A2(new_n542), .ZN(new_n644));
  AND2_X1   g522(.A1(new_n631), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g523(.A1(new_n645), .A2(new_n532), .ZN(new_n646));
  NAND4_X1  g524(.A1(new_n496), .A2(new_n261), .A3(new_n431), .A4(new_n644), .ZN(new_n647));
  OR3_X1    g525(.A1(new_n647), .A2(new_n398), .A3(new_n456), .ZN(new_n648));
  NAND3_X1  g526(.A1(new_n643), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g527(.A(new_n630), .B1(new_n636), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g528(.A1(new_n648), .A2(new_n646), .ZN(new_n651));
  AOI21_X1  g529(.A(new_n651), .B1(new_n642), .B2(new_n641), .ZN(new_n652));
  AOI22_X1  g530(.A1(new_n580), .A2(new_n581), .B1(new_n265), .B2(new_n634), .ZN(new_n653));
  OAI211_X1 g531(.A(new_n652), .B(KEYINPUT51), .C1(new_n653), .C2(new_n632), .ZN(new_n654));
  NOR2_X1   g532(.A1(new_n430), .A2(G953), .ZN(new_n655));
  NAND3_X1  g533(.A1(new_n631), .A2(new_n527), .A3(new_n517), .ZN(new_n656));
  OAI211_X1 g534(.A(new_n655), .B(new_n656), .C1(new_n647), .C2(new_n457), .ZN(new_n657));
  NAND2_X1  g535(.A1(new_n645), .A2(new_n550), .ZN(new_n658));
  OR2_X1    g536(.A1(new_n658), .A2(KEYINPUT48), .ZN(RLL_wire_A_116));
  XOR2_X1 RLL_XOR_116 (.A(RLL_wire_A_116), .B(KEYINPUT116), .Z(new_n659) );
  NAND2_X1  g537(.A1(new_n658), .A2(KEYINPUT48), .ZN(new_n660));
  AOI21_X1  g538(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g539(.A1(new_n650), .A2(new_n654), .A3(new_n661), .ZN(new_n662));
  NOR2_X1   g540(.A1(new_n629), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g541(.A1(G952), .A2(G953), .ZN(new_n664));
  OAI21_X1  g542(.A(new_n590), .B1(new_n663), .B2(new_n664), .ZN(G75));
  NAND2_X1  g543(.A1(new_n328), .A2(new_n330), .ZN(new_n666));
  XOR2_X1   g544(.A(new_n666), .B(new_n337), .Z(new_n667));
  XNOR2_X1  g545(.A(new_n667), .B(KEYINPUT55), .ZN(new_n668));
  AOI211_X1 g546(.A(new_n209), .B(new_n354), .C1(new_n622), .C2(new_n626), .ZN(new_n669));
  OAI21_X1  g547(.A(new_n668), .B1(new_n669), .B2(KEYINPUT56), .ZN(new_n670));
  AOI21_X1  g548(.A(new_n209), .B1(new_n622), .B2(new_n626), .ZN(new_n671));
  NAND2_X1  g549(.A1(new_n671), .A2(new_n355), .ZN(new_n672));
  INV_X1    g550(.A(KEYINPUT56), .ZN(new_n673));
  INV_X1    g551(.A(new_n668), .ZN(new_n674));
  NAND3_X1  g552(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g553(.A1(new_n179), .A2(G952), .ZN(RLL_wire_A_117));
  XNOR2_X1 RLL_XNOR_117 (.A(RLL_wire_A_117), .B(KEYINPUT117), .ZN(new_n676) );
  INV_X1    g554(.A(new_n676), .ZN(new_n677));
  AND3_X1   g555(.A1(new_n670), .A2(new_n675), .A3(new_n677), .ZN(G51));
  XOR2_X1   g556(.A(new_n536), .B(KEYINPUT57), .Z(new_n679));
  AND3_X1   g557(.A1(new_n622), .A2(new_n627), .A3(new_n626), .ZN(new_n680));
  AOI21_X1  g558(.A(new_n627), .B1(new_n622), .B2(new_n626), .ZN(RLL_wire_A_118));
  XNOR2_X1 RLL_XNOR_118 (.A(RLL_wire_A_118), .B(KEYINPUT118), .ZN(new_n681) );
  OAI21_X1  g559(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(RLL_wire_A_119));
  XOR2_X1 RLL_XOR_119 (.A(RLL_wire_A_119), .B(KEYINPUT119), .Z(new_n682) );
  OR2_X1    g560(.A1(new_n312), .A2(new_n313), .ZN(new_n683));
  NAND2_X1  g561(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g562(.A(new_n559), .ZN(new_n685));
  NAND2_X1  g563(.A1(new_n671), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g564(.A(new_n676), .B1(new_n684), .B2(new_n686), .ZN(G54));
  AND2_X1   g565(.A1(KEYINPUT58), .A2(G475), .ZN(new_n688));
  AND3_X1   g566(.A1(new_n671), .A2(new_n389), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g567(.A(new_n389), .B1(new_n671), .B2(new_n688), .ZN(RLL_wire_A_120));
  XOR2_X1 RLL_XOR_120 (.A(RLL_wire_A_120), .B(KEYINPUT120), .Z(new_n690) );
  NOR3_X1   g568(.A1(new_n689), .A2(new_n690), .A3(new_n676), .ZN(G60));
  AND2_X1   g569(.A1(new_n447), .A2(new_n452), .ZN(new_n692));
  NAND2_X1  g570(.A1(G478), .A2(G902), .ZN(new_n693));
  XNOR2_X1  g571(.A(new_n693), .B(KEYINPUT59), .ZN(new_n694));
  OAI211_X1 g572(.A(new_n692), .B(new_n694), .C1(new_n680), .C2(new_n681), .ZN(new_n695));
  NAND2_X1  g573(.A1(new_n695), .A2(new_n677), .ZN(new_n696));
  AOI21_X1  g574(.A(new_n692), .B1(new_n629), .B2(new_n694), .ZN(new_n697));
  NOR2_X1   g575(.A1(new_n696), .A2(new_n697), .ZN(G63));
  INV_X1    g576(.A(KEYINPUT61), .ZN(new_n699));
  NAND2_X1  g577(.A1(G217), .A2(G902), .ZN(new_n700));
  XOR2_X1   g578(.A(new_n700), .B(KEYINPUT60), .Z(new_n701));
  INV_X1    g579(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g580(.A(new_n702), .B1(new_n622), .B2(new_n626), .ZN(new_n703));
  INV_X1    g581(.A(new_n473), .ZN(new_n704));
  NAND2_X1  g582(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g583(.A(new_n705), .ZN(new_n706));
  INV_X1    g584(.A(new_n257), .ZN(new_n707));
  OAI21_X1  g585(.A(new_n677), .B1(new_n703), .B2(new_n707), .ZN(RLL_wire_A_121));
  XNOR2_X1 RLL_XNOR_121 (.A(RLL_wire_A_121), .B(KEYINPUT121), .ZN(new_n708) );
  OAI21_X1  g586(.A(new_n699), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  OR2_X1    g587(.A1(new_n703), .A2(new_n707), .ZN(new_n710));
  NAND4_X1  g588(.A1(new_n710), .A2(KEYINPUT61), .A3(new_n677), .A4(new_n705), .ZN(new_n711));
  NAND2_X1  g589(.A1(new_n709), .A2(new_n711), .ZN(G66));
  NAND2_X1  g590(.A1(new_n591), .A2(new_n599), .ZN(new_n713));
  NAND2_X1  g591(.A1(new_n713), .A2(new_n179), .ZN(new_n714));
  OAI21_X1  g592(.A(G953), .B1(new_n433), .B2(new_n335), .ZN(new_n715));
  NAND2_X1  g593(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g594(.A(new_n666), .B1(G898), .B2(new_n179), .ZN(new_n717));
  XNOR2_X1  g595(.A(new_n716), .B(new_n717), .ZN(RLL_wire_A_122));
  XNOR2_X1 RLL_XNOR_122 (.A(RLL_wire_A_122), .B(KEYINPUT122), .ZN(G69) );
  NAND2_X1  g596(.A1(new_n156), .A2(new_n174), .ZN(new_n719));
  AND2_X1   g597(.A1(new_n374), .A2(new_n376), .ZN(new_n720));
  XNOR2_X1  g598(.A(new_n719), .B(new_n720), .ZN(new_n721));
  INV_X1    g599(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g600(.A1(new_n607), .A2(new_n506), .ZN(RLL_wire_A_123));
  XNOR2_X1 RLL_XNOR_123 (.A(RLL_wire_A_123), .B(KEYINPUT123), .ZN(new_n723) );
  OR3_X1    g601(.A1(new_n502), .A2(new_n723), .A3(KEYINPUT62), .ZN(RLL_wire_A_124));
  XNOR2_X1 RLL_XNOR_124 (.A(RLL_wire_A_124), .B(KEYINPUT124), .ZN(new_n724) );
  OAI21_X1  g602(.A(KEYINPUT62), .B1(new_n502), .B2(new_n723), .ZN(new_n725));
  NOR2_X1   g603(.A1(new_n592), .A2(new_n596), .ZN(new_n726));
  NOR4_X1   g604(.A1(new_n262), .A2(new_n500), .A3(new_n726), .A4(new_n542), .ZN(new_n727));
  AOI21_X1  g605(.A(new_n727), .B1(new_n564), .B2(new_n576), .ZN(new_n728));
  NAND4_X1  g606(.A1(new_n724), .A2(new_n725), .A3(new_n583), .A4(new_n728), .ZN(new_n729));
  AOI21_X1  g607(.A(new_n722), .B1(new_n729), .B2(new_n179), .ZN(new_n730));
  INV_X1    g608(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g609(.A(new_n179), .B1(G227), .B2(G900), .ZN(new_n732));
  INV_X1    g610(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g611(.A1(new_n179), .A2(G900), .ZN(new_n734));
  AOI21_X1  g612(.A(new_n723), .B1(new_n576), .B2(new_n564), .ZN(new_n735));
  NAND3_X1  g613(.A1(new_n564), .A2(new_n550), .A3(new_n529), .ZN(new_n736));
  AND2_X1   g614(.A1(new_n552), .A2(new_n555), .ZN(new_n737));
  NAND4_X1  g615(.A1(new_n583), .A2(new_n735), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  AOI21_X1  g616(.A(new_n734), .B1(new_n738), .B2(new_n179), .ZN(new_n739));
  OAI211_X1 g617(.A(new_n731), .B(new_n733), .C1(new_n721), .C2(new_n739), .ZN(new_n740));
  NOR2_X1   g618(.A1(new_n739), .A2(new_n721), .ZN(new_n741));
  OAI21_X1  g619(.A(new_n732), .B1(new_n741), .B2(new_n730), .ZN(RLL_wire_A_125));
  XOR2_X1 RLL_XOR_125 (.A(RLL_wire_A_125), .B(KEYINPUT125), .Z(new_n742) );
  NAND2_X1  g620(.A1(new_n740), .A2(new_n742), .ZN(G72));
  NAND2_X1  g621(.A1(G472), .A2(G902), .ZN(new_n744));
  XNOR2_X1  g622(.A(new_n744), .B(KEYINPUT63), .ZN(new_n745));
  INV_X1    g623(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g624(.A(new_n746), .B1(new_n729), .B2(new_n713), .ZN(RLL_wire_A_126));
  XOR2_X1 RLL_XOR_126 (.A(RLL_wire_A_126), .B(KEYINPUT126), .Z(new_n747) );
  NAND2_X1  g625(.A1(new_n175), .A2(new_n177), .ZN(new_n748));
  NAND3_X1  g626(.A1(new_n747), .A2(new_n183), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g627(.A(new_n746), .B1(new_n738), .B2(new_n713), .ZN(RLL_wire_A_127));
  XOR2_X1 RLL_XOR_127 (.A(RLL_wire_A_127), .B(KEYINPUT127), .Z(new_n750) );
  NOR2_X1   g628(.A1(new_n748), .A2(new_n183), .ZN(new_n751));
  AOI21_X1  g629(.A(new_n676), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g630(.A(new_n202), .ZN(new_n753));
  AOI21_X1  g631(.A(new_n745), .B1(new_n753), .B2(new_n185), .ZN(new_n754));
  OAI21_X1  g632(.A(new_n754), .B1(new_n617), .B2(new_n620), .ZN(new_n755));
  AND3_X1   g633(.A1(new_n749), .A2(new_n752), .A3(new_n755), .ZN(G57));

endmodule
