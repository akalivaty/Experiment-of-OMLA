

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U548 ( .A1(n600), .A2(n599), .ZN(n997) );
  NAND2_X2 U549 ( .A1(G8), .A2(n649), .ZN(n682) );
  AND2_X1 U550 ( .A1(n514), .A2(n670), .ZN(n671) );
  NOR2_X1 U551 ( .A1(n644), .A2(n643), .ZN(n646) );
  NOR2_X1 U552 ( .A1(G543), .A2(n536), .ZN(n524) );
  XNOR2_X2 U553 ( .A(n519), .B(n518), .ZN(n584) );
  XOR2_X1 U554 ( .A(n631), .B(KEYINPUT29), .Z(n511) );
  XOR2_X1 U555 ( .A(KEYINPUT98), .B(n992), .Z(n512) );
  NOR2_X1 U556 ( .A1(n682), .A2(n681), .ZN(n513) );
  NOR2_X1 U557 ( .A1(n682), .A2(n590), .ZN(n514) );
  INV_X1 U558 ( .A(KEYINPUT26), .ZN(n601) );
  XNOR2_X1 U559 ( .A(n602), .B(n601), .ZN(n603) );
  NOR2_X1 U560 ( .A1(n619), .A2(n1000), .ZN(n613) );
  INV_X1 U561 ( .A(n649), .ZN(n614) );
  BUF_X1 U562 ( .A(n614), .Z(n633) );
  XNOR2_X1 U563 ( .A(KEYINPUT97), .B(KEYINPUT32), .ZN(n658) );
  XNOR2_X1 U564 ( .A(n659), .B(n658), .ZN(n667) );
  NAND2_X2 U565 ( .A1(n588), .A2(n687), .ZN(n649) );
  AND2_X1 U566 ( .A1(n736), .A2(G40), .ZN(n587) );
  NAND2_X1 U567 ( .A1(n737), .A2(n587), .ZN(n686) );
  XNOR2_X1 U568 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n519) );
  INV_X1 U569 ( .A(KEYINPUT23), .ZN(n580) );
  NOR2_X1 U570 ( .A1(G651), .A2(n537), .ZN(n767) );
  NOR2_X1 U571 ( .A1(n537), .A2(n536), .ZN(n774) );
  NAND2_X1 U572 ( .A1(n734), .A2(n733), .ZN(n735) );
  AND2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n873) );
  NAND2_X1 U574 ( .A1(G114), .A2(n873), .ZN(n516) );
  XOR2_X1 U575 ( .A(G2104), .B(KEYINPUT64), .Z(n517) );
  NOR2_X2 U576 ( .A1(n517), .A2(G2105), .ZN(n869) );
  NAND2_X1 U577 ( .A1(G102), .A2(n869), .ZN(n515) );
  NAND2_X1 U578 ( .A1(n516), .A2(n515), .ZN(n523) );
  AND2_X2 U579 ( .A1(n517), .A2(G2105), .ZN(n872) );
  NAND2_X1 U580 ( .A1(n872), .A2(G126), .ZN(n521) );
  NOR2_X1 U581 ( .A1(G2105), .A2(G2104), .ZN(n518) );
  NAND2_X1 U582 ( .A1(n584), .A2(G138), .ZN(n520) );
  NAND2_X1 U583 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U584 ( .A1(n523), .A2(n522), .ZN(G164) );
  INV_X1 U585 ( .A(G651), .ZN(n536) );
  XOR2_X1 U586 ( .A(KEYINPUT1), .B(n524), .Z(n766) );
  XOR2_X1 U587 ( .A(KEYINPUT0), .B(G543), .Z(n537) );
  NAND2_X1 U588 ( .A1(G49), .A2(n767), .ZN(n526) );
  NAND2_X1 U589 ( .A1(G74), .A2(G651), .ZN(n525) );
  NAND2_X1 U590 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U591 ( .A1(n766), .A2(n527), .ZN(n530) );
  NAND2_X1 U592 ( .A1(G87), .A2(n537), .ZN(n528) );
  XOR2_X1 U593 ( .A(KEYINPUT77), .B(n528), .Z(n529) );
  NAND2_X1 U594 ( .A1(n530), .A2(n529), .ZN(G288) );
  NAND2_X1 U595 ( .A1(G65), .A2(n766), .ZN(n532) );
  NOR2_X1 U596 ( .A1(G651), .A2(G543), .ZN(n770) );
  NAND2_X1 U597 ( .A1(G91), .A2(n770), .ZN(n531) );
  NAND2_X1 U598 ( .A1(n532), .A2(n531), .ZN(n535) );
  NAND2_X1 U599 ( .A1(G53), .A2(n767), .ZN(n533) );
  XNOR2_X1 U600 ( .A(KEYINPUT67), .B(n533), .ZN(n534) );
  NOR2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n539) );
  NAND2_X1 U602 ( .A1(n774), .A2(G78), .ZN(n538) );
  NAND2_X1 U603 ( .A1(n539), .A2(n538), .ZN(G299) );
  NAND2_X1 U604 ( .A1(n774), .A2(G77), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n540), .B(KEYINPUT66), .ZN(n542) );
  NAND2_X1 U606 ( .A1(G90), .A2(n770), .ZN(n541) );
  NAND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U608 ( .A(KEYINPUT9), .B(n543), .ZN(n547) );
  NAND2_X1 U609 ( .A1(G64), .A2(n766), .ZN(n545) );
  NAND2_X1 U610 ( .A1(G52), .A2(n767), .ZN(n544) );
  AND2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U612 ( .A1(n547), .A2(n546), .ZN(G301) );
  INV_X1 U613 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U614 ( .A(KEYINPUT72), .B(KEYINPUT6), .ZN(n551) );
  NAND2_X1 U615 ( .A1(G63), .A2(n766), .ZN(n549) );
  NAND2_X1 U616 ( .A1(G51), .A2(n767), .ZN(n548) );
  NAND2_X1 U617 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(n557) );
  NAND2_X1 U619 ( .A1(n770), .A2(G89), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n552), .B(KEYINPUT4), .ZN(n554) );
  NAND2_X1 U621 ( .A1(G76), .A2(n774), .ZN(n553) );
  NAND2_X1 U622 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U623 ( .A(KEYINPUT5), .B(n555), .Z(n556) );
  NOR2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n559) );
  XNOR2_X1 U625 ( .A(KEYINPUT7), .B(KEYINPUT73), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G88), .A2(n770), .ZN(n561) );
  NAND2_X1 U629 ( .A1(G75), .A2(n774), .ZN(n560) );
  NAND2_X1 U630 ( .A1(n561), .A2(n560), .ZN(n565) );
  NAND2_X1 U631 ( .A1(G62), .A2(n766), .ZN(n563) );
  NAND2_X1 U632 ( .A1(G50), .A2(n767), .ZN(n562) );
  NAND2_X1 U633 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U634 ( .A1(n565), .A2(n564), .ZN(G166) );
  INV_X1 U635 ( .A(G166), .ZN(G303) );
  NAND2_X1 U636 ( .A1(G61), .A2(n766), .ZN(n567) );
  NAND2_X1 U637 ( .A1(G86), .A2(n770), .ZN(n566) );
  NAND2_X1 U638 ( .A1(n567), .A2(n566), .ZN(n570) );
  NAND2_X1 U639 ( .A1(n774), .A2(G73), .ZN(n568) );
  XOR2_X1 U640 ( .A(KEYINPUT2), .B(n568), .Z(n569) );
  NOR2_X1 U641 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U642 ( .A(n571), .B(KEYINPUT78), .ZN(n573) );
  NAND2_X1 U643 ( .A1(G48), .A2(n767), .ZN(n572) );
  NAND2_X1 U644 ( .A1(n573), .A2(n572), .ZN(G305) );
  NAND2_X1 U645 ( .A1(G85), .A2(n770), .ZN(n575) );
  NAND2_X1 U646 ( .A1(G72), .A2(n774), .ZN(n574) );
  NAND2_X1 U647 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U648 ( .A1(G60), .A2(n766), .ZN(n577) );
  NAND2_X1 U649 ( .A1(G47), .A2(n767), .ZN(n576) );
  NAND2_X1 U650 ( .A1(n577), .A2(n576), .ZN(n578) );
  OR2_X1 U651 ( .A1(n579), .A2(n578), .ZN(G290) );
  NAND2_X1 U652 ( .A1(n869), .A2(G101), .ZN(n581) );
  XNOR2_X1 U653 ( .A(n581), .B(n580), .ZN(n583) );
  NAND2_X1 U654 ( .A1(n873), .A2(G113), .ZN(n582) );
  AND2_X1 U655 ( .A1(n583), .A2(n582), .ZN(n737) );
  NAND2_X1 U656 ( .A1(G137), .A2(n584), .ZN(n586) );
  NAND2_X1 U657 ( .A1(G125), .A2(n872), .ZN(n585) );
  AND2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n736) );
  INV_X1 U659 ( .A(n686), .ZN(n588) );
  NOR2_X1 U660 ( .A1(G164), .A2(G1384), .ZN(n687) );
  NOR2_X1 U661 ( .A1(G1976), .A2(G288), .ZN(n669) );
  NAND2_X1 U662 ( .A1(n669), .A2(KEYINPUT33), .ZN(n589) );
  NOR2_X1 U663 ( .A1(n682), .A2(n589), .ZN(n673) );
  NAND2_X1 U664 ( .A1(G1976), .A2(G288), .ZN(n986) );
  INV_X1 U665 ( .A(n986), .ZN(n590) );
  NAND2_X1 U666 ( .A1(n766), .A2(G56), .ZN(n591) );
  XNOR2_X1 U667 ( .A(n591), .B(KEYINPUT14), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n770), .A2(G81), .ZN(n592) );
  XNOR2_X1 U669 ( .A(n592), .B(KEYINPUT12), .ZN(n594) );
  NAND2_X1 U670 ( .A1(G68), .A2(n774), .ZN(n593) );
  NAND2_X1 U671 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U672 ( .A(KEYINPUT13), .B(n595), .ZN(n596) );
  NAND2_X1 U673 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U674 ( .A(n598), .B(KEYINPUT71), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n767), .A2(G43), .ZN(n599) );
  NAND2_X1 U676 ( .A1(G1996), .A2(n614), .ZN(n602) );
  NOR2_X1 U677 ( .A1(n997), .A2(n603), .ZN(n605) );
  NAND2_X1 U678 ( .A1(G1341), .A2(n649), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n619) );
  NAND2_X1 U680 ( .A1(G79), .A2(n774), .ZN(n607) );
  NAND2_X1 U681 ( .A1(G54), .A2(n767), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U683 ( .A1(G66), .A2(n766), .ZN(n609) );
  NAND2_X1 U684 ( .A1(G92), .A2(n770), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U686 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U687 ( .A(n612), .B(KEYINPUT15), .ZN(n1000) );
  XNOR2_X1 U688 ( .A(n613), .B(KEYINPUT93), .ZN(n618) );
  NOR2_X1 U689 ( .A1(n633), .A2(G1348), .ZN(n616) );
  NOR2_X1 U690 ( .A1(G2067), .A2(n649), .ZN(n615) );
  NOR2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U693 ( .A1(n619), .A2(n1000), .ZN(n620) );
  NAND2_X1 U694 ( .A1(n621), .A2(n620), .ZN(n626) );
  INV_X1 U695 ( .A(G299), .ZN(n987) );
  NAND2_X1 U696 ( .A1(n633), .A2(G2072), .ZN(n622) );
  XNOR2_X1 U697 ( .A(n622), .B(KEYINPUT27), .ZN(n624) );
  INV_X1 U698 ( .A(G1956), .ZN(n926) );
  NOR2_X1 U699 ( .A1(n926), .A2(n633), .ZN(n623) );
  NOR2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U701 ( .A1(n987), .A2(n627), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n626), .A2(n625), .ZN(n630) );
  NOR2_X1 U703 ( .A1(n987), .A2(n627), .ZN(n628) );
  XOR2_X1 U704 ( .A(n628), .B(KEYINPUT28), .Z(n629) );
  NAND2_X1 U705 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U706 ( .A1(n633), .A2(G1961), .ZN(n632) );
  XNOR2_X1 U707 ( .A(n632), .B(KEYINPUT91), .ZN(n635) );
  XNOR2_X1 U708 ( .A(KEYINPUT25), .B(G2078), .ZN(n903) );
  NAND2_X1 U709 ( .A1(n633), .A2(n903), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n642) );
  NAND2_X1 U711 ( .A1(G171), .A2(n642), .ZN(n636) );
  XNOR2_X1 U712 ( .A(KEYINPUT92), .B(n636), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n511), .A2(n637), .ZN(n648) );
  NOR2_X1 U714 ( .A1(G2084), .A2(n649), .ZN(n661) );
  NOR2_X1 U715 ( .A1(G1966), .A2(n682), .ZN(n638) );
  XOR2_X1 U716 ( .A(KEYINPUT90), .B(n638), .Z(n660) );
  NAND2_X1 U717 ( .A1(G8), .A2(n660), .ZN(n639) );
  NOR2_X1 U718 ( .A1(n661), .A2(n639), .ZN(n640) );
  XOR2_X1 U719 ( .A(KEYINPUT30), .B(n640), .Z(n641) );
  NOR2_X1 U720 ( .A1(G168), .A2(n641), .ZN(n644) );
  NOR2_X1 U721 ( .A1(G171), .A2(n642), .ZN(n643) );
  XOR2_X1 U722 ( .A(KEYINPUT94), .B(KEYINPUT31), .Z(n645) );
  XNOR2_X1 U723 ( .A(n646), .B(n645), .ZN(n647) );
  NAND2_X1 U724 ( .A1(n648), .A2(n647), .ZN(n663) );
  NAND2_X1 U725 ( .A1(n663), .A2(G286), .ZN(n655) );
  NOR2_X1 U726 ( .A1(G2090), .A2(n649), .ZN(n650) );
  XOR2_X1 U727 ( .A(KEYINPUT95), .B(n650), .Z(n652) );
  NOR2_X1 U728 ( .A1(G1971), .A2(n682), .ZN(n651) );
  NOR2_X1 U729 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U730 ( .A1(n653), .A2(G303), .ZN(n654) );
  NAND2_X1 U731 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U732 ( .A(n656), .B(KEYINPUT96), .ZN(n657) );
  NAND2_X1 U733 ( .A1(n657), .A2(G8), .ZN(n659) );
  INV_X1 U734 ( .A(n660), .ZN(n665) );
  NAND2_X1 U735 ( .A1(G8), .A2(n661), .ZN(n662) );
  NAND2_X1 U736 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U737 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X2 U738 ( .A1(n667), .A2(n666), .ZN(n677) );
  NOR2_X1 U739 ( .A1(G1971), .A2(G303), .ZN(n668) );
  NOR2_X1 U740 ( .A1(n669), .A2(n668), .ZN(n992) );
  OR2_X1 U741 ( .A1(n677), .A2(n512), .ZN(n670) );
  NOR2_X1 U742 ( .A1(KEYINPUT33), .A2(n671), .ZN(n672) );
  NOR2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U744 ( .A(G1981), .B(G305), .Z(n982) );
  NAND2_X1 U745 ( .A1(n674), .A2(n982), .ZN(n685) );
  NAND2_X1 U746 ( .A1(G166), .A2(G8), .ZN(n675) );
  NOR2_X1 U747 ( .A1(G2090), .A2(n675), .ZN(n676) );
  NOR2_X1 U748 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U749 ( .A(n678), .B(KEYINPUT99), .ZN(n679) );
  AND2_X1 U750 ( .A1(n679), .A2(n682), .ZN(n683) );
  NOR2_X1 U751 ( .A1(G1981), .A2(G305), .ZN(n680) );
  XOR2_X1 U752 ( .A(n680), .B(KEYINPUT24), .Z(n681) );
  NOR2_X1 U753 ( .A1(n683), .A2(n513), .ZN(n684) );
  AND2_X1 U754 ( .A1(n685), .A2(n684), .ZN(n699) );
  NOR2_X1 U755 ( .A1(n687), .A2(n686), .ZN(n731) );
  NAND2_X1 U756 ( .A1(G140), .A2(n584), .ZN(n689) );
  NAND2_X1 U757 ( .A1(G104), .A2(n869), .ZN(n688) );
  NAND2_X1 U758 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U759 ( .A(KEYINPUT34), .B(n690), .ZN(n696) );
  NAND2_X1 U760 ( .A1(G128), .A2(n872), .ZN(n692) );
  NAND2_X1 U761 ( .A1(G116), .A2(n873), .ZN(n691) );
  NAND2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U763 ( .A(KEYINPUT35), .B(n693), .Z(n694) );
  XNOR2_X1 U764 ( .A(KEYINPUT86), .B(n694), .ZN(n695) );
  NOR2_X1 U765 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U766 ( .A(KEYINPUT36), .B(n697), .ZN(n885) );
  XNOR2_X1 U767 ( .A(G2067), .B(KEYINPUT37), .ZN(n729) );
  NOR2_X1 U768 ( .A1(n885), .A2(n729), .ZN(n959) );
  NAND2_X1 U769 ( .A1(n731), .A2(n959), .ZN(n727) );
  INV_X1 U770 ( .A(n727), .ZN(n698) );
  NOR2_X1 U771 ( .A1(n699), .A2(n698), .ZN(n720) );
  NAND2_X1 U772 ( .A1(n872), .A2(G129), .ZN(n706) );
  NAND2_X1 U773 ( .A1(G141), .A2(n584), .ZN(n701) );
  NAND2_X1 U774 ( .A1(G117), .A2(n873), .ZN(n700) );
  NAND2_X1 U775 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U776 ( .A1(n869), .A2(G105), .ZN(n702) );
  XOR2_X1 U777 ( .A(KEYINPUT38), .B(n702), .Z(n703) );
  NOR2_X1 U778 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U779 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U780 ( .A(KEYINPUT87), .B(n707), .Z(n879) );
  NAND2_X1 U781 ( .A1(G1996), .A2(n879), .ZN(n708) );
  XNOR2_X1 U782 ( .A(n708), .B(KEYINPUT88), .ZN(n716) );
  NAND2_X1 U783 ( .A1(G131), .A2(n584), .ZN(n710) );
  NAND2_X1 U784 ( .A1(G107), .A2(n873), .ZN(n709) );
  NAND2_X1 U785 ( .A1(n710), .A2(n709), .ZN(n714) );
  NAND2_X1 U786 ( .A1(G119), .A2(n872), .ZN(n712) );
  NAND2_X1 U787 ( .A1(G95), .A2(n869), .ZN(n711) );
  NAND2_X1 U788 ( .A1(n712), .A2(n711), .ZN(n713) );
  OR2_X1 U789 ( .A1(n714), .A2(n713), .ZN(n855) );
  NAND2_X1 U790 ( .A1(G1991), .A2(n855), .ZN(n715) );
  NAND2_X1 U791 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U792 ( .A(KEYINPUT89), .B(n717), .ZN(n723) );
  XOR2_X1 U793 ( .A(G1986), .B(G290), .Z(n988) );
  NAND2_X1 U794 ( .A1(n723), .A2(n988), .ZN(n718) );
  NAND2_X1 U795 ( .A1(n718), .A2(n731), .ZN(n719) );
  NAND2_X1 U796 ( .A1(n720), .A2(n719), .ZN(n734) );
  NOR2_X1 U797 ( .A1(G1996), .A2(n879), .ZN(n948) );
  NOR2_X1 U798 ( .A1(G1991), .A2(n855), .ZN(n968) );
  NOR2_X1 U799 ( .A1(G1986), .A2(G290), .ZN(n721) );
  XNOR2_X1 U800 ( .A(KEYINPUT100), .B(n721), .ZN(n722) );
  NOR2_X1 U801 ( .A1(n968), .A2(n722), .ZN(n724) );
  INV_X1 U802 ( .A(n723), .ZN(n963) );
  NOR2_X1 U803 ( .A1(n724), .A2(n963), .ZN(n725) );
  NOR2_X1 U804 ( .A1(n948), .A2(n725), .ZN(n726) );
  XNOR2_X1 U805 ( .A(n726), .B(KEYINPUT39), .ZN(n728) );
  NAND2_X1 U806 ( .A1(n728), .A2(n727), .ZN(n730) );
  NAND2_X1 U807 ( .A1(n885), .A2(n729), .ZN(n966) );
  NAND2_X1 U808 ( .A1(n730), .A2(n966), .ZN(n732) );
  NAND2_X1 U809 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U810 ( .A(n735), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U811 ( .A1(n737), .A2(n736), .ZN(G160) );
  AND2_X1 U812 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U813 ( .A(G57), .ZN(G237) );
  INV_X1 U814 ( .A(G132), .ZN(G219) );
  INV_X1 U815 ( .A(G82), .ZN(G220) );
  NAND2_X1 U816 ( .A1(G7), .A2(G661), .ZN(n738) );
  XNOR2_X1 U817 ( .A(n738), .B(KEYINPUT68), .ZN(n739) );
  XNOR2_X1 U818 ( .A(KEYINPUT10), .B(n739), .ZN(G223) );
  XOR2_X1 U819 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n741) );
  INV_X1 U820 ( .A(G223), .ZN(n817) );
  NAND2_X1 U821 ( .A1(n817), .A2(G567), .ZN(n740) );
  XNOR2_X1 U822 ( .A(n741), .B(n740), .ZN(n742) );
  XOR2_X1 U823 ( .A(KEYINPUT69), .B(n742), .Z(G234) );
  INV_X1 U824 ( .A(G860), .ZN(n765) );
  OR2_X1 U825 ( .A1(n997), .A2(n765), .ZN(G153) );
  NAND2_X1 U826 ( .A1(G868), .A2(G301), .ZN(n744) );
  INV_X1 U827 ( .A(G868), .ZN(n788) );
  NAND2_X1 U828 ( .A1(n1000), .A2(n788), .ZN(n743) );
  NAND2_X1 U829 ( .A1(n744), .A2(n743), .ZN(G284) );
  NOR2_X1 U830 ( .A1(G286), .A2(n788), .ZN(n745) );
  XNOR2_X1 U831 ( .A(n745), .B(KEYINPUT74), .ZN(n747) );
  NOR2_X1 U832 ( .A1(G299), .A2(G868), .ZN(n746) );
  NOR2_X1 U833 ( .A1(n747), .A2(n746), .ZN(G297) );
  NAND2_X1 U834 ( .A1(G559), .A2(n765), .ZN(n748) );
  XOR2_X1 U835 ( .A(KEYINPUT75), .B(n748), .Z(n749) );
  INV_X1 U836 ( .A(n1000), .ZN(n763) );
  NAND2_X1 U837 ( .A1(n749), .A2(n763), .ZN(n750) );
  XNOR2_X1 U838 ( .A(n750), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U839 ( .A1(G868), .A2(n997), .ZN(n753) );
  NAND2_X1 U840 ( .A1(n763), .A2(G868), .ZN(n751) );
  NOR2_X1 U841 ( .A1(G559), .A2(n751), .ZN(n752) );
  NOR2_X1 U842 ( .A1(n753), .A2(n752), .ZN(G282) );
  NAND2_X1 U843 ( .A1(G135), .A2(n584), .ZN(n755) );
  NAND2_X1 U844 ( .A1(G111), .A2(n873), .ZN(n754) );
  NAND2_X1 U845 ( .A1(n755), .A2(n754), .ZN(n760) );
  NAND2_X1 U846 ( .A1(n872), .A2(G123), .ZN(n756) );
  XNOR2_X1 U847 ( .A(n756), .B(KEYINPUT18), .ZN(n758) );
  NAND2_X1 U848 ( .A1(G99), .A2(n869), .ZN(n757) );
  NAND2_X1 U849 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U850 ( .A1(n760), .A2(n759), .ZN(n965) );
  XNOR2_X1 U851 ( .A(n965), .B(G2096), .ZN(n762) );
  INV_X1 U852 ( .A(G2100), .ZN(n761) );
  NAND2_X1 U853 ( .A1(n762), .A2(n761), .ZN(G156) );
  NAND2_X1 U854 ( .A1(G559), .A2(n763), .ZN(n764) );
  XOR2_X1 U855 ( .A(n997), .B(n764), .Z(n785) );
  NAND2_X1 U856 ( .A1(n765), .A2(n785), .ZN(n777) );
  NAND2_X1 U857 ( .A1(G67), .A2(n766), .ZN(n769) );
  NAND2_X1 U858 ( .A1(G55), .A2(n767), .ZN(n768) );
  NAND2_X1 U859 ( .A1(n769), .A2(n768), .ZN(n773) );
  NAND2_X1 U860 ( .A1(n770), .A2(G93), .ZN(n771) );
  XOR2_X1 U861 ( .A(KEYINPUT76), .B(n771), .Z(n772) );
  NOR2_X1 U862 ( .A1(n773), .A2(n772), .ZN(n776) );
  NAND2_X1 U863 ( .A1(n774), .A2(G80), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n789) );
  XNOR2_X1 U865 ( .A(n777), .B(n789), .ZN(G145) );
  XNOR2_X1 U866 ( .A(KEYINPUT80), .B(KEYINPUT19), .ZN(n779) );
  XNOR2_X1 U867 ( .A(G288), .B(KEYINPUT79), .ZN(n778) );
  XNOR2_X1 U868 ( .A(n779), .B(n778), .ZN(n782) );
  XNOR2_X1 U869 ( .A(n987), .B(G305), .ZN(n780) );
  XNOR2_X1 U870 ( .A(n780), .B(n789), .ZN(n781) );
  XNOR2_X1 U871 ( .A(n782), .B(n781), .ZN(n784) );
  XNOR2_X1 U872 ( .A(G290), .B(G166), .ZN(n783) );
  XNOR2_X1 U873 ( .A(n784), .B(n783), .ZN(n890) );
  XNOR2_X1 U874 ( .A(n785), .B(n890), .ZN(n786) );
  XNOR2_X1 U875 ( .A(KEYINPUT81), .B(n786), .ZN(n787) );
  NOR2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n791) );
  NOR2_X1 U877 ( .A1(G868), .A2(n789), .ZN(n790) );
  NOR2_X1 U878 ( .A1(n791), .A2(n790), .ZN(G295) );
  NAND2_X1 U879 ( .A1(G2084), .A2(G2078), .ZN(n792) );
  XOR2_X1 U880 ( .A(KEYINPUT20), .B(n792), .Z(n793) );
  NAND2_X1 U881 ( .A1(G2090), .A2(n793), .ZN(n794) );
  XNOR2_X1 U882 ( .A(n794), .B(KEYINPUT83), .ZN(n796) );
  XOR2_X1 U883 ( .A(KEYINPUT21), .B(KEYINPUT82), .Z(n795) );
  XNOR2_X1 U884 ( .A(n796), .B(n795), .ZN(n797) );
  NAND2_X1 U885 ( .A1(n797), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U886 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U887 ( .A1(G220), .A2(G219), .ZN(n798) );
  XOR2_X1 U888 ( .A(KEYINPUT22), .B(n798), .Z(n799) );
  NOR2_X1 U889 ( .A1(G218), .A2(n799), .ZN(n800) );
  NAND2_X1 U890 ( .A1(G96), .A2(n800), .ZN(n822) );
  NAND2_X1 U891 ( .A1(n822), .A2(G2106), .ZN(n804) );
  NAND2_X1 U892 ( .A1(G120), .A2(G108), .ZN(n801) );
  NOR2_X1 U893 ( .A1(G237), .A2(n801), .ZN(n802) );
  NAND2_X1 U894 ( .A1(G69), .A2(n802), .ZN(n823) );
  NAND2_X1 U895 ( .A1(n823), .A2(G567), .ZN(n803) );
  NAND2_X1 U896 ( .A1(n804), .A2(n803), .ZN(n824) );
  NAND2_X1 U897 ( .A1(G661), .A2(G483), .ZN(n805) );
  XNOR2_X1 U898 ( .A(KEYINPUT84), .B(n805), .ZN(n806) );
  NOR2_X1 U899 ( .A1(n824), .A2(n806), .ZN(n821) );
  NAND2_X1 U900 ( .A1(n821), .A2(G36), .ZN(n807) );
  XOR2_X1 U901 ( .A(KEYINPUT85), .B(n807), .Z(G176) );
  XNOR2_X1 U902 ( .A(G1348), .B(G2454), .ZN(n808) );
  XNOR2_X1 U903 ( .A(n808), .B(G2430), .ZN(n809) );
  XNOR2_X1 U904 ( .A(n809), .B(G1341), .ZN(n815) );
  XOR2_X1 U905 ( .A(G2443), .B(G2427), .Z(n811) );
  XNOR2_X1 U906 ( .A(G2438), .B(G2446), .ZN(n810) );
  XNOR2_X1 U907 ( .A(n811), .B(n810), .ZN(n813) );
  XOR2_X1 U908 ( .A(G2451), .B(G2435), .Z(n812) );
  XNOR2_X1 U909 ( .A(n813), .B(n812), .ZN(n814) );
  XNOR2_X1 U910 ( .A(n815), .B(n814), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n816), .A2(G14), .ZN(n894) );
  XNOR2_X1 U912 ( .A(KEYINPUT101), .B(n894), .ZN(G401) );
  NAND2_X1 U913 ( .A1(n817), .A2(G2106), .ZN(n818) );
  XNOR2_X1 U914 ( .A(n818), .B(KEYINPUT102), .ZN(G217) );
  AND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n819) );
  NAND2_X1 U916 ( .A1(G661), .A2(n819), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n820) );
  NAND2_X1 U918 ( .A1(n821), .A2(n820), .ZN(G188) );
  XNOR2_X1 U919 ( .A(G96), .B(KEYINPUT103), .ZN(G221) );
  NOR2_X1 U920 ( .A1(n823), .A2(n822), .ZN(G325) );
  XOR2_X1 U921 ( .A(KEYINPUT104), .B(G325), .Z(G261) );
  XOR2_X1 U922 ( .A(G108), .B(KEYINPUT114), .Z(G238) );
  INV_X1 U924 ( .A(G120), .ZN(G236) );
  INV_X1 U925 ( .A(n824), .ZN(G319) );
  XOR2_X1 U926 ( .A(G2474), .B(G1981), .Z(n826) );
  XNOR2_X1 U927 ( .A(G1996), .B(G1991), .ZN(n825) );
  XNOR2_X1 U928 ( .A(n826), .B(n825), .ZN(n827) );
  XOR2_X1 U929 ( .A(n827), .B(KEYINPUT107), .Z(n829) );
  XNOR2_X1 U930 ( .A(G1956), .B(G1976), .ZN(n828) );
  XNOR2_X1 U931 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U932 ( .A(G1971), .B(G1961), .Z(n831) );
  XNOR2_X1 U933 ( .A(G1986), .B(G1966), .ZN(n830) );
  XNOR2_X1 U934 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U935 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U936 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n834) );
  XNOR2_X1 U937 ( .A(n835), .B(n834), .ZN(G229) );
  XOR2_X1 U938 ( .A(G2678), .B(KEYINPUT43), .Z(n837) );
  XNOR2_X1 U939 ( .A(KEYINPUT106), .B(KEYINPUT105), .ZN(n836) );
  XNOR2_X1 U940 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U941 ( .A(KEYINPUT42), .B(G2090), .Z(n839) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2072), .ZN(n838) );
  XNOR2_X1 U943 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U944 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U945 ( .A(G2096), .B(G2100), .ZN(n842) );
  XNOR2_X1 U946 ( .A(n843), .B(n842), .ZN(n845) );
  XOR2_X1 U947 ( .A(G2084), .B(G2078), .Z(n844) );
  XNOR2_X1 U948 ( .A(n845), .B(n844), .ZN(G227) );
  NAND2_X1 U949 ( .A1(G100), .A2(n869), .ZN(n852) );
  NAND2_X1 U950 ( .A1(G136), .A2(n584), .ZN(n847) );
  NAND2_X1 U951 ( .A1(G112), .A2(n873), .ZN(n846) );
  NAND2_X1 U952 ( .A1(n847), .A2(n846), .ZN(n850) );
  NAND2_X1 U953 ( .A1(n872), .A2(G124), .ZN(n848) );
  XOR2_X1 U954 ( .A(KEYINPUT44), .B(n848), .Z(n849) );
  NOR2_X1 U955 ( .A1(n850), .A2(n849), .ZN(n851) );
  NAND2_X1 U956 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U957 ( .A(n853), .B(KEYINPUT109), .ZN(G162) );
  XOR2_X1 U958 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n854) );
  XNOR2_X1 U959 ( .A(n855), .B(n854), .ZN(n868) );
  NAND2_X1 U960 ( .A1(n873), .A2(G118), .ZN(n856) );
  XNOR2_X1 U961 ( .A(KEYINPUT111), .B(n856), .ZN(n859) );
  NAND2_X1 U962 ( .A1(n872), .A2(G130), .ZN(n857) );
  XOR2_X1 U963 ( .A(KEYINPUT110), .B(n857), .Z(n858) );
  NOR2_X1 U964 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U965 ( .A(n860), .B(KEYINPUT112), .ZN(n865) );
  NAND2_X1 U966 ( .A1(G142), .A2(n584), .ZN(n862) );
  NAND2_X1 U967 ( .A1(G106), .A2(n869), .ZN(n861) );
  NAND2_X1 U968 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U969 ( .A(KEYINPUT45), .B(n863), .ZN(n864) );
  NAND2_X1 U970 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U971 ( .A(n866), .B(n965), .ZN(n867) );
  XNOR2_X1 U972 ( .A(n868), .B(n867), .ZN(n881) );
  NAND2_X1 U973 ( .A1(G139), .A2(n584), .ZN(n871) );
  NAND2_X1 U974 ( .A1(G103), .A2(n869), .ZN(n870) );
  NAND2_X1 U975 ( .A1(n871), .A2(n870), .ZN(n878) );
  NAND2_X1 U976 ( .A1(G127), .A2(n872), .ZN(n875) );
  NAND2_X1 U977 ( .A1(G115), .A2(n873), .ZN(n874) );
  NAND2_X1 U978 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n876), .Z(n877) );
  NOR2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n951) );
  XNOR2_X1 U981 ( .A(n879), .B(n951), .ZN(n880) );
  XNOR2_X1 U982 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U983 ( .A(n882), .B(G162), .Z(n884) );
  XNOR2_X1 U984 ( .A(G164), .B(G160), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n884), .B(n883), .ZN(n886) );
  XOR2_X1 U986 ( .A(n886), .B(n885), .Z(n887) );
  NOR2_X1 U987 ( .A1(G37), .A2(n887), .ZN(G395) );
  XNOR2_X1 U988 ( .A(KEYINPUT113), .B(G301), .ZN(n888) );
  XNOR2_X1 U989 ( .A(n888), .B(n1000), .ZN(n889) );
  XNOR2_X1 U990 ( .A(n890), .B(n889), .ZN(n892) );
  XNOR2_X1 U991 ( .A(n997), .B(G286), .ZN(n891) );
  XNOR2_X1 U992 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U993 ( .A1(G37), .A2(n893), .ZN(G397) );
  NAND2_X1 U994 ( .A1(G319), .A2(n894), .ZN(n897) );
  NOR2_X1 U995 ( .A1(G229), .A2(G227), .ZN(n895) );
  XNOR2_X1 U996 ( .A(KEYINPUT49), .B(n895), .ZN(n896) );
  NOR2_X1 U997 ( .A1(n897), .A2(n896), .ZN(n899) );
  NOR2_X1 U998 ( .A1(G395), .A2(G397), .ZN(n898) );
  NAND2_X1 U999 ( .A1(n899), .A2(n898), .ZN(G225) );
  INV_X1 U1000 ( .A(G225), .ZN(G308) );
  INV_X1 U1001 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1002 ( .A(KEYINPUT121), .B(G29), .ZN(n919) );
  XNOR2_X1 U1003 ( .A(G2067), .B(G26), .ZN(n901) );
  XNOR2_X1 U1004 ( .A(G33), .B(G2072), .ZN(n900) );
  NOR2_X1 U1005 ( .A1(n901), .A2(n900), .ZN(n908) );
  XOR2_X1 U1006 ( .A(G1996), .B(G32), .Z(n902) );
  NAND2_X1 U1007 ( .A1(n902), .A2(G28), .ZN(n906) );
  XOR2_X1 U1008 ( .A(G27), .B(n903), .Z(n904) );
  XNOR2_X1 U1009 ( .A(KEYINPUT120), .B(n904), .ZN(n905) );
  NOR2_X1 U1010 ( .A1(n906), .A2(n905), .ZN(n907) );
  NAND2_X1 U1011 ( .A1(n908), .A2(n907), .ZN(n910) );
  XNOR2_X1 U1012 ( .A(G25), .B(G1991), .ZN(n909) );
  NOR2_X1 U1013 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1014 ( .A(KEYINPUT53), .B(n911), .Z(n914) );
  XOR2_X1 U1015 ( .A(KEYINPUT54), .B(G34), .Z(n912) );
  XNOR2_X1 U1016 ( .A(G2084), .B(n912), .ZN(n913) );
  NAND2_X1 U1017 ( .A1(n914), .A2(n913), .ZN(n916) );
  XNOR2_X1 U1018 ( .A(G35), .B(G2090), .ZN(n915) );
  NOR2_X1 U1019 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1020 ( .A(KEYINPUT55), .B(n917), .ZN(n918) );
  NAND2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1022 ( .A(KEYINPUT122), .B(n920), .ZN(n980) );
  XNOR2_X1 U1023 ( .A(G1348), .B(KEYINPUT59), .ZN(n921) );
  XNOR2_X1 U1024 ( .A(n921), .B(G4), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(G1341), .B(G19), .ZN(n923) );
  XNOR2_X1 U1026 ( .A(G1981), .B(G6), .ZN(n922) );
  NOR2_X1 U1027 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1028 ( .A1(n925), .A2(n924), .ZN(n929) );
  XOR2_X1 U1029 ( .A(G20), .B(n926), .Z(n927) );
  XNOR2_X1 U1030 ( .A(KEYINPUT126), .B(n927), .ZN(n928) );
  NOR2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1032 ( .A(KEYINPUT60), .B(n930), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(G1966), .B(G21), .ZN(n932) );
  XNOR2_X1 U1034 ( .A(G1961), .B(G5), .ZN(n931) );
  NOR2_X1 U1035 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1036 ( .A1(n934), .A2(n933), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(G1986), .B(G24), .ZN(n936) );
  XNOR2_X1 U1038 ( .A(G22), .B(G1971), .ZN(n935) );
  NOR2_X1 U1039 ( .A1(n936), .A2(n935), .ZN(n939) );
  XNOR2_X1 U1040 ( .A(G1976), .B(KEYINPUT127), .ZN(n937) );
  XNOR2_X1 U1041 ( .A(n937), .B(G23), .ZN(n938) );
  NAND2_X1 U1042 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1043 ( .A(KEYINPUT58), .B(n940), .ZN(n941) );
  NOR2_X1 U1044 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1045 ( .A(KEYINPUT61), .B(n943), .ZN(n945) );
  INV_X1 U1046 ( .A(G16), .ZN(n944) );
  NAND2_X1 U1047 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1048 ( .A1(n946), .A2(G11), .ZN(n978) );
  XOR2_X1 U1049 ( .A(G2090), .B(G162), .Z(n947) );
  NOR2_X1 U1050 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1051 ( .A(KEYINPUT115), .B(n949), .ZN(n950) );
  XNOR2_X1 U1052 ( .A(n950), .B(KEYINPUT51), .ZN(n961) );
  XOR2_X1 U1053 ( .A(G2072), .B(n951), .Z(n952) );
  XNOR2_X1 U1054 ( .A(KEYINPUT116), .B(n952), .ZN(n955) );
  XNOR2_X1 U1055 ( .A(G2078), .B(G164), .ZN(n953) );
  XNOR2_X1 U1056 ( .A(KEYINPUT117), .B(n953), .ZN(n954) );
  NOR2_X1 U1057 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1058 ( .A(n956), .B(KEYINPUT118), .Z(n957) );
  XNOR2_X1 U1059 ( .A(KEYINPUT50), .B(n957), .ZN(n958) );
  NOR2_X1 U1060 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1061 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1062 ( .A1(n963), .A2(n962), .ZN(n971) );
  XOR2_X1 U1063 ( .A(G2084), .B(G160), .Z(n964) );
  NOR2_X1 U1064 ( .A1(n965), .A2(n964), .ZN(n967) );
  NAND2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n969) );
  NOR2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1068 ( .A(KEYINPUT52), .B(n972), .ZN(n973) );
  XOR2_X1 U1069 ( .A(KEYINPUT119), .B(n973), .Z(n974) );
  NOR2_X1 U1070 ( .A1(KEYINPUT55), .A2(n974), .ZN(n976) );
  INV_X1 U1071 ( .A(G29), .ZN(n975) );
  NOR2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n1009) );
  XNOR2_X1 U1075 ( .A(G16), .B(KEYINPUT56), .ZN(n1006) );
  XOR2_X1 U1076 ( .A(G1966), .B(G168), .Z(n981) );
  XNOR2_X1 U1077 ( .A(KEYINPUT123), .B(n981), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1079 ( .A(n984), .B(KEYINPUT57), .ZN(n996) );
  NAND2_X1 U1080 ( .A1(G1971), .A2(G303), .ZN(n985) );
  NAND2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(n987), .B(G1956), .ZN(n989) );
  NAND2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1086 ( .A(KEYINPUT124), .B(n994), .Z(n995) );
  NAND2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(G1341), .B(n997), .ZN(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1004) );
  XNOR2_X1 U1090 ( .A(G301), .B(G1961), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(n1000), .B(G1348), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(KEYINPUT125), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(n1010), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1098 ( .A(G311), .ZN(G150) );
endmodule

