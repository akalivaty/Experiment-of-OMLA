//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011, new_n1012;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT88), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(G8gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  AOI21_X1  g005(.A(G1gat), .B1(new_n202), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n205), .B(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n210));
  NAND2_X1  g009(.A1(G29gat), .A2(G36gat), .ZN(new_n211));
  XOR2_X1   g010(.A(new_n211), .B(KEYINPUT84), .Z(new_n212));
  NOR2_X1   g011(.A1(G29gat), .A2(G36gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(KEYINPUT14), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT85), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n209), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218));
  INV_X1    g017(.A(G50gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G43gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n217), .B(new_n218), .C1(new_n216), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n215), .B1(new_n221), .B2(KEYINPUT86), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n218), .B1(new_n220), .B2(new_n216), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n223), .B1(new_n216), .B2(new_n209), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT86), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n210), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  NOR3_X1   g026(.A1(new_n212), .A2(new_n214), .A3(new_n210), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n208), .B1(new_n230), .B2(KEYINPUT17), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT87), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n221), .A2(KEYINPUT86), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n224), .A2(new_n225), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n234), .A3(new_n215), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n228), .B1(new_n235), .B2(new_n210), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT17), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n232), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AND4_X1   g037(.A1(new_n232), .A2(new_n227), .A3(new_n237), .A4(new_n229), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n231), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n208), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n241), .A2(new_n230), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G229gat), .A2(G233gat), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n240), .A2(KEYINPUT18), .A3(new_n243), .A4(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n236), .B(new_n208), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n244), .B(KEYINPUT13), .Z(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT87), .B1(new_n230), .B2(KEYINPUT17), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n236), .A2(new_n232), .A3(new_n237), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n242), .B1(new_n252), .B2(new_n231), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n244), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT18), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT89), .ZN(new_n257));
  XNOR2_X1  g056(.A(G113gat), .B(G141gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(G197gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT11), .B(G169gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT12), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n249), .B(new_n256), .C1(new_n257), .C2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n245), .A2(new_n257), .A3(new_n248), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT18), .B1(new_n253), .B2(new_n244), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n245), .A2(new_n248), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n265), .B(new_n262), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G228gat), .A2(G233gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(G211gat), .B(G218gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G218gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT70), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G218gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT22), .B1(new_n278), .B2(G211gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(G197gat), .B(G204gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n273), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G211gat), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n283), .B1(new_n275), .B2(new_n277), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n280), .B(new_n272), .C1(new_n284), .C2(KEYINPUT22), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  AND2_X1   g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(G155gat), .A2(G162gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G141gat), .B(G148gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT2), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n291), .B1(G155gat), .B2(G162gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n289), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G141gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G148gat), .ZN(new_n295));
  INV_X1    g094(.A(G148gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G141gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G155gat), .B(G162gat), .ZN(new_n299));
  INV_X1    g098(.A(G155gat), .ZN(new_n300));
  INV_X1    g099(.A(G162gat), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT2), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n298), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT3), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n293), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT73), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n293), .A2(new_n303), .A3(KEYINPUT73), .A4(new_n304), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT29), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n286), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n293), .A2(new_n303), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n285), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT22), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT70), .B(G218gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n315), .B1(new_n316), .B2(new_n283), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n272), .B1(new_n317), .B2(new_n280), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n310), .B1(new_n314), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n313), .B1(new_n319), .B2(new_n304), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n271), .B1(new_n311), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G22gat), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n293), .A2(new_n303), .A3(KEYINPUT72), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT72), .B1(new_n293), .B2(new_n303), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT29), .B1(new_n282), .B2(new_n285), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n325), .B1(new_n326), .B2(KEYINPUT3), .ZN(new_n327));
  INV_X1    g126(.A(new_n271), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT29), .B1(new_n307), .B2(new_n308), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n327), .B(new_n328), .C1(new_n286), .C2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n321), .A2(new_n322), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT79), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n321), .A2(new_n330), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(G22gat), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n321), .A2(new_n330), .A3(KEYINPUT79), .A4(new_n322), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G78gat), .B(G106gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT31), .B(G50gat), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n338), .B(new_n339), .Z(new_n340));
  XOR2_X1   g139(.A(new_n340), .B(KEYINPUT78), .Z(new_n341));
  NAND2_X1  g140(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n340), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n335), .A2(new_n331), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G120gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G113gat), .ZN(new_n348));
  INV_X1    g147(.A(G113gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G120gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT1), .ZN(new_n352));
  INV_X1    g151(.A(G134gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G127gat), .ZN(new_n354));
  INV_X1    g153(.A(G127gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G134gat), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n351), .A2(new_n352), .A3(new_n354), .A4(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n356), .ZN(new_n358));
  XNOR2_X1  g157(.A(G113gat), .B(G120gat), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n358), .B1(new_n359), .B2(KEYINPUT1), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT66), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT65), .B(KEYINPUT24), .ZN(new_n363));
  NAND2_X1  g162(.A1(G183gat), .A2(G190gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n362), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G183gat), .ZN(new_n367));
  INV_X1    g166(.A(G190gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT65), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n373), .A2(KEYINPUT24), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT24), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n375), .A2(KEYINPUT65), .ZN(new_n376));
  OAI211_X1 g175(.A(KEYINPUT66), .B(new_n364), .C1(new_n374), .C2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n366), .A2(new_n372), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT23), .ZN(new_n379));
  INV_X1    g178(.A(G169gat), .ZN(new_n380));
  INV_X1    g179(.A(G176gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(G169gat), .A2(G176gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT64), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT64), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(G169gat), .A3(G176gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(new_n389), .A3(KEYINPUT25), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n369), .B(new_n370), .C1(new_n365), .C2(KEYINPUT24), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n392), .A2(new_n389), .A3(new_n384), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT25), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n378), .A2(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n367), .A2(KEYINPUT27), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT27), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G183gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n398), .A3(new_n368), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT67), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n400), .A3(KEYINPUT28), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n402));
  OR3_X1    g201(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n389), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n401), .A2(new_n404), .A3(new_n364), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT28), .B1(new_n399), .B2(new_n400), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n361), .B1(new_n395), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n399), .A2(new_n400), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT28), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n411), .A2(new_n364), .A3(new_n401), .A4(new_n404), .ZN(new_n412));
  INV_X1    g211(.A(new_n361), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n364), .B1(new_n374), .B2(new_n376), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n371), .B1(new_n414), .B2(new_n362), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n390), .B1(new_n415), .B2(new_n377), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n393), .A2(new_n394), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n412), .B(new_n413), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n408), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G227gat), .A2(G233gat), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT32), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT33), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  XOR2_X1   g224(.A(G15gat), .B(G43gat), .Z(new_n426));
  XNOR2_X1  g225(.A(G71gat), .B(G99gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n423), .A2(new_n425), .A3(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT34), .B1(new_n419), .B2(new_n421), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT34), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n408), .A2(new_n431), .A3(new_n418), .A4(new_n420), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT68), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n420), .B1(new_n408), .B2(new_n418), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n428), .B1(new_n436), .B2(KEYINPUT33), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT32), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n432), .A2(new_n433), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n429), .A2(new_n435), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n430), .A3(new_n434), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n437), .A2(new_n439), .ZN(new_n444));
  AOI221_X4 g243(.A(new_n438), .B1(KEYINPUT33), .B2(new_n428), .C1(new_n419), .C2(new_n421), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT82), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n442), .A2(new_n446), .A3(KEYINPUT82), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n346), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT35), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT72), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n312), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n293), .A2(new_n303), .A3(KEYINPUT72), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(KEYINPUT3), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n309), .A2(new_n455), .A3(new_n361), .ZN(new_n456));
  NAND2_X1  g255(.A1(G225gat), .A2(G233gat), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n293), .A2(new_n357), .A3(new_n360), .A4(new_n303), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(KEYINPUT4), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n456), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT75), .ZN(new_n461));
  XNOR2_X1  g260(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n462));
  INV_X1    g261(.A(new_n458), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n463), .B1(new_n325), .B2(new_n361), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n462), .B1(new_n464), .B2(new_n457), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  XOR2_X1   g266(.A(G1gat), .B(G29gat), .Z(new_n468));
  XNOR2_X1  g267(.A(G57gat), .B(G85gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n470), .B(new_n471), .Z(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n465), .A2(new_n460), .A3(KEYINPUT75), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n467), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(KEYINPUT77), .B(KEYINPUT6), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n465), .A2(new_n460), .A3(KEYINPUT75), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n465), .B1(KEYINPUT75), .B2(new_n460), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n476), .B1(new_n481), .B2(new_n473), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n472), .B1(new_n479), .B2(new_n480), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n478), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n286), .ZN(new_n485));
  INV_X1    g284(.A(G226gat), .ZN(new_n486));
  INV_X1    g285(.A(G233gat), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n412), .B1(new_n416), .B2(new_n417), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n488), .B1(new_n489), .B2(new_n310), .ZN(new_n490));
  INV_X1    g289(.A(new_n488), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n378), .A2(new_n391), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n393), .A2(new_n394), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n491), .B1(new_n494), .B2(new_n412), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n485), .B1(new_n490), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G8gat), .B(G36gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(G64gat), .B(G92gat), .ZN(new_n498));
  XOR2_X1   g297(.A(new_n497), .B(new_n498), .Z(new_n499));
  NAND2_X1  g298(.A1(new_n489), .A2(new_n488), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT29), .B1(new_n494), .B2(new_n412), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n500), .B(new_n286), .C1(new_n501), .C2(new_n488), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n496), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT71), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT30), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n496), .A2(new_n502), .A3(KEYINPUT71), .A4(new_n499), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n499), .B1(new_n496), .B2(new_n502), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n496), .A2(new_n499), .A3(new_n502), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n509), .B1(new_n510), .B2(KEYINPUT30), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n484), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n450), .A2(KEYINPUT83), .A3(new_n451), .A4(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT69), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n442), .A2(new_n446), .A3(new_n515), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n443), .B(KEYINPUT69), .C1(new_n444), .C2(new_n445), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n345), .ZN(new_n519));
  INV_X1    g318(.A(new_n512), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n483), .A2(new_n475), .A3(new_n477), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n481), .A2(new_n473), .A3(new_n476), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT35), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT83), .ZN(new_n526));
  INV_X1    g325(.A(new_n449), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n345), .B1(new_n527), .B2(new_n447), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n520), .A2(new_n523), .A3(new_n451), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n525), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT36), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n532), .B1(new_n516), .B2(new_n517), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT36), .B1(new_n442), .B2(new_n446), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n534), .A2(new_n536), .B1(new_n346), .B2(new_n524), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT40), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n456), .A2(new_n459), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT39), .ZN(new_n540));
  INV_X1    g339(.A(new_n457), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n472), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n453), .A2(new_n361), .A3(new_n454), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n458), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT39), .B1(new_n545), .B2(new_n541), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n546), .B1(new_n541), .B2(new_n539), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n538), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n539), .A2(new_n541), .ZN(new_n549));
  INV_X1    g348(.A(new_n546), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n551), .A2(KEYINPUT40), .A3(new_n472), .A4(new_n542), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n548), .A2(new_n475), .A3(new_n552), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n512), .A2(new_n553), .B1(new_n342), .B2(new_n344), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT81), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT80), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT37), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n496), .A2(new_n557), .A3(new_n502), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n496), .B2(new_n502), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n558), .A2(new_n559), .A3(new_n499), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT38), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n556), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n559), .ZN(new_n563));
  INV_X1    g362(.A(new_n499), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n496), .A2(new_n557), .A3(new_n502), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n566), .A2(KEYINPUT80), .A3(KEYINPUT38), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n505), .A2(new_n507), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n563), .A2(new_n561), .A3(new_n564), .A4(new_n565), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n570), .A2(new_n521), .A3(new_n522), .A4(new_n571), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n554), .B(new_n555), .C1(new_n568), .C2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n569), .B1(new_n560), .B2(new_n561), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n484), .A2(new_n575), .A3(new_n562), .A4(new_n567), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n555), .B1(new_n576), .B2(new_n554), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n537), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n270), .B1(new_n531), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT99), .ZN(new_n580));
  NAND2_X1  g379(.A1(G230gat), .A2(G233gat), .ZN(new_n581));
  XOR2_X1   g380(.A(G99gat), .B(G106gat), .Z(new_n582));
  NAND2_X1  g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583));
  INV_X1    g382(.A(G85gat), .ZN(new_n584));
  INV_X1    g383(.A(G92gat), .ZN(new_n585));
  AOI22_X1  g384(.A1(KEYINPUT8), .A2(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT97), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT96), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(G85gat), .A3(G92gat), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n589), .B(KEYINPUT7), .Z(new_n590));
  OAI21_X1  g389(.A(new_n582), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT97), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n586), .B(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n582), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n589), .B(KEYINPUT7), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G57gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(G64gat), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n599), .A2(KEYINPUT92), .ZN(new_n600));
  INV_X1    g399(.A(G64gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(G57gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n599), .A2(KEYINPUT92), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(G71gat), .ZN(new_n605));
  INV_X1    g404(.A(G78gat), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(new_n606), .A3(KEYINPUT9), .ZN(new_n607));
  NAND2_X1  g406(.A1(G71gat), .A2(G78gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n599), .A2(new_n602), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT9), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n611), .A2(new_n613), .B1(new_n605), .B2(new_n606), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT91), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n608), .B(KEYINPUT90), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n615), .B1(new_n614), .B2(new_n616), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n610), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT98), .B1(new_n597), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n614), .A2(new_n616), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT91), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n622), .A2(new_n623), .B1(new_n609), .B2(new_n604), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(new_n596), .A3(new_n591), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n597), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n627), .A2(KEYINPUT98), .A3(new_n624), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT10), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT10), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n581), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n581), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n626), .A2(new_n628), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(G176gat), .B(G204gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n580), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n632), .A2(new_n634), .A3(KEYINPUT99), .A4(new_n638), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n635), .A2(new_n639), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n645));
  NOR2_X1   g444(.A1(new_n624), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(G127gat), .B(G155gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n208), .B1(KEYINPUT21), .B2(new_n624), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n648), .B(new_n649), .Z(new_n650));
  NAND2_X1  g449(.A1(G231gat), .A2(G233gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT94), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G183gat), .B(G211gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n650), .A2(new_n656), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(G232gat), .A2(G233gat), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(KEYINPUT41), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT95), .ZN(new_n663));
  XNOR2_X1  g462(.A(G134gat), .B(G162gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n627), .B1(new_n230), .B2(KEYINPUT17), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n667), .B1(new_n238), .B2(new_n239), .ZN(new_n668));
  XOR2_X1   g467(.A(G190gat), .B(G218gat), .Z(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  AOI22_X1  g469(.A1(new_n236), .A2(new_n627), .B1(KEYINPUT41), .B2(new_n661), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n668), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n670), .B1(new_n668), .B2(new_n671), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n666), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n674), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n676), .A2(new_n665), .A3(new_n672), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n644), .A2(new_n659), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n579), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(new_n523), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g481(.A1(new_n680), .A2(new_n520), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n684), .A2(G8gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT16), .B(G8gat), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT42), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n688), .B1(KEYINPUT42), .B2(new_n687), .ZN(G1325gat));
  NAND2_X1  g488(.A1(new_n534), .A2(new_n536), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n690), .A2(KEYINPUT100), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(KEYINPUT100), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(G15gat), .B1(new_n680), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n527), .A2(new_n447), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n695), .A2(G15gat), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n680), .B2(new_n696), .ZN(G1326gat));
  NAND3_X1  g496(.A1(new_n579), .A2(new_n346), .A3(new_n679), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT43), .B(G22gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  NAND2_X1  g499(.A1(new_n531), .A2(new_n578), .ZN(new_n701));
  INV_X1    g500(.A(new_n644), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n659), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(new_n270), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n701), .A2(new_n678), .A3(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n705), .A2(G29gat), .A3(new_n523), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT45), .Z(new_n707));
  XOR2_X1   g506(.A(new_n704), .B(KEYINPUT101), .Z(new_n708));
  INV_X1    g507(.A(KEYINPUT102), .ZN(new_n709));
  OAI22_X1  g508(.A1(new_n513), .A2(new_n345), .B1(new_n533), .B2(new_n535), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n554), .B1(new_n568), .B2(new_n572), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT81), .ZN(new_n712));
  AOI211_X1 g511(.A(new_n709), .B(new_n710), .C1(new_n712), .C2(new_n573), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n573), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT102), .B1(new_n714), .B2(new_n537), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n531), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n675), .A2(new_n677), .A3(KEYINPUT103), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT103), .B1(new_n675), .B2(new_n677), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n716), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n720), .B1(new_n701), .B2(new_n678), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n708), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n484), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G29gat), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n707), .A2(new_n728), .ZN(G1328gat));
  NAND2_X1  g528(.A1(new_n726), .A2(new_n512), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G36gat), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n705), .A2(G36gat), .A3(new_n520), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT46), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(G1329gat));
  NOR3_X1   g533(.A1(new_n705), .A2(G43gat), .A3(new_n695), .ZN(new_n735));
  INV_X1    g534(.A(new_n693), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n726), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n735), .B1(new_n737), .B2(G43gat), .ZN(new_n738));
  INV_X1    g537(.A(G43gat), .ZN(new_n739));
  INV_X1    g538(.A(new_n690), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(new_n726), .B2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n742));
  OR2_X1    g541(.A1(new_n735), .A2(new_n742), .ZN(new_n743));
  OAI22_X1  g542(.A1(new_n738), .A2(KEYINPUT47), .B1(new_n741), .B2(new_n743), .ZN(G1330gat));
  NAND2_X1  g543(.A1(new_n579), .A2(new_n346), .ZN(new_n745));
  INV_X1    g544(.A(new_n678), .ZN(new_n746));
  NOR4_X1   g545(.A1(new_n745), .A2(G50gat), .A3(new_n746), .A4(new_n703), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n726), .A2(new_n346), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(G50gat), .ZN(new_n749));
  XNOR2_X1  g548(.A(KEYINPUT104), .B(KEYINPUT48), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n749), .B(new_n750), .Z(G1331gat));
  AND3_X1   g550(.A1(new_n514), .A2(new_n525), .A3(new_n530), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n578), .A2(new_n709), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n714), .A2(KEYINPUT102), .A3(new_n537), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n659), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n270), .A2(new_n756), .A3(new_n746), .A4(new_n644), .ZN(new_n757));
  OR3_X1    g556(.A1(new_n755), .A2(KEYINPUT105), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT105), .B1(new_n755), .B2(new_n757), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n523), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(new_n598), .ZN(G1332gat));
  NOR2_X1   g561(.A1(new_n760), .A2(new_n520), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  AND2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n763), .B2(new_n764), .ZN(G1333gat));
  NAND4_X1  g566(.A1(new_n758), .A2(G71gat), .A3(new_n736), .A4(new_n759), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT106), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n605), .B1(new_n760), .B2(new_n695), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT50), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n769), .A2(new_n773), .A3(new_n770), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(G1334gat));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n345), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(new_n606), .ZN(G1335gat));
  OAI21_X1  g576(.A(KEYINPUT107), .B1(new_n755), .B2(new_n746), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT107), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n716), .A2(new_n779), .A3(new_n678), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n756), .A2(new_n269), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n778), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n778), .A2(new_n780), .A3(KEYINPUT51), .A4(new_n781), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n702), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n786), .A2(new_n584), .A3(new_n484), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n781), .A2(new_n644), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n788), .B1(new_n723), .B2(new_n725), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(G85gat), .B1(new_n790), .B2(new_n523), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n787), .A2(new_n791), .ZN(G1336gat));
  AOI21_X1  g591(.A(new_n585), .B1(new_n789), .B2(new_n512), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT109), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n795), .B(new_n796), .C1(new_n793), .C2(KEYINPUT108), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n702), .A2(G92gat), .A3(new_n520), .ZN(new_n798));
  INV_X1    g597(.A(new_n781), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n755), .A2(new_n746), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n799), .B1(new_n800), .B2(new_n779), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT51), .B1(new_n801), .B2(new_n778), .ZN(new_n802));
  INV_X1    g601(.A(new_n785), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n798), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n788), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n753), .A2(new_n754), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n721), .B1(new_n806), .B2(new_n531), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n512), .B(new_n805), .C1(new_n807), .C2(new_n724), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT108), .B1(new_n808), .B2(G92gat), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT109), .B1(new_n809), .B2(KEYINPUT52), .ZN(new_n810));
  AND4_X1   g609(.A1(new_n794), .A2(new_n797), .A3(new_n804), .A4(new_n810), .ZN(new_n811));
  AOI22_X1  g610(.A1(new_n810), .A2(new_n797), .B1(new_n804), .B2(new_n794), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(G1337gat));
  XOR2_X1   g612(.A(KEYINPUT110), .B(G99gat), .Z(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n695), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n815), .B1(new_n786), .B2(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n790), .A2(new_n693), .A3(new_n814), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT111), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n820));
  INV_X1    g619(.A(new_n818), .ZN(new_n821));
  AOI211_X1 g620(.A(new_n695), .B(new_n702), .C1(new_n784), .C2(new_n785), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n820), .B(new_n821), .C1(new_n822), .C2(new_n815), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n823), .ZN(G1338gat));
  NOR2_X1   g623(.A1(new_n345), .A2(G106gat), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n644), .B(new_n825), .C1(new_n802), .C2(new_n803), .ZN(new_n826));
  OR2_X1    g625(.A1(KEYINPUT113), .A2(KEYINPUT53), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n789), .A2(new_n346), .ZN(new_n828));
  XOR2_X1   g627(.A(KEYINPUT112), .B(G106gat), .Z(new_n829));
  AOI22_X1  g628(.A1(new_n828), .A2(new_n829), .B1(KEYINPUT113), .B2(KEYINPUT53), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n826), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n827), .B1(new_n826), .B2(new_n830), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(G1339gat));
  NOR2_X1   g632(.A1(new_n270), .A2(G113gat), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n835), .B(new_n581), .C1(new_n629), .C2(new_n631), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n639), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n626), .A2(new_n628), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n631), .B1(new_n839), .B2(new_n630), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n633), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(KEYINPUT54), .A3(new_n632), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n843), .A2(new_n844), .B1(new_n640), .B2(new_n641), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n632), .A2(KEYINPUT54), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n837), .B1(new_n847), .B2(new_n841), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n846), .B1(new_n848), .B2(KEYINPUT55), .ZN(new_n849));
  AND4_X1   g648(.A1(new_n846), .A2(new_n838), .A3(new_n842), .A4(KEYINPUT55), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n845), .B(new_n269), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n266), .A2(new_n267), .A3(new_n262), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n253), .A2(new_n244), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n246), .A2(new_n247), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n261), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n644), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n719), .B1(new_n851), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n848), .A2(new_n846), .A3(KEYINPUT55), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n838), .A2(new_n842), .A3(KEYINPUT55), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT114), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  AND4_X1   g661(.A1(new_n719), .A2(new_n862), .A3(new_n856), .A4(new_n845), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n659), .B1(new_n858), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n679), .A2(new_n270), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT115), .ZN(new_n867));
  INV_X1    g666(.A(new_n519), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT115), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n864), .A2(new_n869), .A3(new_n865), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n867), .A2(new_n484), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT116), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n520), .B(new_n834), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n867), .A2(new_n870), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n523), .A2(new_n512), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n450), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(G113gat), .B1(new_n878), .B2(new_n270), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT117), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n875), .A2(new_n882), .A3(new_n879), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(G1340gat));
  NOR2_X1   g683(.A1(new_n702), .A2(G120gat), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n520), .B(new_n885), .C1(new_n873), .C2(new_n874), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n887));
  OAI21_X1  g686(.A(G120gat), .B1(new_n878), .B2(new_n702), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n887), .B1(new_n886), .B2(new_n888), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(G1341gat));
  NOR2_X1   g690(.A1(new_n659), .A2(G127gat), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n520), .B(new_n892), .C1(new_n873), .C2(new_n874), .ZN(new_n893));
  OAI21_X1  g692(.A(G127gat), .B1(new_n878), .B2(new_n659), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT119), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n893), .A2(KEYINPUT119), .A3(new_n894), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1342gat));
  NAND2_X1  g698(.A1(new_n678), .A2(new_n520), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(G134gat), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n901), .B1(new_n873), .B2(new_n874), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n902), .A2(KEYINPUT56), .ZN(new_n903));
  OAI21_X1  g702(.A(G134gat), .B1(new_n878), .B2(new_n746), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(KEYINPUT56), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(G1343gat));
  NOR2_X1   g705(.A1(new_n736), .A2(new_n345), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n867), .A2(new_n870), .A3(new_n877), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n269), .A2(new_n294), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n851), .A2(new_n857), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT120), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n851), .A2(new_n913), .A3(new_n857), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n912), .A2(new_n746), .A3(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n863), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n756), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(new_n865), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n346), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT57), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT57), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n867), .A2(new_n921), .A3(new_n346), .A4(new_n870), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n690), .A2(new_n877), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n920), .A2(new_n269), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n910), .B1(new_n924), .B2(G141gat), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT121), .B1(new_n908), .B2(new_n909), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT58), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT122), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n926), .A2(new_n929), .A3(KEYINPUT58), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n925), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n924), .A2(G141gat), .ZN(new_n932));
  INV_X1    g731(.A(new_n910), .ZN(new_n933));
  AOI22_X1  g732(.A1(new_n928), .A2(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n931), .A2(new_n934), .ZN(G1344gat));
  INV_X1    g734(.A(new_n908), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n936), .A2(new_n296), .A3(new_n644), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n938), .A2(new_n702), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n939), .A2(KEYINPUT59), .A3(new_n296), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT59), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n867), .A2(new_n870), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT57), .B1(new_n942), .B2(new_n345), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n862), .A2(new_n678), .A3(new_n856), .A4(new_n845), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n756), .B1(new_n915), .B2(new_n944), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n921), .B(new_n346), .C1(new_n945), .C2(new_n918), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n943), .A2(new_n644), .A3(new_n923), .A4(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n941), .B1(new_n947), .B2(G148gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n937), .B1(new_n940), .B2(new_n948), .ZN(G1345gat));
  OAI21_X1  g748(.A(G155gat), .B1(new_n938), .B2(new_n659), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n936), .A2(new_n300), .A3(new_n756), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(G1346gat));
  INV_X1    g751(.A(new_n719), .ZN(new_n953));
  OAI21_X1  g752(.A(G162gat), .B1(new_n938), .B2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(new_n907), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n955), .A2(G162gat), .A3(new_n900), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n876), .A2(new_n956), .A3(new_n484), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n954), .A2(new_n957), .ZN(G1347gat));
  NOR2_X1   g757(.A1(new_n484), .A2(new_n520), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n876), .A2(new_n450), .A3(new_n959), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n960), .A2(new_n380), .A3(new_n270), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n942), .A2(new_n484), .A3(new_n520), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n963), .A2(new_n519), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(new_n269), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n961), .B1(new_n965), .B2(new_n380), .ZN(G1348gat));
  NAND3_X1  g765(.A1(new_n964), .A2(new_n381), .A3(new_n644), .ZN(new_n967));
  OAI21_X1  g766(.A(G176gat), .B1(new_n960), .B2(new_n702), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(G1349gat));
  INV_X1    g768(.A(KEYINPUT123), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n970), .A2(KEYINPUT60), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n970), .A2(KEYINPUT60), .ZN(new_n972));
  OAI21_X1  g771(.A(G183gat), .B1(new_n960), .B2(new_n659), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n756), .A2(new_n396), .A3(new_n398), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n962), .A2(new_n868), .A3(new_n974), .ZN(new_n975));
  AOI211_X1 g774(.A(new_n971), .B(new_n972), .C1(new_n973), .C2(new_n975), .ZN(new_n976));
  AND4_X1   g775(.A1(new_n970), .A2(new_n973), .A3(KEYINPUT60), .A4(new_n975), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n976), .A2(new_n977), .ZN(G1350gat));
  NAND3_X1  g777(.A1(new_n964), .A2(new_n368), .A3(new_n719), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n962), .A2(new_n450), .A3(new_n678), .ZN(new_n980));
  NOR2_X1   g779(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n368), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n981), .B1(new_n980), .B2(new_n982), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n979), .B1(new_n984), .B2(new_n985), .ZN(G1351gat));
  INV_X1    g785(.A(G197gat), .ZN(new_n987));
  AND2_X1   g786(.A1(new_n693), .A2(new_n959), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n943), .A2(new_n269), .A3(new_n946), .A4(new_n988), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n987), .B1(new_n989), .B2(KEYINPUT125), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n990), .B1(KEYINPUT125), .B2(new_n989), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n876), .A2(new_n907), .A3(new_n959), .ZN(new_n992));
  INV_X1    g791(.A(new_n992), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n993), .A2(new_n987), .A3(new_n269), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n991), .A2(new_n994), .ZN(G1352gat));
  INV_X1    g794(.A(KEYINPUT126), .ZN(new_n996));
  AOI211_X1 g795(.A(G204gat), .B(new_n702), .C1(new_n996), .C2(KEYINPUT62), .ZN(new_n997));
  INV_X1    g796(.A(new_n997), .ZN(new_n998));
  OR4_X1    g797(.A1(new_n996), .A2(new_n992), .A3(KEYINPUT62), .A4(new_n998), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n943), .A2(new_n946), .A3(new_n988), .ZN(new_n1000));
  OAI21_X1  g799(.A(G204gat), .B1(new_n1000), .B2(new_n702), .ZN(new_n1001));
  OAI22_X1  g800(.A1(new_n992), .A2(new_n998), .B1(new_n996), .B2(KEYINPUT62), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n999), .A2(new_n1001), .A3(new_n1002), .ZN(G1353gat));
  NAND3_X1  g802(.A1(new_n993), .A2(new_n283), .A3(new_n756), .ZN(new_n1004));
  NAND4_X1  g803(.A1(new_n943), .A2(new_n756), .A3(new_n946), .A4(new_n988), .ZN(new_n1005));
  AND3_X1   g804(.A1(new_n1005), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1006));
  AOI21_X1  g805(.A(KEYINPUT63), .B1(new_n1005), .B2(G211gat), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(G1354gat));
  OAI21_X1  g807(.A(new_n274), .B1(new_n992), .B2(new_n953), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT127), .ZN(new_n1010));
  XNOR2_X1  g809(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  NOR3_X1   g810(.A1(new_n1000), .A2(new_n316), .A3(new_n746), .ZN(new_n1012));
  NOR2_X1   g811(.A1(new_n1011), .A2(new_n1012), .ZN(G1355gat));
endmodule


