//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G110), .B(G140), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G227), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n191), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT66), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT66), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G134), .ZN(new_n198));
  INV_X1    g012(.A(G137), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT68), .B(G131), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n200), .A2(KEYINPUT67), .A3(new_n201), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n199), .A2(KEYINPUT11), .A3(G134), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n196), .A2(new_n198), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G137), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n204), .A2(new_n206), .A3(new_n207), .A4(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT69), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n204), .A2(new_n213), .A3(new_n207), .A4(new_n211), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G131), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT67), .B1(new_n200), .B2(new_n201), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT66), .B(G134), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n208), .B1(new_n217), .B2(new_n199), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n213), .B1(new_n219), .B2(new_n207), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n212), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G101), .ZN(new_n222));
  INV_X1    g036(.A(G104), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G107), .ZN(new_n224));
  INV_X1    g038(.A(G107), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G104), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n222), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n228), .B1(new_n223), .B2(G107), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n225), .A2(KEYINPUT3), .A3(G104), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n229), .A2(new_n230), .B1(new_n223), .B2(G107), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n227), .B1(new_n231), .B2(new_n222), .ZN(new_n232));
  INV_X1    g046(.A(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G143), .ZN(new_n234));
  INV_X1    g048(.A(G143), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G146), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT1), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n234), .A2(new_n236), .A3(new_n237), .A4(G128), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n234), .A2(new_n236), .ZN(new_n239));
  INV_X1    g053(.A(G128), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(new_n234), .B2(KEYINPUT1), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n238), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n232), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT64), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n236), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n235), .A2(KEYINPUT64), .A3(G146), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n245), .A2(new_n246), .B1(G143), .B2(new_n233), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n238), .B1(new_n247), .B2(new_n241), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n243), .B1(new_n248), .B2(new_n232), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n221), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT12), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT0), .B(G128), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n245), .A2(new_n246), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n253), .B1(new_n254), .B2(new_n234), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT65), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n234), .A2(new_n236), .A3(G128), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n255), .A2(new_n256), .B1(KEYINPUT0), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n259), .B1(new_n231), .B2(new_n222), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n260), .B1(new_n222), .B2(new_n231), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT65), .B1(new_n247), .B2(new_n253), .ZN(new_n262));
  OR3_X1    g076(.A1(new_n231), .A2(KEYINPUT4), .A3(new_n222), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n258), .A2(new_n261), .A3(new_n262), .A4(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n248), .A2(KEYINPUT10), .A3(new_n232), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT10), .B1(new_n232), .B2(new_n242), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n266), .A2(KEYINPUT79), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(KEYINPUT79), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n264), .B(new_n265), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT80), .B1(new_n269), .B2(new_n221), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n264), .A2(new_n265), .ZN(new_n271));
  INV_X1    g085(.A(new_n221), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT80), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n266), .B(KEYINPUT79), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n271), .A2(new_n272), .A3(new_n273), .A4(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n194), .B1(new_n252), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n272), .B1(new_n274), .B2(new_n271), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n194), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n280), .B1(new_n270), .B2(new_n275), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n277), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(G469), .B1(new_n282), .B2(G902), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n276), .A2(new_n279), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(KEYINPUT81), .A3(new_n280), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT81), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n278), .B1(new_n275), .B2(new_n270), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n286), .B1(new_n287), .B2(new_n194), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n281), .A2(new_n252), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n285), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G469), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n190), .B1(new_n283), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G214), .B1(G237), .B2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n255), .A2(new_n256), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n257), .A2(KEYINPUT0), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n262), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G125), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(G125), .B2(new_n248), .ZN(new_n301));
  INV_X1    g115(.A(G224), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(G953), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G113), .ZN(new_n305));
  INV_X1    g119(.A(G116), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(G119), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT5), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OR3_X1    g123(.A1(new_n306), .A2(KEYINPUT71), .A3(G119), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT71), .B1(new_n306), .B2(G119), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(new_n307), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n309), .B1(new_n312), .B2(new_n308), .ZN(new_n313));
  NOR2_X1   g127(.A1(KEYINPUT2), .A2(G113), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT2), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT70), .B1(new_n315), .B2(new_n305), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT70), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(KEYINPUT2), .A3(G113), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n314), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n319), .B(new_n310), .C1(new_n307), .C2(new_n311), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n232), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OR2_X1    g137(.A1(new_n323), .A2(KEYINPUT85), .ZN(new_n324));
  OR2_X1    g138(.A1(new_n312), .A2(new_n308), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  XOR2_X1   g140(.A(new_n309), .B(KEYINPUT84), .Z(new_n327));
  OAI211_X1 g141(.A(new_n232), .B(new_n320), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(KEYINPUT85), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n324), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  XOR2_X1   g144(.A(G110), .B(G122), .Z(new_n331));
  XOR2_X1   g145(.A(new_n331), .B(KEYINPUT8), .Z(new_n332));
  AOI22_X1  g146(.A1(new_n304), .A2(KEYINPUT7), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n301), .A2(new_n303), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT7), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n301), .A2(new_n335), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n316), .A2(new_n318), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n312), .B1(new_n337), .B2(new_n314), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n320), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n261), .A3(new_n263), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n313), .A2(new_n320), .A3(new_n232), .ZN(new_n341));
  INV_X1    g155(.A(new_n331), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n334), .A2(new_n336), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(G902), .B1(new_n333), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n301), .B(new_n303), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n343), .A2(KEYINPUT6), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n340), .A2(new_n341), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n331), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(KEYINPUT82), .A3(new_n349), .ZN(new_n350));
  XOR2_X1   g164(.A(KEYINPUT83), .B(KEYINPUT6), .Z(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n348), .A2(KEYINPUT82), .A3(new_n331), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n352), .B1(new_n347), .B2(new_n353), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n346), .B(new_n350), .C1(new_n354), .C2(new_n349), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n345), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(G210), .B1(G237), .B2(G902), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n345), .A2(new_n355), .A3(new_n357), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n296), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G237), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(new_n192), .A3(G214), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(new_n235), .ZN(new_n364));
  NAND2_X1  g178(.A1(KEYINPUT18), .A2(G131), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n364), .B(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(G125), .B(G140), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(new_n233), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(KEYINPUT16), .ZN(new_n370));
  INV_X1    g184(.A(G125), .ZN(new_n371));
  OR3_X1    g185(.A1(new_n371), .A2(KEYINPUT16), .A3(G140), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(G146), .A3(new_n372), .ZN(new_n373));
  XOR2_X1   g187(.A(new_n367), .B(KEYINPUT19), .Z(new_n374));
  NAND2_X1  g188(.A1(new_n364), .A2(new_n205), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n363), .B(G143), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n206), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT86), .ZN(new_n379));
  OAI221_X1 g193(.A(new_n373), .B1(G146), .B2(new_n374), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT86), .B1(new_n375), .B2(new_n377), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n369), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(G113), .B(G122), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n383), .B(new_n223), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n378), .A2(KEYINPUT17), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n370), .A2(new_n372), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n233), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT17), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n373), .B(new_n389), .C1(new_n375), .C2(new_n390), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n369), .B(new_n384), .C1(new_n387), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT20), .ZN(new_n394));
  NOR2_X1   g208(.A1(G475), .A2(G902), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n395), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n393), .A2(KEYINPUT87), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT87), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n386), .A2(new_n399), .A3(new_n392), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n397), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n396), .B1(new_n401), .B2(new_n394), .ZN(new_n402));
  INV_X1    g216(.A(G475), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n369), .B1(new_n387), .B2(new_n391), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n385), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n392), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n403), .B1(new_n406), .B2(new_n292), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(G116), .B(G122), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(new_n225), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n306), .A2(G122), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(KEYINPUT14), .A3(G107), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n410), .A2(KEYINPUT14), .A3(new_n412), .A4(G107), .ZN(new_n415));
  XOR2_X1   g229(.A(G128), .B(G143), .Z(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(new_n217), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT89), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT13), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n240), .B2(G143), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(G128), .B2(new_n235), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n421), .A2(new_n240), .A3(G143), .ZN(new_n424));
  OAI21_X1  g238(.A(G134), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT88), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n416), .A2(new_n217), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n426), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n427), .A2(new_n411), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n420), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G217), .ZN(new_n432));
  NOR3_X1   g246(.A1(new_n188), .A2(new_n432), .A3(G953), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n433), .B1(new_n420), .B2(new_n430), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n292), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT15), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G478), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n437), .A2(new_n439), .A3(G478), .ZN(new_n442));
  INV_X1    g256(.A(G952), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n443), .A2(KEYINPUT90), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n443), .A2(KEYINPUT90), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n192), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(G234), .B2(G237), .ZN(new_n447));
  XOR2_X1   g261(.A(KEYINPUT21), .B(G898), .Z(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(KEYINPUT92), .ZN(new_n449));
  NAND2_X1  g263(.A1(G234), .A2(G237), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(G902), .A3(G953), .ZN(new_n451));
  XOR2_X1   g265(.A(new_n451), .B(KEYINPUT91), .Z(new_n452));
  AOI21_X1  g266(.A(new_n447), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n441), .A2(new_n442), .A3(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n409), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n294), .A2(new_n361), .A3(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(KEYINPUT93), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT73), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT30), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT11), .B1(new_n217), .B2(new_n199), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n211), .B1(new_n461), .B2(KEYINPUT67), .ZN(new_n462));
  INV_X1    g276(.A(new_n207), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT69), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(G131), .A3(new_n214), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n299), .B1(new_n465), .B2(new_n212), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n200), .B1(G134), .B2(new_n199), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G131), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n212), .A2(new_n248), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n460), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n299), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n221), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(KEYINPUT30), .A3(new_n469), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n471), .A2(new_n339), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n362), .A2(new_n192), .A3(G210), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n476), .B(new_n222), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n478));
  XOR2_X1   g292(.A(new_n477), .B(new_n478), .Z(new_n479));
  INV_X1    g293(.A(KEYINPUT72), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n470), .B1(new_n221), .B2(new_n472), .ZN(new_n481));
  INV_X1    g295(.A(new_n339), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR4_X1   g297(.A1(new_n466), .A2(KEYINPUT72), .A3(new_n339), .A4(new_n470), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n475), .B(new_n479), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT31), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n473), .A2(new_n482), .A3(new_n469), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT72), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n481), .A2(new_n480), .A3(new_n482), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT31), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n479), .A4(new_n475), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n339), .B1(new_n466), .B2(new_n470), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n494), .B1(new_n484), .B2(new_n483), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT28), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT28), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n487), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n479), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n459), .B1(new_n493), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n481), .A2(new_n482), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n501), .B1(new_n488), .B2(new_n489), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n498), .B1(new_n502), .B2(new_n497), .ZN(new_n503));
  INV_X1    g317(.A(new_n479), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n505), .A2(KEYINPUT73), .A3(new_n486), .A4(new_n492), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(G472), .A2(G902), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT74), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT32), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n507), .A2(KEYINPUT32), .A3(new_n509), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT29), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n490), .A2(new_n475), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n504), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n514), .B(new_n516), .C1(new_n503), .C2(new_n504), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n496), .A2(KEYINPUT75), .B1(new_n497), .B2(new_n487), .ZN(new_n518));
  OR3_X1    g332(.A1(new_n502), .A2(KEYINPUT75), .A3(new_n497), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n479), .A2(KEYINPUT29), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n517), .B(new_n292), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G472), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n512), .A2(new_n513), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT23), .B1(new_n240), .B2(G119), .ZN(new_n525));
  INV_X1    g339(.A(G119), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT76), .B1(new_n526), .B2(G128), .ZN(new_n527));
  XOR2_X1   g341(.A(new_n525), .B(new_n527), .Z(new_n528));
  XNOR2_X1  g342(.A(G119), .B(G128), .ZN(new_n529));
  XOR2_X1   g343(.A(KEYINPUT24), .B(G110), .Z(new_n530));
  OAI22_X1  g344(.A1(new_n528), .A2(G110), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n367), .A2(new_n233), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(new_n373), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n528), .A2(G110), .B1(new_n529), .B2(new_n530), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n389), .A2(new_n373), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(KEYINPUT77), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT22), .B(G137), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n533), .A2(new_n536), .A3(new_n541), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(G902), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT78), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT25), .ZN(new_n548));
  OR2_X1    g362(.A1(new_n547), .A2(KEYINPUT25), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n432), .B1(G234), .B2(new_n292), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n550), .B(new_n551), .C1(new_n546), .C2(new_n548), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n545), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n551), .A2(G902), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n458), .A2(new_n524), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(G101), .ZN(G3));
  AOI21_X1  g372(.A(G902), .B1(new_n500), .B2(new_n506), .ZN(new_n559));
  INV_X1    g373(.A(G472), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(new_n507), .B2(new_n509), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(new_n294), .A3(new_n556), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT94), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n435), .A2(KEYINPUT33), .A3(new_n436), .ZN(new_n565));
  INV_X1    g379(.A(new_n435), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n431), .A2(KEYINPUT96), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n434), .A2(KEYINPUT95), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n566), .A2(KEYINPUT96), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n567), .B2(new_n568), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n565), .B1(new_n570), .B2(KEYINPUT33), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n292), .A2(G478), .ZN(new_n572));
  OAI22_X1  g386(.A1(new_n571), .A2(new_n572), .B1(G478), .B2(new_n438), .ZN(new_n573));
  AND4_X1   g387(.A1(new_n361), .A2(new_n573), .A3(new_n409), .A4(new_n454), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n564), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g389(.A(KEYINPUT34), .B(G104), .Z(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(G6));
  NOR2_X1   g391(.A1(new_n401), .A2(new_n394), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n401), .A2(new_n394), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n407), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT97), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n441), .A2(new_n442), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n581), .A2(new_n582), .A3(new_n583), .A4(new_n454), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n401), .A2(new_n394), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n408), .B(new_n583), .C1(new_n585), .C2(new_n578), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT97), .B1(new_n586), .B2(new_n453), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n584), .A2(new_n587), .A3(new_n361), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n564), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(KEYINPUT98), .ZN(new_n590));
  XOR2_X1   g404(.A(KEYINPUT35), .B(G107), .Z(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G9));
  INV_X1    g406(.A(KEYINPUT99), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n533), .A2(new_n593), .A3(new_n536), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n593), .B1(new_n533), .B2(new_n536), .ZN(new_n596));
  OAI22_X1  g410(.A1(new_n595), .A2(new_n596), .B1(KEYINPUT36), .B2(new_n542), .ZN(new_n597));
  INV_X1    g411(.A(new_n596), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n542), .A2(KEYINPUT36), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n599), .A3(new_n594), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(KEYINPUT100), .A3(new_n555), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT100), .ZN(new_n603));
  INV_X1    g417(.A(new_n601), .ZN(new_n604));
  INV_X1    g418(.A(new_n555), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n552), .A2(new_n602), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n458), .A2(new_n562), .A3(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT37), .B(G110), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G12));
  AND3_X1   g424(.A1(new_n294), .A2(new_n361), .A3(new_n607), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n524), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(G900), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n447), .B1(new_n452), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n586), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(G128), .ZN(G30));
  XOR2_X1   g431(.A(new_n614), .B(KEYINPUT39), .Z(new_n618));
  NAND2_X1  g432(.A1(new_n294), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n619), .B(KEYINPUT102), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT40), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n622), .B1(new_n502), .B2(new_n479), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n495), .A2(KEYINPUT101), .A3(new_n504), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n623), .A2(new_n485), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(G472), .B1(new_n625), .B2(G902), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n512), .A2(new_n513), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n359), .A2(new_n360), .ZN(new_n628));
  XOR2_X1   g442(.A(new_n628), .B(KEYINPUT38), .Z(new_n629));
  NAND2_X1  g443(.A1(new_n409), .A2(new_n583), .ZN(new_n630));
  NOR4_X1   g444(.A1(new_n629), .A2(new_n296), .A3(new_n607), .A4(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n621), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G143), .ZN(G45));
  NAND2_X1  g447(.A1(new_n573), .A2(new_n409), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(new_n614), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n612), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G146), .ZN(G48));
  AND3_X1   g451(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n291), .B1(new_n290), .B2(new_n292), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n190), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n524), .A2(new_n556), .A3(new_n574), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT103), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT41), .B(G113), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G15));
  NAND4_X1  g460(.A1(new_n524), .A2(new_n556), .A3(new_n588), .A4(new_n642), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G116), .ZN(G18));
  NAND2_X1  g462(.A1(new_n456), .A2(new_n607), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n640), .A2(KEYINPUT104), .A3(new_n361), .A4(new_n189), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n290), .A2(new_n292), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(G469), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n652), .A2(new_n361), .A3(new_n189), .A4(new_n293), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n649), .B1(new_n650), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n524), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G119), .ZN(G21));
  AOI21_X1  g472(.A(new_n479), .B1(new_n518), .B2(new_n519), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n509), .B1(new_n659), .B2(new_n493), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n556), .B(new_n660), .C1(new_n559), .C2(new_n560), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n653), .A2(new_n453), .A3(new_n630), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G122), .ZN(G24));
  OAI211_X1 g479(.A(new_n607), .B(new_n660), .C1(new_n559), .C2(new_n560), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n650), .A2(new_n655), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n667), .A2(new_n668), .A3(new_n635), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G125), .ZN(G27));
  NOR2_X1   g484(.A1(new_n628), .A2(new_n296), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n294), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n524), .A2(new_n556), .A3(new_n635), .A4(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G131), .ZN(G33));
  XNOR2_X1  g493(.A(new_n615), .B(KEYINPUT105), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n524), .A2(new_n680), .A3(new_n556), .A4(new_n673), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G134), .ZN(G36));
  NAND3_X1  g496(.A1(new_n573), .A2(new_n408), .A3(new_n402), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT43), .Z(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n607), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n562), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT44), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n671), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n282), .A2(KEYINPUT45), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n282), .A2(KEYINPUT45), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n689), .A2(G469), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(G469), .A2(G902), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n691), .A2(KEYINPUT46), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(KEYINPUT46), .B1(new_n691), .B2(new_n692), .ZN(new_n694));
  OR3_X1    g508(.A1(new_n693), .A2(new_n694), .A3(new_n638), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n189), .A3(new_n618), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT106), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n686), .A2(KEYINPUT44), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n688), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(new_n199), .ZN(G39));
  NAND2_X1  g514(.A1(new_n695), .A2(new_n189), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT47), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n512), .A2(new_n513), .ZN(new_n703));
  INV_X1    g517(.A(new_n671), .ZN(new_n704));
  NOR4_X1   g518(.A1(new_n634), .A2(new_n704), .A3(new_n556), .A4(new_n614), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n703), .A2(new_n705), .A3(new_n523), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT107), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n708), .B(G140), .Z(G42));
  NAND2_X1  g523(.A1(new_n684), .A2(new_n447), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n642), .A2(new_n671), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n524), .A2(new_n556), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OR2_X1    g528(.A1(new_n714), .A2(KEYINPUT48), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(KEYINPUT48), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n710), .A2(new_n661), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n446), .B1(new_n717), .B2(new_n668), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n715), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n703), .A2(new_n556), .A3(new_n626), .ZN(new_n720));
  INV_X1    g534(.A(new_n447), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n720), .A2(new_n721), .A3(new_n711), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT120), .ZN(new_n723));
  OR3_X1    g537(.A1(new_n723), .A2(new_n409), .A3(new_n573), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n642), .A2(new_n296), .A3(new_n629), .ZN(new_n725));
  XOR2_X1   g539(.A(new_n725), .B(KEYINPUT118), .Z(new_n726));
  NAND2_X1  g540(.A1(new_n717), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(new_n727), .B(KEYINPUT50), .Z(new_n728));
  NAND2_X1  g542(.A1(new_n712), .A2(new_n667), .ZN(new_n729));
  XOR2_X1   g543(.A(new_n729), .B(KEYINPUT119), .Z(new_n730));
  NAND3_X1  g544(.A1(new_n724), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n717), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n704), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n640), .A2(new_n190), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n702), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT51), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  OAI221_X1 g551(.A(new_n719), .B1(new_n634), .B2(new_n723), .C1(new_n731), .C2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT121), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n731), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n724), .A2(new_n728), .A3(new_n730), .A4(KEYINPUT121), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n702), .A2(KEYINPUT116), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n735), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n702), .A2(KEYINPUT116), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n733), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n745), .A2(KEYINPUT117), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(KEYINPUT117), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n740), .A2(new_n741), .A3(new_n746), .A4(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n738), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n524), .B(new_n611), .C1(new_n615), .C2(new_n635), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n614), .B(KEYINPUT111), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n607), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n294), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n294), .A2(KEYINPUT112), .A3(new_n753), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n361), .A2(new_n409), .A3(new_n583), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n627), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n751), .A2(new_n669), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT113), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(KEYINPUT52), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT114), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n751), .A2(new_n766), .A3(new_n761), .A4(new_n669), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n764), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n765), .B1(new_n764), .B2(new_n767), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n763), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n764), .A2(new_n767), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT114), .ZN(new_n773));
  INV_X1    g587(.A(new_n763), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n774), .A3(new_n768), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n583), .A2(new_n614), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n581), .A2(new_n607), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n524), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n667), .A2(new_n635), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n672), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AND4_X1   g596(.A1(new_n524), .A2(new_n680), .A3(new_n556), .A4(new_n673), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n777), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI22_X1  g598(.A1(new_n524), .A2(new_n779), .B1(new_n667), .B2(new_n635), .ZN(new_n785));
  OAI211_X1 g599(.A(KEYINPUT110), .B(new_n681), .C1(new_n785), .C2(new_n672), .ZN(new_n786));
  AOI22_X1  g600(.A1(new_n784), .A2(new_n786), .B1(new_n677), .B2(new_n676), .ZN(new_n787));
  INV_X1    g601(.A(new_n583), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n634), .B1(new_n409), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n361), .A3(new_n454), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n608), .B(new_n557), .C1(new_n563), .C2(new_n790), .ZN(new_n791));
  AOI22_X1  g605(.A1(new_n656), .A2(new_n524), .B1(new_n662), .B2(new_n663), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n643), .A3(new_n647), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT109), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT109), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n792), .A2(new_n643), .A3(new_n647), .A4(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n791), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n787), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n764), .A2(new_n767), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n787), .A2(new_n797), .A3(new_n800), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n776), .A2(new_n799), .B1(KEYINPUT53), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT54), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n791), .A2(new_n798), .A3(new_n793), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n787), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n769), .A2(new_n770), .A3(new_n763), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n774), .B1(new_n773), .B2(new_n768), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n801), .A2(new_n810), .A3(new_n798), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n810), .B1(new_n801), .B2(new_n798), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n809), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n814), .A2(KEYINPUT54), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n750), .A2(new_n803), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n816), .B1(G952), .B2(G953), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n683), .A2(new_n296), .A3(new_n190), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n641), .A2(KEYINPUT49), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n629), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n641), .A2(KEYINPUT49), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n720), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT108), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n817), .A2(new_n823), .ZN(G75));
  OR2_X1    g638(.A1(new_n354), .A2(new_n349), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n825), .A2(new_n350), .ZN(new_n826));
  XOR2_X1   g640(.A(new_n826), .B(new_n346), .Z(new_n827));
  XNOR2_X1  g641(.A(KEYINPUT122), .B(KEYINPUT55), .ZN(new_n828));
  XOR2_X1   g642(.A(new_n827), .B(new_n828), .Z(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT56), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT123), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n801), .A2(new_n798), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT115), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n835), .A2(new_n811), .B1(new_n776), .B2(new_n806), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n833), .B1(new_n836), .B2(new_n292), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n814), .A2(KEYINPUT123), .A3(G902), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n832), .B1(new_n839), .B2(new_n358), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n192), .A2(G952), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n835), .A2(new_n811), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n292), .B1(new_n843), .B2(new_n809), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT56), .B1(new_n844), .B2(G210), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n842), .B1(new_n845), .B2(new_n830), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT124), .B1(new_n840), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n814), .A2(G210), .A3(G902), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n831), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n841), .B1(new_n849), .B2(new_n829), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT124), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n357), .B1(new_n837), .B2(new_n838), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n850), .B(new_n851), .C1(new_n852), .C2(new_n832), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n847), .A2(new_n853), .ZN(G51));
  XNOR2_X1  g668(.A(new_n814), .B(KEYINPUT54), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n692), .B(KEYINPUT57), .Z(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n290), .ZN(new_n858));
  INV_X1    g672(.A(new_n691), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n839), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n841), .B1(new_n858), .B2(new_n860), .ZN(G54));
  AND2_X1   g675(.A1(KEYINPUT58), .A2(G475), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n836), .A2(new_n833), .A3(new_n292), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT123), .B1(new_n814), .B2(G902), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n398), .A2(new_n400), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n841), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n839), .A2(new_n869), .A3(new_n866), .A4(new_n862), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n866), .B(new_n862), .C1(new_n863), .C2(new_n864), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT125), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n868), .A2(new_n870), .A3(new_n872), .ZN(G60));
  INV_X1    g687(.A(new_n571), .ZN(new_n874));
  XOR2_X1   g688(.A(KEYINPUT126), .B(KEYINPUT59), .Z(new_n875));
  NAND2_X1  g689(.A1(G478), .A2(G902), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n875), .B(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n855), .A2(new_n874), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n815), .A2(new_n803), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n874), .B1(new_n879), .B2(new_n877), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n878), .A2(new_n880), .A3(new_n841), .ZN(G63));
  NAND2_X1  g695(.A1(G217), .A2(G902), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT60), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n836), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n601), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n545), .B1(new_n836), .B2(new_n883), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n885), .A2(new_n842), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT61), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n887), .B(new_n888), .ZN(G66));
  NOR2_X1   g703(.A1(new_n449), .A2(new_n302), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n890), .A2(new_n192), .ZN(new_n891));
  INV_X1    g705(.A(new_n797), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n891), .B1(new_n892), .B2(new_n192), .ZN(new_n893));
  INV_X1    g707(.A(G898), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n826), .B1(new_n894), .B2(G953), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n893), .B(new_n895), .ZN(G69));
  NAND3_X1  g710(.A1(new_n632), .A2(new_n669), .A3(new_n751), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT62), .Z(new_n898));
  NOR2_X1   g712(.A1(new_n699), .A2(new_n708), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n713), .A2(new_n620), .A3(new_n671), .A4(new_n789), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n471), .A2(new_n474), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n374), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n901), .A2(G953), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(G900), .A2(G953), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n713), .A2(new_n760), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n681), .B1(new_n697), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n751), .A2(new_n669), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n899), .A2(new_n678), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n905), .B1(new_n910), .B2(G953), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n904), .B1(new_n911), .B2(new_n903), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n912), .B(new_n913), .ZN(G72));
  NAND2_X1  g728(.A1(G472), .A2(G902), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT63), .Z(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(new_n910), .B2(new_n892), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n917), .A2(new_n490), .A3(new_n504), .A4(new_n475), .ZN(new_n918));
  INV_X1    g732(.A(new_n916), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n901), .B2(new_n797), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n515), .A2(new_n479), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n918), .B(new_n842), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n919), .B1(new_n516), .B2(new_n485), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n922), .B1(new_n802), .B2(new_n923), .ZN(G57));
endmodule


