//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n800,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(KEYINPUT22), .B2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G211gat), .B(G218gat), .Z(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT29), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT3), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G141gat), .B(G148gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n212), .B1(G155gat), .B2(G162gat), .ZN(new_n213));
  INV_X1    g012(.A(G155gat), .ZN(new_n214));
  INV_X1    g013(.A(G162gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI22_X1  g015(.A1(new_n211), .A2(new_n213), .B1(KEYINPUT80), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G155gat), .B(G162gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n210), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n209), .B1(new_n219), .B2(KEYINPUT3), .ZN(new_n222));
  INV_X1    g021(.A(new_n208), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G78gat), .B(G106gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G228gat), .A2(G233gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n227), .B(G22gat), .ZN(new_n228));
  XOR2_X1   g027(.A(KEYINPUT31), .B(G50gat), .Z(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n226), .B(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n232), .B(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT26), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT71), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G169gat), .ZN(new_n239));
  INV_X1    g038(.A(G176gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n240), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n241), .B1(KEYINPUT26), .B2(new_n242), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n238), .A2(new_n243), .B1(G183gat), .B2(G190gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT28), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT27), .B(G183gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G183gat), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n247), .B1(new_n249), .B2(KEYINPUT27), .ZN(new_n250));
  INV_X1    g049(.A(G190gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n245), .B1(new_n248), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n246), .A2(KEYINPUT28), .A3(new_n251), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n244), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g057(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n259));
  NOR2_X1   g058(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n242), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT66), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT66), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n242), .B(new_n263), .C1(new_n259), .C2(new_n260), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n266), .B1(new_n249), .B2(new_n251), .ZN(new_n267));
  NAND3_X1  g066(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n241), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n232), .A2(KEYINPUT23), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n265), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT25), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n272), .B1(new_n234), .B2(KEYINPUT23), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n274), .A2(new_n269), .A3(new_n265), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n258), .A2(new_n276), .ZN(new_n277));
  AND2_X1   g076(.A1(G226gat), .A2(G233gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(KEYINPUT29), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n273), .A2(KEYINPUT68), .A3(new_n275), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n284), .A2(new_n278), .A3(new_n258), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n280), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n208), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n284), .A2(new_n258), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(new_n279), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n258), .A2(new_n278), .A3(new_n276), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(new_n223), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G8gat), .B(G36gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(KEYINPUT78), .ZN(new_n294));
  XNOR2_X1  g093(.A(G64gat), .B(G92gat), .ZN(new_n295));
  XOR2_X1   g094(.A(new_n294), .B(new_n295), .Z(new_n296));
  NAND2_X1  g095(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n296), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n287), .A2(new_n291), .A3(KEYINPUT30), .A4(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n287), .A2(new_n291), .A3(new_n298), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT30), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(KEYINPUT79), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT79), .B1(new_n300), .B2(new_n301), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n297), .B(new_n299), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G134gat), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT72), .B1(new_n306), .B2(G127gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(G127gat), .B(G134gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n307), .B1(new_n308), .B2(KEYINPUT72), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(KEYINPUT73), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n311));
  INV_X1    g110(.A(G113gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(G120gat), .ZN(new_n313));
  INV_X1    g112(.A(G120gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n314), .A2(G113gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(KEYINPUT74), .A3(G113gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n318), .B1(G113gat), .B2(new_n314), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n313), .A2(KEYINPUT74), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n311), .B(new_n308), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT75), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n317), .A2(new_n323), .A3(new_n220), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n324), .A2(KEYINPUT4), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(KEYINPUT4), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n219), .B(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n317), .A2(new_n323), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n325), .A2(new_n326), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G225gat), .A2(G233gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n329), .A2(new_n219), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n333), .A2(KEYINPUT81), .A3(new_n324), .ZN(new_n334));
  INV_X1    g133(.A(new_n331), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT81), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n329), .A2(new_n336), .A3(new_n219), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT5), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n330), .A2(KEYINPUT5), .A3(new_n331), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(G1gat), .B(G29gat), .Z(new_n344));
  XNOR2_X1  g143(.A(G57gat), .B(G85gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT86), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n343), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n330), .A2(new_n331), .ZN(new_n352));
  XOR2_X1   g151(.A(KEYINPUT87), .B(KEYINPUT39), .Z(new_n353));
  AOI21_X1  g152(.A(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n334), .A2(new_n337), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n331), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n356), .B(KEYINPUT39), .C1(new_n331), .C2(new_n330), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT40), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n354), .A2(new_n357), .A3(KEYINPUT40), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n351), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n231), .B1(new_n305), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n300), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT37), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n287), .A2(new_n291), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT88), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n287), .A2(new_n291), .A3(KEYINPUT88), .A4(new_n365), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n365), .B1(new_n286), .B2(new_n223), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n289), .A2(new_n208), .A3(new_n290), .ZN(new_n372));
  AOI211_X1 g171(.A(KEYINPUT38), .B(new_n298), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n364), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n298), .B1(new_n292), .B2(KEYINPUT37), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT38), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n374), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n348), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n340), .A2(KEYINPUT6), .A3(new_n379), .A4(new_n341), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT84), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n380), .A2(new_n381), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT89), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OR2_X1    g183(.A1(new_n380), .A2(new_n381), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT89), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n380), .A2(new_n381), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT6), .B1(new_n342), .B2(new_n348), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n351), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n384), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n363), .B1(new_n378), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT77), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT76), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n395), .B1(new_n288), .B2(new_n329), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n288), .A2(new_n329), .ZN(new_n397));
  INV_X1    g196(.A(new_n329), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n284), .A2(new_n258), .A3(KEYINPUT76), .A4(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n396), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(G227gat), .A2(G233gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n401), .B(KEYINPUT64), .Z(new_n402));
  OR2_X1    g201(.A1(new_n402), .A2(KEYINPUT34), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n401), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT34), .B1(new_n400), .B2(new_n405), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT33), .B1(new_n400), .B2(new_n402), .ZN(new_n408));
  XOR2_X1   g207(.A(G15gat), .B(G43gat), .Z(new_n409));
  XNOR2_X1  g208(.A(G71gat), .B(G99gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT32), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n414), .B1(new_n400), .B2(new_n402), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  AOI221_X4 g216(.A(new_n414), .B1(KEYINPUT33), .B2(new_n411), .C1(new_n400), .C2(new_n402), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n407), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n415), .A2(new_n408), .A3(new_n412), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n421), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n394), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT36), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n417), .A2(new_n407), .A3(new_n419), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT77), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n424), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n382), .A2(new_n383), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n343), .A2(KEYINPUT83), .A3(new_n379), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT83), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n431), .B1(new_n342), .B2(new_n348), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n389), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n297), .A2(new_n299), .ZN(new_n435));
  INV_X1    g234(.A(new_n304), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n435), .B1(new_n436), .B2(new_n302), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n231), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT36), .B1(new_n420), .B2(new_n423), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n428), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n393), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n428), .A2(KEYINPUT85), .A3(new_n439), .A4(new_n440), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n422), .B1(new_n421), .B2(new_n418), .ZN(new_n445));
  INV_X1    g244(.A(new_n231), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(new_n426), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT35), .B1(new_n438), .B2(new_n447), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n305), .A2(KEYINPUT35), .A3(new_n231), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n424), .A2(new_n449), .A3(new_n427), .A4(new_n391), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n443), .A2(new_n444), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G15gat), .B(G22gat), .ZN(new_n452));
  INV_X1    g251(.A(G1gat), .ZN(new_n453));
  OR2_X1    g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(KEYINPUT16), .A3(new_n453), .ZN(new_n455));
  INV_X1    g254(.A(G8gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT92), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n456), .A2(KEYINPUT92), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n459), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT90), .ZN(new_n463));
  INV_X1    g262(.A(G29gat), .ZN(new_n464));
  INV_X1    g263(.A(G36gat), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(KEYINPUT90), .A2(G29gat), .A3(G36gat), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT14), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n468), .A2(new_n464), .A3(new_n465), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n466), .A2(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G43gat), .B(G50gat), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n471), .B1(KEYINPUT91), .B2(new_n472), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n473), .A2(KEYINPUT15), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n473), .B(KEYINPUT15), .C1(new_n472), .C2(new_n471), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n476), .A2(KEYINPUT17), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT17), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n478), .B1(new_n474), .B2(new_n475), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n462), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(G229gat), .A2(G233gat), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT93), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n462), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n460), .A2(KEYINPUT93), .A3(new_n461), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n484), .A3(new_n476), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n480), .A2(new_n481), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT18), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n481), .B(KEYINPUT13), .Z(new_n489));
  INV_X1    g288(.A(new_n485), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n476), .B1(new_n483), .B2(new_n484), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n480), .A2(KEYINPUT18), .A3(new_n485), .A4(new_n481), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n488), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G113gat), .B(G141gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(G197gat), .ZN(new_n496));
  XOR2_X1   g295(.A(KEYINPUT11), .B(G169gat), .Z(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(KEYINPUT12), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n488), .A2(new_n492), .A3(new_n499), .A4(new_n493), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n451), .A2(new_n504), .ZN(new_n505));
  XOR2_X1   g304(.A(G71gat), .B(G78gat), .Z(new_n506));
  AOI21_X1  g305(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT94), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G57gat), .B(G64gat), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n507), .B(KEYINPUT94), .ZN(new_n512));
  INV_X1    g311(.A(new_n506), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT95), .ZN(new_n514));
  INV_X1    g313(.A(G57gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n514), .B1(new_n515), .B2(G64gat), .ZN(new_n516));
  INV_X1    g315(.A(G64gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(KEYINPUT95), .A3(G57gat), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n516), .B(new_n518), .C1(G57gat), .C2(new_n517), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n512), .A2(new_n513), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n511), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT21), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G231gat), .A2(G233gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(G127gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n483), .A2(new_n484), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(new_n522), .B2(new_n521), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n527), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(new_n214), .ZN(new_n532));
  XNOR2_X1  g331(.A(G183gat), .B(G211gat), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n532), .B(new_n533), .Z(new_n534));
  OR2_X1    g333(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n530), .A2(new_n534), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G190gat), .B(G218gat), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT100), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g339(.A1(G232gat), .A2(G233gat), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n541), .A2(KEYINPUT41), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n540), .B(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G99gat), .A2(G106gat), .ZN(new_n545));
  INV_X1    g344(.A(G85gat), .ZN(new_n546));
  INV_X1    g345(.A(G92gat), .ZN(new_n547));
  AOI22_X1  g346(.A1(KEYINPUT8), .A2(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(KEYINPUT96), .A2(G85gat), .A3(G92gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT97), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT7), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT97), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n552), .A2(KEYINPUT96), .A3(G85gat), .A4(G92gat), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n551), .B1(new_n550), .B2(new_n553), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n548), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(G99gat), .ZN(new_n557));
  INV_X1    g356(.A(G106gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n545), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT98), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT98), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n559), .A2(new_n562), .A3(new_n545), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n556), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n564), .B(new_n548), .C1(new_n554), .C2(new_n555), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(KEYINPUT99), .A3(new_n567), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n554), .A2(new_n555), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT99), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n569), .A2(new_n570), .A3(new_n564), .A4(new_n548), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n572), .A2(new_n476), .B1(KEYINPUT41), .B2(new_n541), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n477), .A2(new_n479), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(new_n572), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n538), .A2(new_n539), .ZN(new_n576));
  XNOR2_X1  g375(.A(G134gat), .B(G162gat), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n578), .B1(new_n575), .B2(new_n576), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n544), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n581), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n583), .A2(new_n543), .A3(new_n579), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n521), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n556), .A2(new_n565), .A3(KEYINPUT101), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT101), .B1(new_n556), .B2(new_n565), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n586), .B(new_n567), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n568), .A2(new_n521), .A3(new_n571), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G230gat), .A2(G233gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT103), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT104), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n591), .A2(KEYINPUT104), .A3(new_n593), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT10), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n589), .A2(new_n590), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n511), .A2(KEYINPUT10), .A3(new_n520), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT102), .B1(new_n572), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT102), .ZN(new_n604));
  AOI211_X1 g403(.A(new_n604), .B(new_n601), .C1(new_n568), .C2(new_n571), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n600), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n593), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(G176gat), .B(G204gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  NAND3_X1  g410(.A1(new_n598), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT105), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n598), .A2(KEYINPUT105), .A3(new_n608), .A4(new_n611), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n608), .A2(new_n594), .ZN(new_n617));
  INV_X1    g416(.A(new_n611), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NOR3_X1   g419(.A1(new_n537), .A2(new_n585), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n505), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n622), .A2(new_n434), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(new_n453), .ZN(G1324gat));
  NOR2_X1   g423(.A1(new_n622), .A2(new_n437), .ZN(new_n625));
  XOR2_X1   g424(.A(KEYINPUT16), .B(G8gat), .Z(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT42), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n625), .A2(KEYINPUT42), .A3(new_n626), .ZN(new_n630));
  OAI21_X1  g429(.A(G8gat), .B1(new_n622), .B2(new_n437), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(G1325gat));
  AND2_X1   g431(.A1(new_n428), .A2(new_n440), .ZN(new_n633));
  OAI21_X1  g432(.A(G15gat), .B1(new_n622), .B2(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n424), .A2(new_n427), .ZN(new_n635));
  INV_X1    g434(.A(G15gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n634), .B1(new_n622), .B2(new_n637), .ZN(G1326gat));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n446), .ZN(new_n639));
  XOR2_X1   g438(.A(KEYINPUT43), .B(G22gat), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(G1327gat));
  NAND2_X1  g440(.A1(new_n441), .A2(new_n442), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n642), .A2(new_n444), .A3(new_n392), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n450), .A2(new_n448), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n620), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n537), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n585), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n645), .A2(new_n503), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n434), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(new_n464), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT45), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n428), .A2(new_n392), .A3(new_n439), .A4(new_n440), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n644), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n585), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n647), .A2(new_n504), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n648), .A2(new_n658), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n659), .B(new_n660), .C1(new_n451), .C2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(G29gat), .B1(new_n663), .B2(new_n434), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n652), .A2(new_n653), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n654), .A2(new_n664), .A3(new_n665), .ZN(G1328gat));
  NAND3_X1  g465(.A1(new_n650), .A2(new_n465), .A3(new_n305), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n667), .A2(KEYINPUT46), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(KEYINPUT46), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n663), .A2(KEYINPUT106), .A3(new_n437), .ZN(new_n670));
  OAI21_X1  g469(.A(KEYINPUT106), .B1(new_n663), .B2(new_n437), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(G36gat), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n668), .B(new_n669), .C1(new_n670), .C2(new_n672), .ZN(G1329gat));
  NAND4_X1  g472(.A1(new_n645), .A2(new_n503), .A3(new_n635), .A4(new_n649), .ZN(new_n674));
  INV_X1    g473(.A(G43gat), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(KEYINPUT47), .ZN(new_n678));
  INV_X1    g477(.A(new_n633), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(G43gat), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n676), .B(new_n678), .C1(new_n663), .C2(new_n680), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n677), .A2(KEYINPUT47), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1330gat));
  NOR2_X1   g482(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n446), .A2(G50gat), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n684), .B1(new_n650), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(G50gat), .B1(new_n663), .B2(new_n446), .ZN(new_n687));
  NAND2_X1  g486(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n686), .B2(new_n687), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(G1331gat));
  NOR4_X1   g490(.A1(new_n537), .A2(new_n646), .A3(new_n503), .A4(new_n585), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n656), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(new_n434), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(new_n515), .ZN(G1332gat));
  XNOR2_X1  g494(.A(new_n437), .B(KEYINPUT109), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n698));
  AND2_X1   g497(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n700), .B1(new_n697), .B2(new_n698), .ZN(G1333gat));
  OAI21_X1  g500(.A(G71gat), .B1(new_n693), .B2(new_n633), .ZN(new_n702));
  INV_X1    g501(.A(G71gat), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n635), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n693), .B2(new_n704), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g505(.A1(new_n693), .A2(new_n446), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(G78gat), .Z(G1335gat));
  INV_X1    g507(.A(new_n537), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(new_n503), .A3(new_n646), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n659), .B(new_n710), .C1(new_n451), .C2(new_n662), .ZN(new_n711));
  OAI21_X1  g510(.A(G85gat), .B1(new_n711), .B2(new_n434), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT51), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n709), .A2(new_n503), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n713), .B1(new_n657), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n648), .B1(new_n655), .B2(new_n644), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(KEYINPUT51), .A3(new_n714), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n651), .A2(new_n546), .A3(new_n620), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT110), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n712), .B1(new_n720), .B2(new_n722), .ZN(G1336gat));
  OAI21_X1  g522(.A(G92gat), .B1(new_n711), .B2(new_n437), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n696), .A2(G92gat), .A3(new_n646), .ZN(new_n725));
  INV_X1    g524(.A(new_n718), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT51), .B1(new_n717), .B2(new_n714), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n719), .A2(KEYINPUT111), .A3(new_n725), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n724), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT52), .ZN(new_n733));
  OAI21_X1  g532(.A(G92gat), .B1(new_n711), .B2(new_n696), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT52), .B1(new_n719), .B2(new_n725), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n735), .B1(new_n734), .B2(new_n736), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n733), .B1(new_n737), .B2(new_n738), .ZN(G1337gat));
  OAI21_X1  g538(.A(G99gat), .B1(new_n711), .B2(new_n633), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n635), .A2(new_n557), .A3(new_n620), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n720), .B2(new_n741), .ZN(G1338gat));
  OAI21_X1  g541(.A(G106gat), .B1(new_n711), .B2(new_n446), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n719), .A2(new_n558), .A3(new_n231), .A4(new_n620), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n745), .A2(new_n747), .A3(KEYINPUT53), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT53), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n743), .B(new_n744), .C1(new_n746), .C2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(G1339gat));
  NOR4_X1   g550(.A1(new_n537), .A2(new_n503), .A3(new_n585), .A4(new_n620), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT54), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n753), .B1(new_n606), .B2(new_n607), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n607), .B2(new_n606), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n606), .A2(new_n753), .A3(new_n607), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n756), .A2(KEYINPUT114), .A3(new_n618), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT114), .B1(new_n756), .B2(new_n618), .ZN(new_n758));
  OAI211_X1 g557(.A(KEYINPUT55), .B(new_n755), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n759), .A2(new_n616), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n755), .B1(new_n757), .B2(new_n758), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n490), .A2(new_n491), .A3(new_n489), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n481), .B1(new_n480), .B2(new_n485), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n498), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AND4_X1   g565(.A1(new_n502), .A2(new_n582), .A3(new_n584), .A4(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n760), .A2(new_n763), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n502), .A2(new_n766), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n769), .B1(new_n616), .B2(new_n619), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n759), .A2(new_n503), .A3(new_n616), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(new_n763), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n768), .B1(new_n772), .B2(new_n585), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n752), .B1(new_n773), .B2(new_n537), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(new_n434), .ZN(new_n775));
  INV_X1    g574(.A(new_n447), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n775), .A2(new_n776), .A3(new_n696), .ZN(new_n777));
  AOI21_X1  g576(.A(G113gat), .B1(new_n777), .B2(new_n503), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n763), .A2(new_n503), .A3(new_n616), .A4(new_n759), .ZN(new_n779));
  INV_X1    g578(.A(new_n770), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n585), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n760), .A2(new_n763), .A3(new_n767), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n537), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n752), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n446), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT115), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n696), .A2(new_n651), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(new_n635), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n504), .A2(new_n312), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n778), .B1(new_n790), .B2(new_n791), .ZN(G1340gat));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n314), .A3(new_n620), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(new_n620), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(new_n795), .A3(G120gat), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n795), .B1(new_n794), .B2(G120gat), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n793), .B1(new_n797), .B2(new_n798), .ZN(G1341gat));
  OAI21_X1  g598(.A(G127gat), .B1(new_n789), .B2(new_n537), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n777), .A2(new_n526), .A3(new_n709), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(G1342gat));
  OAI21_X1  g601(.A(G134gat), .B1(new_n789), .B2(new_n648), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n305), .A2(new_n648), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n775), .A2(new_n306), .A3(new_n776), .A4(new_n804), .ZN(new_n805));
  XOR2_X1   g604(.A(new_n805), .B(KEYINPUT56), .Z(new_n806));
  NAND2_X1  g605(.A1(new_n803), .A2(new_n806), .ZN(G1343gat));
  NAND2_X1  g606(.A1(new_n633), .A2(new_n788), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n446), .B1(new_n783), .B2(new_n784), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n810), .B1(new_n811), .B2(KEYINPUT57), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813));
  OAI211_X1 g612(.A(KEYINPUT117), .B(new_n813), .C1(new_n774), .C2(new_n446), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n446), .A2(new_n813), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n761), .A2(KEYINPUT118), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n819), .B(new_n755), .C1(new_n757), .C2(new_n758), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(new_n762), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT119), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n818), .A2(new_n823), .A3(new_n762), .A4(new_n820), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n822), .A2(new_n771), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n585), .B1(new_n825), .B2(new_n780), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n537), .B1(new_n826), .B2(new_n782), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n817), .B1(new_n827), .B2(new_n784), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n809), .B1(new_n815), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(G141gat), .B1(new_n829), .B2(new_n504), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT58), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n428), .A2(new_n231), .A3(new_n440), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n775), .A2(new_n696), .A3(new_n832), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n833), .A2(G141gat), .A3(new_n504), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n830), .A2(new_n831), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n829), .A2(KEYINPUT120), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n838), .B(new_n809), .C1(new_n815), .C2(new_n828), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(new_n503), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n834), .B1(new_n840), .B2(G141gat), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n836), .B1(new_n841), .B2(new_n831), .ZN(G1344gat));
  AND2_X1   g641(.A1(new_n827), .A2(new_n784), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n813), .B1(new_n843), .B2(new_n446), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n785), .A2(new_n816), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT121), .ZN(new_n846));
  AOI211_X1 g645(.A(new_n646), .B(new_n808), .C1(new_n844), .C2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(G148gat), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT59), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n837), .ZN(new_n850));
  INV_X1    g649(.A(new_n839), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n850), .A2(new_n851), .A3(new_n646), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n848), .A2(KEYINPUT59), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n849), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n775), .A2(new_n832), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n855), .A2(new_n848), .A3(new_n620), .A4(new_n696), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(G1345gat));
  INV_X1    g656(.A(KEYINPUT123), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n837), .A2(new_n709), .A3(new_n839), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(G155gat), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT122), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n855), .A2(new_n861), .A3(new_n709), .A4(new_n696), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT122), .B1(new_n833), .B2(new_n537), .ZN(new_n863));
  AOI21_X1  g662(.A(G155gat), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n858), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  AOI211_X1 g665(.A(KEYINPUT123), .B(new_n864), .C1(new_n859), .C2(G155gat), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(G1346gat));
  NAND3_X1  g667(.A1(new_n855), .A2(new_n215), .A3(new_n804), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n850), .A2(new_n851), .A3(new_n648), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(new_n215), .ZN(G1347gat));
  NOR2_X1   g670(.A1(new_n651), .A2(new_n437), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n787), .A2(new_n635), .A3(new_n872), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n873), .A2(new_n239), .A3(new_n504), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n696), .A2(new_n651), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n785), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n876), .A2(new_n776), .ZN(new_n877));
  AOI21_X1  g676(.A(G169gat), .B1(new_n877), .B2(new_n503), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n874), .A2(new_n878), .ZN(G1348gat));
  OAI21_X1  g678(.A(G176gat), .B1(new_n873), .B2(new_n646), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n877), .A2(new_n240), .A3(new_n620), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n882), .B(KEYINPUT124), .Z(G1349gat));
  OAI21_X1  g682(.A(G183gat), .B1(new_n873), .B2(new_n537), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n877), .A2(new_n246), .A3(new_n709), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g686(.A1(new_n877), .A2(new_n251), .A3(new_n585), .ZN(new_n888));
  OAI21_X1  g687(.A(G190gat), .B1(new_n873), .B2(new_n648), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n889), .A2(KEYINPUT61), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n889), .A2(KEYINPUT61), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(G1351gat));
  AND2_X1   g692(.A1(new_n876), .A2(new_n832), .ZN(new_n894));
  INV_X1    g693(.A(G197gat), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n895), .A3(new_n503), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n896), .B(KEYINPUT125), .Z(new_n897));
  NAND2_X1  g696(.A1(new_n633), .A2(new_n872), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n898), .B1(new_n844), .B2(new_n846), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n895), .B1(new_n899), .B2(new_n503), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n897), .A2(new_n900), .ZN(G1352gat));
  INV_X1    g700(.A(G204gat), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n646), .B1(new_n844), .B2(new_n846), .ZN(new_n903));
  INV_X1    g702(.A(new_n898), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n894), .A2(new_n902), .A3(new_n620), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT62), .ZN(new_n907));
  OR3_X1    g706(.A1(new_n905), .A2(new_n907), .A3(KEYINPUT126), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT126), .B1(new_n905), .B2(new_n907), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1353gat));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n203), .A3(new_n709), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n899), .A2(new_n709), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n912), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT63), .B1(new_n912), .B2(G211gat), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(G1354gat));
  AOI21_X1  g714(.A(G218gat), .B1(new_n894), .B2(new_n585), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT127), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n648), .A2(new_n204), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n899), .B2(new_n918), .ZN(G1355gat));
endmodule


