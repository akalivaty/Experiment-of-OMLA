//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n438, new_n439, new_n446, new_n451, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  OR2_X1    g012(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g013(.A1(new_n436), .A2(new_n437), .ZN(new_n439));
  NAND2_X1  g014(.A1(new_n438), .A2(new_n439), .ZN(G220));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g016(.A(G69), .ZN(G235));
  INV_X1    g017(.A(G120), .ZN(G236));
  XNOR2_X1  g018(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g019(.A(G108), .ZN(G238));
  NAND4_X1  g020(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT67), .ZN(G158));
  NAND3_X1  g022(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g023(.A(G452), .Z(G391));
  AND2_X1   g024(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR3_X1   g029(.A1(G221), .A2(G218), .A3(G219), .ZN(new_n455));
  NAND3_X1  g030(.A1(new_n438), .A2(new_n455), .A3(new_n439), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT2), .ZN(new_n457));
  NOR4_X1   g032(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  AOI22_X1  g036(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n463), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT68), .B(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n463), .A2(new_n465), .A3(G137), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n466), .A2(new_n471), .ZN(G160));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(new_n465), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(G2105), .ZN(new_n477));
  AOI22_X1  g052(.A1(G124), .A2(new_n476), .B1(new_n477), .B2(G136), .ZN(new_n478));
  OAI221_X1 g053(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n465), .C2(G112), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n463), .A2(new_n465), .A3(new_n482), .A4(G138), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT70), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n463), .A2(new_n465), .A3(G138), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n482), .B1(new_n485), .B2(KEYINPUT69), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n463), .A2(new_n465), .A3(new_n487), .A4(G138), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n484), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(G138), .B1(new_n473), .B2(new_n474), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n468), .A2(KEYINPUT68), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT69), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n495), .A2(new_n488), .A3(new_n496), .A4(KEYINPUT4), .ZN(new_n497));
  AND2_X1   g072(.A1(G126), .A2(G2105), .ZN(new_n498));
  OR2_X1    g073(.A1(new_n468), .A2(G114), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n463), .A2(new_n498), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n489), .A2(new_n503), .ZN(G164));
  NAND2_X1  g079(.A1(KEYINPUT71), .A2(G651), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  XNOR2_X1  g081(.A(new_n505), .B(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT5), .B(G543), .ZN(new_n510));
  AOI21_X1  g085(.A(KEYINPUT6), .B1(KEYINPUT71), .B2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n505), .A2(new_n506), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n508), .A2(new_n509), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n515), .A2(new_n518), .ZN(G166));
  INV_X1    g094(.A(new_n513), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n520), .A2(G89), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n524));
  INV_X1    g099(.A(G51), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n523), .B(new_n524), .C1(new_n508), .C2(new_n525), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n521), .A2(new_n526), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  NAND2_X1  g103(.A1(G77), .A2(G543), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT5), .B(G543), .Z(new_n530));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n520), .A2(G90), .B1(new_n532), .B2(G651), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n507), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G52), .ZN(new_n535));
  AOI21_X1  g110(.A(KEYINPUT72), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n533), .A2(KEYINPUT72), .A3(new_n535), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(G171));
  NAND2_X1  g114(.A1(new_n534), .A2(G43), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(new_n517), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n520), .A2(G81), .ZN(new_n543));
  AND3_X1   g118(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  NAND3_X1  g124(.A1(new_n507), .A2(G53), .A3(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(KEYINPUT9), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT9), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n507), .A2(new_n552), .A3(G53), .A4(G543), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n513), .A2(KEYINPUT73), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n507), .A2(new_n556), .A3(new_n510), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n555), .A2(new_n557), .A3(G91), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n510), .A2(G65), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT74), .Z(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n554), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT75), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n554), .A2(new_n565), .A3(new_n558), .A4(new_n562), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  INV_X1    g144(.A(G166), .ZN(G303));
  NAND3_X1  g145(.A1(new_n555), .A2(new_n557), .A3(G87), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(KEYINPUT76), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n555), .A2(new_n557), .A3(new_n573), .A4(G87), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n510), .A2(G74), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n534), .A2(G49), .B1(G651), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(G288));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n530), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n534), .A2(G48), .B1(new_n581), .B2(G651), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n555), .A2(new_n557), .A3(G86), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G305));
  NAND2_X1  g159(.A1(new_n520), .A2(G85), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  XOR2_X1   g161(.A(KEYINPUT77), .B(G47), .Z(new_n587));
  OAI221_X1 g162(.A(new_n585), .B1(new_n517), .B2(new_n586), .C1(new_n508), .C2(new_n587), .ZN(G290));
  INV_X1    g163(.A(G868), .ZN(new_n589));
  NOR2_X1   g164(.A1(G171), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT78), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n555), .A2(new_n557), .A3(G92), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT79), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n530), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(G54), .A2(new_n534), .B1(new_n598), .B2(G651), .ZN(new_n599));
  AND3_X1   g174(.A1(new_n594), .A2(KEYINPUT80), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(KEYINPUT80), .B1(new_n594), .B2(new_n599), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n591), .B1(G868), .B2(new_n603), .ZN(G284));
  OAI21_X1  g179(.A(new_n591), .B1(G868), .B2(new_n603), .ZN(G321));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n567), .B2(G868), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(new_n567), .B2(G868), .ZN(G280));
  NOR2_X1   g183(.A1(new_n602), .A2(G559), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(G860), .B2(new_n603), .ZN(G148));
  NAND3_X1  g185(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(new_n589), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n609), .B2(new_n589), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n463), .A2(new_n469), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(KEYINPUT82), .B(KEYINPUT13), .Z(new_n618));
  XOR2_X1   g193(.A(new_n617), .B(new_n618), .Z(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n620), .A2(G2100), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT83), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n476), .A2(G123), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n477), .A2(G135), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n465), .A2(G111), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n626), .A2(KEYINPUT84), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(new_n626), .B2(KEYINPUT84), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n625), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(G2096), .ZN(new_n631));
  AOI22_X1  g206(.A1(new_n620), .A2(G2100), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n622), .B(new_n632), .C1(new_n631), .C2(new_n630), .ZN(G156));
  INV_X1    g208(.A(G14), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  INV_X1    g210(.A(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n635), .B(G2430), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(new_n638), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n640), .A2(new_n642), .A3(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT16), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  INV_X1    g222(.A(new_n645), .ZN(new_n648));
  NAND4_X1  g223(.A1(new_n648), .A2(new_n640), .A3(new_n642), .A4(KEYINPUT14), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n647), .B1(new_n646), .B2(new_n649), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n634), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT85), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n646), .A2(new_n649), .ZN(new_n658));
  INV_X1    g233(.A(new_n647), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(new_n650), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n657), .B1(new_n661), .B2(new_n654), .ZN(new_n662));
  AOI211_X1 g237(.A(KEYINPUT85), .B(new_n655), .C1(new_n660), .C2(new_n650), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n656), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G401));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2072), .B(G2078), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT18), .Z(new_n670));
  INV_X1    g245(.A(KEYINPUT86), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n668), .B1(new_n671), .B2(new_n667), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n671), .B2(new_n667), .ZN(new_n673));
  INV_X1    g248(.A(new_n666), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n667), .B(KEYINPUT17), .Z(new_n675));
  INV_X1    g250(.A(new_n668), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n673), .B(new_n674), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n675), .A2(new_n676), .A3(new_n666), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n670), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(new_n631), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT87), .B(G2100), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(G2096), .ZN(new_n683));
  INV_X1    g258(.A(new_n681), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT89), .Z(new_n688));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT88), .ZN(new_n690));
  XOR2_X1   g265(.A(G1956), .B(G2474), .Z(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1971), .B(G1976), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT19), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n694), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n690), .B2(new_n691), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n695), .B1(new_n692), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n696), .A2(new_n690), .A3(new_n691), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT20), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n688), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(G1991), .B(G1996), .Z(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n698), .A2(new_n700), .A3(new_n688), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n702), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n705), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n703), .B1(new_n707), .B2(new_n701), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1981), .B(G1986), .ZN(new_n709));
  AND3_X1   g284(.A1(new_n706), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n706), .B2(new_n708), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(G229));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G26), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT28), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n476), .A2(G128), .ZN(new_n717));
  OAI221_X1 g292(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n465), .C2(G116), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n477), .A2(G140), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n716), .B1(new_n720), .B2(G29), .ZN(new_n721));
  INV_X1    g296(.A(G2067), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(G21), .B(G286), .S(G16), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1966), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT91), .B(G16), .Z(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(G19), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n544), .B2(new_n727), .ZN(new_n729));
  AOI211_X1 g304(.A(new_n723), .B(new_n725), .C1(G1341), .C2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n726), .A2(G20), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT100), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT23), .Z(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G299), .B2(G16), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT101), .B(G1956), .Z(new_n736));
  OR2_X1    g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n714), .A2(G35), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G162), .B2(new_n714), .ZN(new_n739));
  INV_X1    g314(.A(G2090), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G11), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n744), .A2(KEYINPUT31), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(KEYINPUT31), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT30), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n747), .A2(G28), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n714), .B1(new_n747), .B2(G28), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n745), .B(new_n746), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n630), .B2(G29), .ZN(new_n751));
  INV_X1    g326(.A(G34), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n752), .A2(KEYINPUT24), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n752), .B2(KEYINPUT24), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(KEYINPUT94), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(KEYINPUT94), .B2(new_n754), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT95), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G29), .B2(G160), .ZN(new_n758));
  OAI221_X1 g333(.A(new_n751), .B1(new_n758), .B2(G2084), .C1(G1341), .C2(new_n729), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n714), .A2(G32), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n476), .A2(G129), .ZN(new_n761));
  NAND3_X1  g336(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT26), .Z(new_n763));
  AND2_X1   g338(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT97), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n477), .A2(G141), .B1(G105), .B2(new_n469), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n766), .A2(new_n761), .A3(new_n763), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(KEYINPUT97), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n760), .B1(new_n770), .B2(G29), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT27), .B(G1996), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n759), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n730), .A2(new_n737), .A3(new_n743), .A4(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n736), .B2(new_n735), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT102), .ZN(new_n777));
  NOR2_X1   g352(.A1(G4), .A2(G16), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n603), .B2(G16), .ZN(new_n779));
  INV_X1    g354(.A(G1348), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n758), .A2(G2084), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT96), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n771), .A2(new_n772), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n714), .A2(G33), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT25), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n477), .A2(G139), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n788), .B(new_n789), .C1(new_n465), .C2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n785), .B1(new_n791), .B2(G29), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G2072), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n783), .A2(new_n784), .A3(new_n793), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT98), .Z(new_n795));
  NOR2_X1   g370(.A1(G5), .A2(G16), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G171), .B2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1961), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n714), .A2(G27), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G164), .B2(new_n714), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G2078), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n795), .A2(new_n798), .A3(new_n801), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n776), .A2(new_n777), .A3(new_n781), .A4(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n776), .A2(new_n781), .A3(new_n802), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(KEYINPUT102), .ZN(new_n805));
  MUX2_X1   g380(.A(G6), .B(G305), .S(G16), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT92), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT32), .B(G1981), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  MUX2_X1   g384(.A(G23), .B(G288), .S(G16), .Z(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT33), .B(G1976), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n727), .A2(G22), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G166), .B2(new_n727), .ZN(new_n814));
  INV_X1    g389(.A(G1971), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n809), .A2(new_n812), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT34), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n809), .A2(new_n819), .A3(new_n812), .A4(new_n816), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n714), .A2(G25), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT90), .ZN(new_n822));
  AOI22_X1  g397(.A1(G119), .A2(new_n476), .B1(new_n477), .B2(G131), .ZN(new_n823));
  OAI221_X1 g398(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n465), .C2(G107), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n822), .B1(new_n825), .B2(G29), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT35), .B(G1991), .Z(new_n827));
  XOR2_X1   g402(.A(new_n826), .B(new_n827), .Z(new_n828));
  MUX2_X1   g403(.A(G24), .B(G290), .S(new_n727), .Z(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(G1986), .Z(new_n830));
  NAND4_X1  g405(.A1(new_n818), .A2(new_n820), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT36), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n832), .A2(KEYINPUT93), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n831), .B(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n832), .A2(KEYINPUT93), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n803), .A2(new_n805), .B1(new_n834), .B2(new_n835), .ZN(G311));
  NAND2_X1  g411(.A1(new_n805), .A2(new_n803), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n834), .A2(new_n835), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(G150));
  NAND2_X1  g414(.A1(new_n603), .A2(G559), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT38), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n507), .A2(G55), .A3(G543), .ZN(new_n842));
  INV_X1    g417(.A(G93), .ZN(new_n843));
  AOI22_X1  g418(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n844));
  OAI221_X1 g419(.A(new_n842), .B1(new_n513), .B2(new_n843), .C1(new_n517), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n611), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n611), .A2(new_n845), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n841), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT39), .ZN(new_n852));
  AOI21_X1  g427(.A(G860), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n852), .B2(new_n851), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n845), .A2(G860), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT37), .Z(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(G145));
  XNOR2_X1  g432(.A(G160), .B(KEYINPUT103), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(G162), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n630), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT105), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n791), .B2(KEYINPUT104), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(new_n861), .B2(new_n791), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n765), .B1(new_n764), .B2(new_n766), .ZN(new_n864));
  AND4_X1   g439(.A1(new_n765), .A2(new_n766), .A3(new_n761), .A4(new_n763), .ZN(new_n865));
  INV_X1    g440(.A(new_n720), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n720), .B1(new_n767), .B2(new_n769), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n867), .A2(new_n868), .A3(G164), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n489), .A2(new_n503), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n866), .B1(new_n864), .B2(new_n865), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n767), .A2(new_n769), .A3(new_n720), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n863), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(G164), .B1(new_n867), .B2(new_n868), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n871), .A2(new_n872), .A3(new_n870), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n862), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n617), .ZN(new_n878));
  AOI22_X1  g453(.A1(G130), .A2(new_n476), .B1(new_n477), .B2(G142), .ZN(new_n879));
  OAI221_X1 g454(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n465), .C2(G118), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n881), .A2(new_n824), .A3(new_n823), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n825), .A2(new_n880), .A3(new_n879), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n884), .B1(new_n882), .B2(new_n883), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n878), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n882), .A2(new_n883), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT106), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n617), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n874), .A2(new_n877), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n892), .B1(new_n874), .B2(new_n877), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n860), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT107), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n897), .B(new_n860), .C1(new_n893), .C2(new_n894), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n893), .A2(new_n894), .A3(new_n860), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n900), .A2(G37), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g478(.A(new_n609), .B(new_n849), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n594), .A2(new_n599), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n906), .A2(new_n567), .A3(KEYINPUT108), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT108), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n564), .A2(new_n908), .A3(new_n566), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n908), .B1(new_n564), .B2(new_n566), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n909), .A2(new_n910), .A3(new_n905), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n904), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n911), .B2(new_n907), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n910), .A2(new_n905), .ZN(new_n915));
  INV_X1    g490(.A(new_n909), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(G299), .A2(new_n908), .A3(new_n905), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(KEYINPUT41), .A3(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n914), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n912), .B1(new_n904), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT42), .ZN(new_n922));
  XNOR2_X1  g497(.A(G288), .B(G166), .ZN(new_n923));
  XNOR2_X1  g498(.A(G290), .B(G305), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n923), .B(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n926), .A2(KEYINPUT109), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n912), .B(new_n928), .C1(new_n904), .C2(new_n920), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n922), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n927), .B1(new_n922), .B2(new_n929), .ZN(new_n931));
  OAI21_X1  g506(.A(G868), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n845), .A2(new_n589), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(G295));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n933), .ZN(G331));
  OAI211_X1 g510(.A(new_n538), .B(new_n537), .C1(new_n847), .C2(new_n848), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n611), .A2(new_n845), .ZN(new_n937));
  INV_X1    g512(.A(new_n538), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n937), .B(new_n846), .C1(new_n938), .C2(new_n536), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(G286), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n936), .A2(new_n939), .A3(G168), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n914), .A2(new_n919), .A3(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n941), .A2(new_n917), .A3(new_n918), .A4(new_n942), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(G37), .B1(new_n946), .B2(new_n925), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n926), .A3(new_n945), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n947), .A2(new_n951), .A3(new_n948), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n953), .B(new_n954), .ZN(G397));
  INV_X1    g530(.A(G1384), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(new_n489), .B2(new_n503), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(G160), .A2(G40), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G1996), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(new_n770), .ZN(new_n964));
  XOR2_X1   g539(.A(new_n961), .B(KEYINPUT110), .Z(new_n965));
  NAND2_X1  g540(.A1(new_n866), .A2(new_n722), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n720), .A2(G2067), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n770), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n968), .B1(new_n969), .B2(new_n962), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n964), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n825), .B(new_n827), .Z(new_n972));
  NAND2_X1  g547(.A1(new_n965), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(G290), .B(G1986), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n974), .B1(new_n961), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n977));
  INV_X1    g552(.A(G8), .ZN(new_n978));
  NOR2_X1   g553(.A1(G168), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n957), .A2(KEYINPUT50), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n982), .B(new_n956), .C1(new_n489), .C2(new_n503), .ZN(new_n983));
  INV_X1    g558(.A(new_n960), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n985), .A2(G2084), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n870), .A2(KEYINPUT116), .A3(KEYINPUT45), .A4(new_n956), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n960), .B1(new_n957), .B2(new_n958), .ZN(new_n988));
  OAI211_X1 g563(.A(KEYINPUT45), .B(new_n956), .C1(new_n489), .C2(new_n503), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n987), .A2(new_n988), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1966), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n986), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(G8), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n980), .B1(new_n996), .B2(KEYINPUT122), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n978), .B1(new_n986), .B2(new_n994), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT122), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n977), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n980), .A2(KEYINPUT51), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT121), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1002), .B1(new_n998), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n996), .A2(KEYINPUT121), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n1004), .A2(new_n1005), .B1(new_n995), .B2(new_n979), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1001), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n960), .B1(new_n957), .B2(KEYINPUT50), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT120), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n983), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1009), .B1(new_n1008), .B2(new_n983), .ZN(new_n1011));
  XOR2_X1   g586(.A(KEYINPUT123), .B(G1961), .Z(new_n1012));
  NOR3_X1   g587(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G2078), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n988), .A2(new_n1014), .A3(new_n989), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(G2078), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n987), .A2(new_n988), .A3(new_n991), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(G171), .B1(new_n1013), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT124), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n985), .A2(KEYINPUT120), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1008), .A2(new_n1009), .A3(new_n983), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1012), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1027), .A2(new_n1019), .A3(new_n1017), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT125), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n988), .A2(new_n1030), .A3(new_n989), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1015), .A2(new_n1031), .A3(KEYINPUT53), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1015), .B1(new_n1031), .B2(KEYINPUT53), .ZN(new_n1033));
  OAI211_X1 g608(.A(G301), .B(new_n1027), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1023), .A2(new_n1029), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n563), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n1040), .B(KEYINPUT118), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1039), .B(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G1956), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n985), .A2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT56), .B(G2072), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n988), .A2(new_n989), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1042), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1044), .A2(new_n1042), .A3(new_n1046), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(new_n602), .ZN(new_n1050));
  INV_X1    g625(.A(new_n957), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1051), .A2(new_n722), .A3(new_n984), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1052), .B(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1024), .A2(new_n780), .A3(new_n1025), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1047), .B1(new_n1050), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT61), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n1049), .B2(new_n1047), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n988), .A2(new_n962), .A3(new_n989), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n870), .A2(new_n956), .A3(new_n984), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT58), .B(G1341), .Z(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT59), .B1(new_n1064), .B2(new_n544), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n1066));
  AOI211_X1 g641(.A(new_n1066), .B(new_n611), .C1(new_n1060), .C2(new_n1063), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1042), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1071), .A2(new_n1048), .A3(KEYINPUT61), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1059), .A2(new_n1068), .A3(new_n1072), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1010), .A2(new_n1011), .A3(G1348), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1052), .B(KEYINPUT119), .ZN(new_n1075));
  OAI211_X1 g650(.A(KEYINPUT60), .B(new_n603), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n603), .A2(KEYINPUT60), .ZN(new_n1077));
  OR3_X1    g652(.A1(new_n600), .A2(new_n601), .A3(KEYINPUT60), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1077), .A2(new_n1054), .A3(new_n1055), .A4(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1057), .B1(new_n1073), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT111), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1008), .A2(new_n740), .A3(new_n983), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(G1971), .B1(new_n988), .B2(new_n989), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1082), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(G303), .A2(G8), .ZN(new_n1087));
  XNOR2_X1  g662(.A(new_n1087), .B(KEYINPUT55), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n959), .A2(new_n984), .A3(new_n989), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n815), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1091), .A2(KEYINPUT111), .A3(new_n1083), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1086), .A2(G8), .A3(new_n1089), .A4(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n978), .B1(new_n1051), .B2(new_n984), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n581), .A2(G651), .ZN(new_n1095));
  INV_X1    g670(.A(G48), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1095), .B1(new_n1096), .B2(new_n508), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT113), .B(G86), .Z(new_n1098));
  NOR2_X1   g673(.A1(new_n513), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(G1981), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1981), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n582), .A2(new_n1101), .A3(new_n583), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT49), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1100), .A2(KEYINPUT49), .A3(new_n1102), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1094), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n577), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1108), .B1(new_n572), .B2(new_n574), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT112), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(new_n1110), .A3(G1976), .ZN(new_n1111));
  INV_X1    g686(.A(G1976), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT112), .B1(G288), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1094), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT52), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1109), .B2(G1976), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1107), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  NOR3_X1   g692(.A1(G288), .A2(KEYINPUT112), .A3(new_n1112), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1110), .B1(new_n1109), .B2(G1976), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1115), .B1(new_n1120), .B2(new_n1094), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(G8), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n1088), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1093), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1028), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1036), .B1(new_n1126), .B2(G301), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1027), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(G171), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1125), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1037), .A2(new_n1081), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1125), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1029), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT124), .B1(new_n1028), .B2(G171), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1132), .B(new_n1133), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1007), .B1(new_n1131), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n998), .A2(G168), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT63), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1086), .A2(G8), .A3(new_n1092), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n1088), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1140), .A2(new_n1093), .A3(new_n1122), .A4(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1139), .B1(new_n1125), .B2(new_n1138), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1107), .A2(new_n1112), .A3(new_n1109), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1102), .B(KEYINPUT114), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1094), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1148), .B1(new_n1149), .B2(new_n1093), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT115), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1148), .B(KEYINPUT115), .C1(new_n1149), .C2(new_n1093), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1132), .B(KEYINPUT62), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1001), .A2(new_n1006), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1145), .B(new_n1154), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n976), .B1(new_n1137), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n965), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n971), .A2(new_n827), .A3(new_n824), .A4(new_n823), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1159), .B1(new_n1160), .B2(new_n966), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n963), .B(KEYINPUT46), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n968), .A2(new_n969), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n1159), .B2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g739(.A(new_n1164), .B(KEYINPUT47), .Z(new_n1165));
  INV_X1    g740(.A(new_n974), .ZN(new_n1166));
  NOR2_X1   g741(.A1(G290), .A2(G1986), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n961), .A2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT48), .ZN(new_n1169));
  AOI211_X1 g744(.A(new_n1161), .B(new_n1165), .C1(new_n1166), .C2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1158), .A2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g746(.A(KEYINPUT126), .ZN(new_n1173));
  AND3_X1   g747(.A1(new_n682), .A2(new_n685), .A3(G319), .ZN(new_n1174));
  AND3_X1   g748(.A1(new_n664), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g749(.A(new_n1173), .B1(new_n664), .B2(new_n1174), .ZN(new_n1176));
  OAI21_X1  g750(.A(new_n712), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g751(.A(new_n1177), .B1(new_n899), .B2(new_n901), .ZN(new_n1178));
  AOI21_X1  g752(.A(KEYINPUT127), .B1(new_n953), .B2(new_n1178), .ZN(new_n1179));
  AND3_X1   g753(.A1(new_n947), .A2(new_n951), .A3(new_n948), .ZN(new_n1180));
  AOI21_X1  g754(.A(new_n951), .B1(new_n947), .B2(new_n948), .ZN(new_n1181));
  OAI211_X1 g755(.A(new_n1178), .B(KEYINPUT127), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  INV_X1    g756(.A(new_n1182), .ZN(new_n1183));
  NOR2_X1   g757(.A1(new_n1179), .A2(new_n1183), .ZN(G308));
  NAND2_X1  g758(.A1(new_n953), .A2(new_n1178), .ZN(G225));
endmodule


