//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n841, new_n842,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT26), .ZN(new_n205));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT26), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n202), .B(new_n205), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT27), .B(G183gat), .ZN(new_n212));
  INV_X1    g011(.A(G190gat), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT28), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G183gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT27), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT27), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G183gat), .ZN(new_n218));
  AND4_X1   g017(.A1(KEYINPUT28), .A2(new_n216), .A3(new_n218), .A4(new_n213), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n211), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n206), .B1(new_n202), .B2(KEYINPUT24), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(new_n203), .A3(new_n204), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n221), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n215), .A2(new_n213), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n226), .A2(KEYINPUT24), .A3(new_n202), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT25), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n221), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n224), .A2(new_n222), .ZN(new_n230));
  AND4_X1   g029(.A1(KEYINPUT25), .A2(new_n229), .A3(new_n230), .A4(new_n227), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n220), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT73), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT29), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n220), .B(KEYINPUT73), .C1(new_n228), .C2(new_n231), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G226gat), .A2(G233gat), .ZN(new_n238));
  XOR2_X1   g037(.A(new_n238), .B(KEYINPUT72), .Z(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G197gat), .B(G204gat), .ZN(new_n242));
  AND2_X1   g041(.A1(G211gat), .A2(G218gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n242), .B1(KEYINPUT22), .B2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(G211gat), .A2(G218gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n244), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n220), .A2(KEYINPUT65), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n216), .A2(new_n218), .A3(new_n213), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT28), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n212), .A2(KEYINPUT28), .A3(new_n213), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n254), .A3(new_n211), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n248), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT64), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n257), .B1(new_n228), .B2(new_n231), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n225), .A2(KEYINPUT25), .A3(new_n227), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n229), .A2(new_n230), .A3(new_n227), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT25), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n262), .A3(KEYINPUT64), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n256), .A2(new_n258), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(new_n239), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n241), .A2(new_n247), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n234), .A2(new_n236), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n239), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n239), .A2(KEYINPUT29), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n244), .A2(new_n246), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n244), .A2(new_n246), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n268), .A2(new_n270), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G8gat), .B(G36gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(G64gat), .B(G92gat), .ZN(new_n276));
  XOR2_X1   g075(.A(new_n275), .B(new_n276), .Z(new_n277));
  AND3_X1   g076(.A1(new_n266), .A2(new_n274), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n277), .B1(new_n266), .B2(new_n274), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT30), .ZN(new_n280));
  OR3_X1    g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n274), .ZN(new_n282));
  INV_X1    g081(.A(new_n277), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n282), .A2(KEYINPUT30), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n287));
  XOR2_X1   g086(.A(KEYINPUT74), .B(KEYINPUT2), .Z(new_n288));
  XOR2_X1   g087(.A(G141gat), .B(G148gat), .Z(new_n289));
  INV_X1    g088(.A(G162gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G155gat), .ZN(new_n291));
  INV_X1    g090(.A(G155gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G162gat), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n288), .A2(new_n289), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT78), .ZN(new_n296));
  INV_X1    g095(.A(G141gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(G148gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  XOR2_X1   g098(.A(KEYINPUT75), .B(G141gat), .Z(new_n300));
  INV_X1    g099(.A(G148gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n292), .A2(G162gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n290), .A2(G155gat), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT76), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT76), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n291), .A2(new_n293), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  AND2_X1   g107(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n310));
  OAI21_X1  g109(.A(G155gat), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT2), .ZN(new_n312));
  AND4_X1   g111(.A1(new_n296), .A2(new_n302), .A3(new_n308), .A4(new_n312), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n305), .A2(new_n307), .B1(new_n311), .B2(KEYINPUT2), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n296), .B1(new_n314), .B2(new_n302), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n295), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G113gat), .ZN(new_n317));
  INV_X1    g116(.A(G120gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT68), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n317), .A2(new_n318), .B1(new_n319), .B2(KEYINPUT1), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(new_n319), .B2(KEYINPUT1), .ZN(new_n321));
  XOR2_X1   g120(.A(G127gat), .B(G134gat), .Z(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  XOR2_X1   g122(.A(KEYINPUT67), .B(G113gat), .Z(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G120gat), .ZN(new_n325));
  XOR2_X1   g124(.A(KEYINPUT66), .B(G127gat), .Z(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G134gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(G127gat), .A2(G134gat), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT1), .B1(new_n317), .B2(new_n318), .ZN(new_n329));
  NAND2_X1  g128(.A1(G113gat), .A2(G120gat), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n323), .A2(new_n325), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n295), .B(new_n332), .C1(new_n313), .C2(new_n315), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G225gat), .A2(G233gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n287), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n306), .B1(new_n291), .B2(new_n293), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n291), .A2(new_n293), .A3(new_n306), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n312), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT75), .B(G141gat), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n298), .B1(new_n343), .B2(G148gat), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT78), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n314), .A2(new_n296), .A3(new_n302), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n294), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT79), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .A4(new_n332), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n333), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n316), .A2(KEYINPUT3), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n337), .B(new_n350), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n335), .A2(KEYINPUT4), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n345), .A2(new_n346), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n356), .A2(new_n349), .A3(new_n295), .A4(new_n332), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n355), .A2(KEYINPUT79), .A3(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n339), .B1(new_n354), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT0), .ZN(new_n361));
  XNOR2_X1  g160(.A(G57gat), .B(G85gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  AOI21_X1  g162(.A(new_n332), .B1(new_n316), .B2(KEYINPUT3), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n351), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n338), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n335), .A2(KEYINPUT80), .A3(KEYINPUT4), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT80), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n355), .A2(new_n368), .A3(new_n357), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n366), .A2(new_n287), .A3(new_n367), .A4(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n359), .A2(new_n363), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT6), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n363), .B1(new_n359), .B2(new_n370), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI211_X1 g174(.A(new_n372), .B(new_n363), .C1(new_n359), .C2(new_n370), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n286), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G78gat), .B(G106gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n378), .B(G22gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n316), .A2(new_n235), .A3(new_n247), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n316), .A2(KEYINPUT3), .ZN(new_n382));
  NAND2_X1  g181(.A1(G228gat), .A2(G233gat), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n385), .B(new_n273), .C1(new_n353), .C2(KEYINPUT29), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT29), .B1(new_n347), .B2(new_n351), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT81), .B1(new_n387), .B2(new_n247), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n384), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n387), .A2(new_n247), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n247), .A2(new_n235), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT3), .B1(new_n391), .B2(KEYINPUT82), .ZN(new_n392));
  OR3_X1    g191(.A1(new_n273), .A2(KEYINPUT82), .A3(KEYINPUT29), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n347), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI211_X1 g193(.A(G228gat), .B(G233gat), .C1(new_n390), .C2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT31), .B(G50gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n389), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n397), .B1(new_n389), .B2(new_n395), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n380), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n389), .A2(new_n395), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n396), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n389), .A2(new_n395), .A3(new_n397), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n402), .A2(new_n379), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n258), .A2(new_n263), .ZN(new_n406));
  AOI211_X1 g205(.A(KEYINPUT65), .B(new_n210), .C1(new_n251), .C2(new_n252), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n254), .B1(new_n253), .B2(new_n211), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n332), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(G227gat), .ZN(new_n411));
  INV_X1    g210(.A(G233gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n256), .A2(new_n333), .A3(new_n258), .A4(new_n263), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n410), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT32), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  XOR2_X1   g217(.A(G15gat), .B(G43gat), .Z(new_n419));
  XNOR2_X1  g218(.A(G71gat), .B(G99gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n416), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n421), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n415), .B(KEYINPUT32), .C1(new_n417), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT71), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT71), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n422), .A2(new_n427), .A3(new_n424), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n414), .ZN(new_n429));
  INV_X1    g228(.A(new_n413), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n431), .B1(new_n429), .B2(new_n430), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n426), .A2(new_n428), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT36), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n434), .A2(new_n427), .A3(new_n422), .A4(new_n424), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT70), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n435), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n425), .A2(new_n434), .A3(new_n440), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(KEYINPUT36), .A3(new_n443), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n377), .A2(new_n405), .B1(new_n439), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n241), .A2(new_n273), .A3(new_n265), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n268), .A2(new_n270), .A3(new_n247), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT85), .A4(KEYINPUT37), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT38), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT37), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n239), .A2(new_n267), .B1(new_n264), .B2(new_n269), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n451), .B1(new_n452), .B2(new_n247), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT85), .B1(new_n453), .B2(new_n446), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n283), .B1(new_n282), .B2(KEYINPUT37), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n278), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n374), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n459), .A2(new_n372), .A3(new_n371), .ZN(new_n460));
  INV_X1    g259(.A(new_n376), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n451), .B1(new_n266), .B2(new_n274), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT38), .B1(new_n456), .B2(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n458), .A2(new_n460), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n465));
  NOR3_X1   g264(.A1(new_n465), .A2(new_n374), .A3(new_n284), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n382), .A2(new_n365), .A3(new_n333), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n369), .A2(new_n467), .A3(new_n367), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n338), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n470), .A2(KEYINPUT39), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  XOR2_X1   g271(.A(KEYINPUT83), .B(KEYINPUT39), .Z(new_n473));
  NAND3_X1  g272(.A1(new_n468), .A2(new_n338), .A3(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n472), .A2(KEYINPUT40), .A3(new_n363), .A4(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT84), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n474), .A2(new_n363), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n478), .A2(KEYINPUT84), .A3(KEYINPUT40), .A4(new_n472), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n472), .A2(new_n363), .A3(new_n474), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT40), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n466), .A2(new_n477), .A3(new_n479), .A4(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n405), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n464), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n445), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n442), .A2(new_n400), .A3(new_n404), .A4(new_n443), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT35), .B1(new_n377), .B2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT86), .B(KEYINPUT35), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n400), .A2(new_n404), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n436), .A2(new_n438), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n460), .A2(new_n461), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .A4(new_n286), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n486), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G113gat), .B(G141gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(KEYINPUT87), .B(G197gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  XOR2_X1   g297(.A(KEYINPUT11), .B(G169gat), .Z(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT12), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT89), .ZN(new_n502));
  INV_X1    g301(.A(G43gat), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n502), .B1(new_n503), .B2(G50gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(G50gat), .ZN(new_n505));
  INV_X1    g304(.A(G50gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n506), .A2(KEYINPUT89), .A3(G43gat), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT15), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT90), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n506), .A2(G43gat), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n505), .A2(new_n513), .A3(KEYINPUT15), .ZN(new_n514));
  INV_X1    g313(.A(G29gat), .ZN(new_n515));
  INV_X1    g314(.A(G36gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT14), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT14), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(G29gat), .B2(G36gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n515), .A2(new_n516), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n514), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n508), .A2(KEYINPUT90), .A3(new_n509), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n512), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT88), .ZN(new_n525));
  OAI22_X1  g324(.A1(new_n520), .A2(new_n525), .B1(new_n515), .B2(new_n516), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT88), .B1(new_n517), .B2(new_n519), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n514), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT17), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n524), .A2(new_n531), .A3(new_n528), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(KEYINPUT91), .B(G1gat), .Z(new_n534));
  OR2_X1    g333(.A1(G15gat), .A2(G22gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(G15gat), .A2(G22gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(new_n537), .A3(KEYINPUT16), .ZN(new_n538));
  NAND2_X1  g337(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n539));
  OR2_X1    g338(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n535), .A2(G1gat), .A3(new_n536), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(G15gat), .A2(G22gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(G15gat), .A2(G22gat), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT16), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT91), .B(G1gat), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n540), .B(new_n541), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n539), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n542), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT93), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n542), .A2(new_n549), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n533), .A2(new_n551), .B1(new_n529), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G229gat), .A2(G233gat), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n554), .B(KEYINPUT94), .Z(new_n555));
  AOI21_X1  g354(.A(KEYINPUT18), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT93), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n550), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n552), .A2(KEYINPUT93), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n524), .A2(new_n531), .A3(new_n528), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n531), .B1(new_n524), .B2(new_n528), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n558), .B(new_n559), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n529), .A2(new_n552), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n562), .A2(KEYINPUT18), .A3(new_n555), .A4(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n556), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT95), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n550), .A2(new_n524), .A3(new_n528), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n563), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n555), .B(KEYINPUT13), .Z(new_n570));
  NAND3_X1  g369(.A1(new_n529), .A2(new_n552), .A3(KEYINPUT95), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT96), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT96), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n569), .A2(new_n574), .A3(new_n570), .A4(new_n571), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n501), .B1(new_n566), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n562), .A2(new_n555), .A3(new_n563), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT18), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AND4_X1   g379(.A1(new_n576), .A2(new_n580), .A3(new_n564), .A4(new_n501), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(G71gat), .ZN(new_n584));
  INV_X1    g383(.A(G78gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G71gat), .A2(G78gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT97), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n586), .A2(KEYINPUT97), .A3(new_n587), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT9), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  OR2_X1    g392(.A1(G57gat), .A2(G64gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(G57gat), .A2(G64gat), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n590), .A2(new_n591), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n594), .A2(new_n595), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n586), .A2(new_n587), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n598), .A2(new_n599), .A3(KEYINPUT97), .A4(new_n593), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(G231gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n602), .A2(new_n412), .ZN(new_n603));
  OR3_X1    g402(.A1(new_n601), .A2(KEYINPUT21), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n603), .B1(new_n601), .B2(KEYINPUT21), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(G127gat), .ZN(new_n607));
  INV_X1    g406(.A(new_n601), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT21), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n550), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT98), .Z(new_n611));
  OR2_X1    g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n607), .A2(new_n611), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(new_n292), .ZN(new_n615));
  XOR2_X1   g414(.A(G183gat), .B(G211gat), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n612), .A2(new_n613), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n617), .B1(new_n612), .B2(new_n613), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G85gat), .A2(G92gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT7), .ZN(new_n623));
  INV_X1    g422(.A(G99gat), .ZN(new_n624));
  INV_X1    g423(.A(G106gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G99gat), .A2(G106gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(G85gat), .ZN(new_n629));
  INV_X1    g428(.A(G92gat), .ZN(new_n630));
  AOI22_X1  g429(.A1(KEYINPUT8), .A2(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n623), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n628), .B1(new_n623), .B2(new_n631), .ZN(new_n633));
  OAI22_X1  g432(.A1(new_n560), .A2(new_n561), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT41), .ZN(new_n637));
  INV_X1    g436(.A(G232gat), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n637), .A2(new_n638), .A3(new_n412), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n632), .A2(new_n633), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n639), .B1(new_n529), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n641), .B1(new_n634), .B2(new_n635), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n643));
  XNOR2_X1  g442(.A(G190gat), .B(G218gat), .ZN(new_n644));
  OAI22_X1  g443(.A1(new_n636), .A2(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n643), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n637), .B1(new_n638), .B2(new_n412), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G134gat), .B(G162gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n645), .B(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n621), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT101), .Z(new_n654));
  NAND3_X1  g453(.A1(new_n623), .A2(new_n628), .A3(new_n631), .ZN(new_n655));
  INV_X1    g454(.A(new_n633), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n601), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n600), .B(new_n597), .C1(new_n632), .C2(new_n633), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT10), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n640), .A2(KEYINPUT10), .A3(new_n601), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n654), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n657), .A2(new_n658), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n654), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(G120gat), .B(G148gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(G176gat), .B(G204gat), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n667), .B(new_n668), .Z(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n663), .A2(new_n665), .A3(new_n669), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n495), .A2(new_n583), .A3(new_n652), .A4(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(new_n492), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT102), .B(G1gat), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1324gat));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n675), .A2(new_n286), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT16), .B(G8gat), .Z(new_n681));
  AOI21_X1  g480(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(G8gat), .B1(new_n675), .B2(new_n286), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n679), .A2(KEYINPUT103), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n685), .B1(new_n681), .B2(new_n686), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n682), .A2(new_n683), .B1(new_n680), .B2(new_n687), .ZN(G1325gat));
  NAND2_X1  g487(.A1(new_n439), .A2(new_n444), .ZN(new_n689));
  OAI21_X1  g488(.A(G15gat), .B1(new_n675), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n491), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n691), .A2(G15gat), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n690), .B1(new_n675), .B2(new_n692), .ZN(G1326gat));
  NOR2_X1   g492(.A1(new_n675), .A2(new_n484), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT43), .B(G22gat), .Z(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1327gat));
  AOI22_X1  g495(.A1(new_n485), .A2(new_n445), .B1(new_n488), .B2(new_n493), .ZN(new_n697));
  INV_X1    g496(.A(new_n651), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n582), .A2(new_n620), .A3(new_n673), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n492), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(new_n515), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT45), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n697), .B2(new_n698), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n495), .A2(KEYINPUT44), .A3(new_n651), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n700), .ZN(new_n710));
  OAI21_X1  g509(.A(G29gat), .B1(new_n710), .B2(new_n492), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n705), .A2(new_n711), .ZN(G1328gat));
  NOR3_X1   g511(.A1(new_n701), .A2(G36gat), .A3(new_n286), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT46), .ZN(new_n714));
  OAI21_X1  g513(.A(G36gat), .B1(new_n710), .B2(new_n286), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(G1329gat));
  OAI21_X1  g515(.A(new_n503), .B1(new_n701), .B2(new_n691), .ZN(new_n717));
  INV_X1    g516(.A(new_n689), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G43gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n717), .B1(new_n710), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g520(.A(G50gat), .B1(new_n710), .B2(new_n484), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT48), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n702), .A2(new_n506), .A3(new_n405), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n722), .B(new_n725), .C1(new_n723), .C2(KEYINPUT48), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1331gat));
  NAND3_X1  g528(.A1(new_n652), .A2(new_n582), .A3(new_n673), .ZN(new_n730));
  OR3_X1    g529(.A1(new_n697), .A2(KEYINPUT105), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT105), .B1(new_n697), .B2(new_n730), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n703), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g535(.A1(new_n733), .A2(new_n286), .ZN(new_n737));
  NOR2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  AND2_X1   g537(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(new_n737), .B2(new_n738), .ZN(G1333gat));
  OAI21_X1  g540(.A(G71gat), .B1(new_n733), .B2(new_n689), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n491), .A2(new_n584), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n733), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1334gat));
  NOR2_X1   g545(.A1(new_n733), .A2(new_n484), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(new_n585), .ZN(G1335gat));
  NOR2_X1   g547(.A1(new_n583), .A2(new_n620), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n495), .A2(new_n651), .A3(new_n749), .ZN(new_n750));
  OR2_X1    g549(.A1(new_n750), .A2(KEYINPUT51), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(KEYINPUT51), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n754), .A2(new_n629), .A3(new_n703), .A4(new_n673), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n583), .A2(new_n620), .A3(new_n674), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n709), .A2(new_n703), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n629), .B2(new_n757), .ZN(G1336gat));
  NOR3_X1   g557(.A1(new_n286), .A2(G92gat), .A3(new_n674), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n754), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761));
  INV_X1    g560(.A(new_n286), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n709), .A2(new_n762), .A3(new_n756), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G92gat), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n760), .A2(new_n761), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(KEYINPUT106), .A2(KEYINPUT51), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n766), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n495), .A2(new_n651), .A3(new_n749), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  AOI22_X1  g569(.A1(new_n763), .A2(G92gat), .B1(new_n770), .B2(new_n759), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n765), .B1(new_n771), .B2(new_n761), .ZN(G1337gat));
  NAND3_X1  g571(.A1(new_n709), .A2(new_n718), .A3(new_n756), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n624), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(new_n774), .B2(new_n773), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n754), .A2(new_n624), .A3(new_n491), .A4(new_n673), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(G1338gat));
  NAND4_X1  g577(.A1(new_n707), .A2(new_n708), .A3(new_n405), .A4(new_n756), .ZN(new_n779));
  XOR2_X1   g578(.A(KEYINPUT108), .B(G106gat), .Z(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n405), .A2(new_n625), .A3(new_n673), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n782), .B1(new_n767), .B2(new_n769), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI211_X1 g584(.A(KEYINPUT109), .B(new_n782), .C1(new_n767), .C2(new_n769), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT53), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT110), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n789), .B(KEYINPUT53), .C1(new_n785), .C2(new_n786), .ZN(new_n790));
  XNOR2_X1  g589(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n781), .B(new_n791), .C1(new_n753), .C2(new_n782), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n788), .A2(new_n790), .A3(new_n792), .ZN(G1339gat));
  NAND3_X1  g592(.A1(new_n698), .A2(new_n620), .A3(new_n674), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(new_n583), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n660), .A2(new_n661), .A3(new_n654), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n797), .A2(new_n662), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n660), .A2(new_n661), .ZN(new_n800));
  INV_X1    g599(.A(new_n654), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n800), .A2(new_n798), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n670), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n796), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n660), .A2(new_n661), .A3(new_n654), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n663), .A2(KEYINPUT54), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n669), .B1(new_n662), .B2(new_n798), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n806), .A2(KEYINPUT55), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n804), .A2(new_n672), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n501), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n573), .A2(new_n575), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n580), .A2(new_n564), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n576), .A2(new_n580), .A3(new_n564), .A4(new_n501), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n809), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n553), .A2(new_n555), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n570), .B1(new_n569), .B2(new_n571), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n500), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n814), .A2(new_n673), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n698), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n804), .A2(new_n672), .A3(new_n808), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n651), .A2(new_n814), .A3(new_n821), .A4(new_n818), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n620), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n820), .A2(KEYINPUT112), .A3(new_n822), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n795), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n405), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n691), .A2(new_n492), .A3(new_n762), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n317), .B1(new_n830), .B2(new_n583), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n827), .A2(new_n492), .A3(new_n487), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n832), .A2(new_n286), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n582), .A2(new_n324), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n831), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n835), .B(new_n836), .ZN(G1340gat));
  AOI21_X1  g636(.A(G120gat), .B1(new_n833), .B2(new_n673), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n674), .A2(new_n318), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n830), .B2(new_n839), .ZN(G1341gat));
  INV_X1    g639(.A(new_n830), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n326), .B1(new_n841), .B2(new_n621), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n621), .A2(new_n326), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n833), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(G1342gat));
  OAI21_X1  g644(.A(G134gat), .B1(new_n841), .B2(new_n698), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n286), .A2(new_n651), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT114), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(G134gat), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n832), .A2(new_n849), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n846), .A2(new_n851), .A3(new_n852), .ZN(G1343gat));
  NOR2_X1   g652(.A1(new_n492), .A2(new_n762), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n689), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  OAI211_X1 g656(.A(KEYINPUT115), .B(new_n857), .C1(new_n827), .C2(new_n484), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n405), .A2(KEYINPUT57), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n821), .B1(new_n577), .B2(new_n581), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n814), .A2(new_n673), .A3(new_n818), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(KEYINPUT116), .A3(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n864), .B1(new_n815), .B2(new_n819), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n865), .A3(new_n698), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n620), .B1(new_n866), .B2(new_n822), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n860), .B1(new_n867), .B2(new_n795), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n858), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n651), .B1(new_n861), .B2(new_n862), .ZN(new_n870));
  INV_X1    g669(.A(new_n822), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n824), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n621), .A3(new_n826), .ZN(new_n873));
  INV_X1    g672(.A(new_n795), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n405), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT115), .B1(new_n876), .B2(new_n857), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n856), .B1(new_n869), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n300), .B1(new_n878), .B2(new_n582), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n689), .A2(new_n405), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT117), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n703), .A3(new_n875), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(new_n762), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n583), .A2(new_n297), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(KEYINPUT118), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n879), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT58), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT58), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n879), .A2(new_n889), .A3(new_n886), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1344gat));
  NAND3_X1  g690(.A1(new_n883), .A2(new_n301), .A3(new_n673), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n301), .A2(KEYINPUT59), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n868), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT57), .B1(new_n875), .B2(new_n405), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(KEYINPUT115), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT115), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n827), .A2(new_n484), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(KEYINPUT57), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n855), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n894), .B1(new_n901), .B2(new_n673), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n405), .B1(new_n867), .B2(new_n795), .ZN(new_n903));
  AOI22_X1  g702(.A1(new_n903), .A2(new_n857), .B1(new_n875), .B2(new_n860), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n856), .A2(new_n673), .ZN(new_n905));
  OAI21_X1  g704(.A(G148gat), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n906), .A2(KEYINPUT59), .ZN(new_n907));
  OAI211_X1 g706(.A(KEYINPUT119), .B(new_n892), .C1(new_n902), .C2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n673), .B(new_n856), .C1(new_n869), .C2(new_n877), .ZN(new_n910));
  AOI22_X1  g709(.A1(new_n910), .A2(new_n893), .B1(KEYINPUT59), .B2(new_n906), .ZN(new_n911));
  INV_X1    g710(.A(new_n892), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n908), .A2(new_n913), .ZN(G1345gat));
  OAI21_X1  g713(.A(G155gat), .B1(new_n878), .B2(new_n621), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n883), .A2(new_n292), .A3(new_n620), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1346gat));
  OR2_X1    g716(.A1(new_n309), .A2(new_n310), .ZN(new_n918));
  OR3_X1    g717(.A1(new_n882), .A2(new_n918), .A3(new_n848), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n901), .A2(KEYINPUT120), .A3(new_n651), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n918), .ZN(new_n921));
  AOI21_X1  g720(.A(KEYINPUT120), .B1(new_n901), .B2(new_n651), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(G1347gat));
  NAND4_X1  g722(.A1(new_n828), .A2(new_n492), .A3(new_n762), .A4(new_n491), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n924), .A2(new_n203), .A3(new_n582), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n827), .A2(KEYINPUT121), .A3(new_n703), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n927), .B1(new_n875), .B2(new_n492), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n487), .A2(new_n286), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(new_n583), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n925), .B1(new_n934), .B2(new_n203), .ZN(G1348gat));
  OAI21_X1  g734(.A(G176gat), .B1(new_n924), .B2(new_n674), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n673), .A2(new_n204), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n932), .B2(new_n937), .ZN(G1349gat));
  OAI21_X1  g737(.A(G183gat), .B1(new_n924), .B2(new_n621), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n620), .A2(new_n212), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n932), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g740(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n941), .B(new_n943), .ZN(G1350gat));
  NAND3_X1  g743(.A1(new_n933), .A2(new_n213), .A3(new_n651), .ZN(new_n945));
  OAI21_X1  g744(.A(G190gat), .B1(new_n924), .B2(new_n698), .ZN(new_n946));
  XOR2_X1   g745(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n947));
  AND2_X1   g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G1351gat));
  NOR2_X1   g749(.A1(new_n880), .A2(new_n286), .ZN(new_n951));
  XOR2_X1   g750(.A(new_n951), .B(KEYINPUT124), .Z(new_n952));
  NAND2_X1  g751(.A1(new_n930), .A2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(G197gat), .B1(new_n954), .B2(new_n583), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n689), .A2(new_n492), .A3(new_n762), .ZN(new_n956));
  XOR2_X1   g755(.A(new_n956), .B(KEYINPUT125), .Z(new_n957));
  NOR2_X1   g756(.A1(new_n904), .A2(new_n957), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n583), .A2(G197gat), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  NOR2_X1   g759(.A1(new_n674), .A2(G204gat), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  OR3_X1    g761(.A1(new_n953), .A2(KEYINPUT62), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n958), .A2(new_n673), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G204gat), .ZN(new_n965));
  OAI21_X1  g764(.A(KEYINPUT62), .B1(new_n953), .B2(new_n962), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(G1353gat));
  INV_X1    g766(.A(G211gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n954), .A2(new_n968), .A3(new_n620), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n958), .B2(new_n620), .ZN(new_n970));
  OR2_X1    g769(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n973), .B1(new_n970), .B2(new_n971), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n969), .B1(new_n972), .B2(new_n974), .ZN(G1354gat));
  AOI21_X1  g774(.A(G218gat), .B1(new_n954), .B2(new_n651), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n651), .A2(G218gat), .ZN(new_n977));
  XOR2_X1   g776(.A(new_n977), .B(KEYINPUT127), .Z(new_n978));
  AOI21_X1  g777(.A(new_n976), .B1(new_n958), .B2(new_n978), .ZN(G1355gat));
endmodule


