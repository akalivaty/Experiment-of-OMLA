//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1199;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT67), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  OR2_X1    g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT68), .Z(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n462), .A2(G2105), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n463), .A2(new_n464), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(G160));
  INV_X1    g049(.A(new_n470), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(new_n469), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n476), .A2(G124), .B1(G136), .B2(new_n465), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT69), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n477), .A2(new_n481), .ZN(G162));
  NAND2_X1  g057(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n470), .A2(new_n469), .ZN(new_n484));
  INV_X1    g059(.A(G138), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(G126), .A2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n469), .A2(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(new_n483), .ZN(new_n489));
  OR2_X1    g064(.A1(new_n469), .A2(G114), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n489), .A2(new_n470), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n486), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  AND2_X1   g070(.A1(KEYINPUT6), .A2(G651), .ZN(new_n496));
  NOR2_X1   g071(.A1(KEYINPUT6), .A2(G651), .ZN(new_n497));
  OR2_X1    g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G543), .ZN(new_n499));
  INV_X1    g074(.A(G50), .ZN(new_n500));
  INV_X1    g075(.A(G88), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  OAI22_X1  g078(.A1(new_n502), .A2(new_n503), .B1(new_n496), .B2(new_n497), .ZN(new_n504));
  OAI22_X1  g079(.A1(new_n499), .A2(new_n500), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n505), .A2(new_n513), .ZN(G166));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT7), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT7), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n517), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G89), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n504), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT72), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n524), .B(new_n519), .C1(new_n504), .C2(new_n520), .ZN(new_n525));
  OAI21_X1  g100(.A(KEYINPUT71), .B1(new_n503), .B2(new_n502), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n508), .A2(new_n527), .A3(new_n509), .ZN(new_n528));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n526), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n496), .A2(new_n497), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n507), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G51), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n525), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n523), .A2(new_n534), .ZN(G168));
  NAND3_X1  g110(.A1(new_n526), .A2(new_n528), .A3(G64), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n512), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(G52), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n499), .A2(new_n539), .B1(new_n540), .B2(new_n504), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  NAND3_X1  g117(.A1(new_n526), .A2(new_n528), .A3(G56), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n543), .A2(KEYINPUT73), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(KEYINPUT73), .B1(new_n543), .B2(new_n544), .ZN(new_n546));
  NOR3_X1   g121(.A1(new_n545), .A2(new_n546), .A3(new_n512), .ZN(new_n547));
  INV_X1    g122(.A(new_n504), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n548), .A2(G81), .B1(new_n532), .B2(G43), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g128(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n554));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  OAI211_X1 g132(.A(G53), .B(G543), .C1(new_n496), .C2(new_n497), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n498), .A2(KEYINPUT75), .A3(new_n510), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n504), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n560), .A2(new_n562), .A3(G91), .ZN(new_n563));
  AND2_X1   g138(.A1(new_n510), .A2(G65), .ZN(new_n564));
  AND2_X1   g139(.A1(G78), .A2(G543), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n559), .A2(new_n563), .A3(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  INV_X1    g143(.A(G168), .ZN(G286));
  INV_X1    g144(.A(G166), .ZN(G303));
  AND2_X1   g145(.A1(new_n526), .A2(new_n528), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n571), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n560), .A2(new_n562), .A3(G87), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n532), .A2(G49), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  NAND3_X1  g150(.A1(new_n560), .A2(new_n562), .A3(G86), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT77), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT76), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n503), .A2(new_n502), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(G48), .B2(new_n532), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n577), .A2(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(new_n548), .A2(G85), .B1(new_n532), .B2(G47), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n571), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n586), .B2(new_n512), .ZN(G290));
  INV_X1    g162(.A(G868), .ZN(new_n588));
  NOR2_X1   g163(.A1(G301), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n560), .A2(new_n562), .A3(G92), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT10), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n560), .A2(new_n562), .A3(new_n592), .A4(G92), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n581), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(new_n532), .B2(G54), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n591), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT78), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n589), .B1(new_n599), .B2(new_n588), .ZN(G284));
  AOI21_X1  g175(.A(new_n589), .B1(new_n599), .B2(new_n588), .ZN(G321));
  NAND2_X1  g176(.A1(G299), .A2(new_n588), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G168), .B2(new_n588), .ZN(G297));
  OAI21_X1  g178(.A(new_n602), .B1(G168), .B2(new_n588), .ZN(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n599), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND2_X1  g181(.A1(new_n599), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n470), .A2(new_n466), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  INV_X1    g188(.A(G2100), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n476), .A2(G123), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n465), .A2(G135), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n469), .A2(G111), .ZN(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n616), .B(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2096), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n613), .A2(new_n614), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n615), .A2(new_n621), .A3(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(G2427), .B(G2438), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2430), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n627), .A2(new_n628), .A3(KEYINPUT14), .ZN(new_n629));
  XOR2_X1   g204(.A(G1341), .B(G1348), .Z(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n629), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G14), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n633), .A2(new_n636), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n638), .A2(new_n639), .ZN(G401));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n643), .A2(KEYINPUT17), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  AOI21_X1  g220(.A(KEYINPUT18), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2096), .B(G2100), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT81), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n643), .B2(KEYINPUT18), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT80), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(G227));
  XOR2_X1   g228(.A(G1971), .B(G1976), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1956), .B(G2474), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1961), .B(G1966), .Z(new_n658));
  AND2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT20), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n657), .A2(new_n658), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n655), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n655), .B2(new_n662), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G1991), .B(G1996), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT82), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n667), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1981), .B(G1986), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G229));
  MUX2_X1   g247(.A(G6), .B(G305), .S(G16), .Z(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT32), .B(G1981), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(G16), .A2(G23), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT85), .ZN(new_n677));
  INV_X1    g252(.A(G288), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n677), .B1(new_n678), .B2(G16), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT33), .B(G1976), .Z(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G22), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(G166), .B2(new_n683), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1971), .ZN(new_n686));
  NOR4_X1   g261(.A1(new_n675), .A2(new_n681), .A3(new_n682), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT84), .B(KEYINPUT34), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n476), .A2(G119), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n465), .A2(G131), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n469), .A2(G107), .ZN(new_n693));
  OAI21_X1  g268(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n691), .B(new_n692), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  MUX2_X1   g270(.A(G25), .B(new_n695), .S(G29), .Z(new_n696));
  XOR2_X1   g271(.A(KEYINPUT35), .B(G1991), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n683), .A2(G24), .ZN(new_n699));
  INV_X1    g274(.A(G290), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n683), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT83), .B(G1986), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND4_X1  g278(.A1(new_n689), .A2(new_n690), .A3(new_n698), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT36), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G35), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G162), .B2(new_n706), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G2090), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT93), .Z(new_n711));
  INV_X1    g286(.A(G34), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n712), .A2(KEYINPUT24), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(KEYINPUT24), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n706), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G160), .B2(new_n706), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT90), .Z(new_n717));
  INV_X1    g292(.A(G2084), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n683), .A2(G5), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G171), .B2(new_n683), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n719), .B1(G1961), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n683), .A2(G21), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G168), .B2(new_n683), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT91), .B(G1966), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NOR3_X1   g301(.A1(new_n711), .A2(new_n722), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n706), .A2(G33), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT25), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n731), .A2(new_n469), .ZN(new_n732));
  AOI211_X1 g307(.A(new_n730), .B(new_n732), .C1(G139), .C2(new_n465), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n728), .B1(new_n733), .B2(new_n706), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(G2072), .Z(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT26), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n476), .B2(G129), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n465), .A2(G141), .B1(G105), .B2(new_n466), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(new_n706), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n706), .B2(G32), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT27), .B(G1996), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OAI221_X1 g321(.A(new_n735), .B1(new_n709), .B2(G2090), .C1(new_n744), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n721), .A2(G1961), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n717), .B2(new_n718), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT31), .B(G11), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT92), .B(G28), .Z(new_n751));
  AOI21_X1  g326(.A(G29), .B1(new_n751), .B2(KEYINPUT30), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(KEYINPUT30), .B2(new_n751), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n750), .B(new_n753), .C1(new_n620), .C2(new_n706), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n744), .B2(new_n746), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n476), .A2(G128), .B1(G140), .B2(new_n465), .ZN(new_n756));
  INV_X1    g331(.A(G104), .ZN(new_n757));
  AND3_X1   g332(.A1(new_n757), .A2(new_n469), .A3(KEYINPUT88), .ZN(new_n758));
  AOI21_X1  g333(.A(KEYINPUT88), .B1(new_n757), .B2(new_n469), .ZN(new_n759));
  OAI221_X1 g334(.A(G2104), .B1(G116), .B2(new_n469), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G29), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n706), .A2(G26), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G2067), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n706), .A2(G27), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G164), .B2(new_n706), .ZN(new_n770));
  INV_X1    g345(.A(G2078), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n755), .A2(new_n768), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT94), .B(KEYINPUT23), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n683), .A2(G20), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G299), .B2(G16), .ZN(new_n777));
  INV_X1    g352(.A(G1956), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NOR4_X1   g354(.A1(new_n747), .A2(new_n749), .A3(new_n773), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n683), .A2(G19), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n551), .B2(new_n683), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT86), .B(G1341), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT87), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n782), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n683), .A2(G4), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n599), .B2(new_n683), .ZN(new_n787));
  INV_X1    g362(.A(G1348), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n727), .A2(new_n780), .A3(new_n785), .A4(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT95), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n705), .A2(new_n791), .ZN(G150));
  INV_X1    g367(.A(G150), .ZN(G311));
  AOI22_X1  g368(.A1(new_n548), .A2(G93), .B1(new_n532), .B2(G55), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n526), .A2(new_n528), .A3(G67), .ZN(new_n795));
  NAND2_X1  g370(.A1(G80), .A2(G543), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n512), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT98), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI211_X1 g374(.A(KEYINPUT98), .B(new_n512), .C1(new_n795), .C2(new_n796), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(G860), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT37), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n599), .A2(G559), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT97), .ZN(new_n806));
  OAI22_X1  g381(.A1(new_n547), .A2(new_n550), .B1(new_n799), .B2(new_n800), .ZN(new_n807));
  INV_X1    g382(.A(G55), .ZN(new_n808));
  INV_X1    g383(.A(G93), .ZN(new_n809));
  OAI22_X1  g384(.A1(new_n499), .A2(new_n808), .B1(new_n809), .B2(new_n504), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n795), .A2(new_n796), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G651), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n810), .B1(new_n812), .B2(KEYINPUT98), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n543), .A2(new_n544), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT73), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n543), .A2(KEYINPUT73), .A3(new_n544), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n816), .A2(G651), .A3(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n800), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n813), .A2(new_n818), .A3(new_n549), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n807), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n806), .B(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n824), .A2(KEYINPUT39), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n802), .B1(new_n824), .B2(KEYINPUT39), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n804), .B1(new_n825), .B2(new_n826), .ZN(G145));
  XNOR2_X1  g402(.A(new_n733), .B(new_n740), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n695), .B(new_n612), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n761), .B(G164), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n476), .A2(G130), .B1(G142), .B2(new_n465), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT99), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n833), .A2(new_n469), .A3(G118), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n469), .B2(G118), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n835), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n832), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n831), .B(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n830), .B(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n620), .B(G160), .Z(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(G162), .Z(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(G37), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n839), .A2(new_n841), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT40), .Z(G395));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n807), .A3(new_n820), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n599), .A2(new_n821), .A3(new_n605), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(G299), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n598), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n598), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(G299), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n598), .A2(new_n851), .A3(KEYINPUT100), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT41), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n854), .A2(KEYINPUT41), .A3(new_n856), .A4(new_n857), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n850), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT42), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n848), .A2(new_n849), .A3(new_n858), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n864), .B1(new_n863), .B2(new_n865), .ZN(new_n867));
  XNOR2_X1  g442(.A(G305), .B(new_n700), .ZN(new_n868));
  XNOR2_X1  g443(.A(G303), .B(G288), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  OR3_X1    g446(.A1(new_n866), .A2(new_n867), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n871), .B1(new_n866), .B2(new_n867), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(G868), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n875));
  INV_X1    g450(.A(new_n801), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n875), .B1(new_n876), .B2(new_n588), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n872), .A2(new_n875), .A3(G868), .A4(new_n873), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(G295));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n880), .B(new_n883), .ZN(G331));
  INV_X1    g459(.A(KEYINPUT109), .ZN(new_n885));
  OAI22_X1  g460(.A1(new_n523), .A2(new_n534), .B1(new_n538), .B2(new_n541), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n533), .A2(new_n530), .ZN(new_n887));
  NAND4_X1  g462(.A1(G171), .A2(new_n887), .A3(new_n522), .A4(new_n525), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n807), .A2(new_n820), .A3(new_n886), .A4(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT104), .ZN(new_n890));
  AOI221_X4 g465(.A(new_n890), .B1(new_n888), .B2(new_n886), .C1(new_n807), .C2(new_n820), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n886), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT104), .B1(new_n821), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n889), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n862), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n858), .A2(new_n889), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n821), .A2(new_n892), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT105), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n821), .A2(new_n900), .A3(new_n892), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n843), .B1(new_n903), .B2(new_n870), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n899), .A2(new_n889), .A3(new_n901), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n860), .A2(new_n907), .A3(new_n861), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n861), .A2(new_n907), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n891), .A2(new_n893), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT107), .B1(new_n911), .B2(new_n896), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n897), .B(new_n913), .C1(new_n893), .C2(new_n891), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n910), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n915), .A2(KEYINPUT108), .A3(new_n870), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT108), .B1(new_n915), .B2(new_n870), .ZN(new_n917));
  OAI211_X1 g492(.A(KEYINPUT43), .B(new_n905), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n871), .B1(new_n895), .B2(new_n902), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n919), .B1(new_n904), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT44), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n919), .B(new_n905), .C1(new_n916), .C2(new_n917), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT43), .B1(new_n904), .B2(new_n920), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n885), .B1(new_n923), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n927), .B1(new_n918), .B2(new_n921), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT44), .B1(new_n924), .B2(new_n925), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT109), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n929), .A2(new_n932), .ZN(G397));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n934));
  AOI21_X1  g509(.A(G1384), .B1(new_n486), .B2(new_n493), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n934), .B1(new_n935), .B2(KEYINPUT110), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(KEYINPUT110), .B2(new_n935), .ZN(new_n937));
  INV_X1    g512(.A(G40), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n468), .A2(new_n473), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G1996), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n940), .A2(new_n941), .A3(new_n741), .ZN(new_n942));
  OR2_X1    g517(.A1(new_n942), .A2(KEYINPUT112), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(KEYINPUT112), .ZN(new_n944));
  INV_X1    g519(.A(new_n940), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n761), .B(new_n767), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(G1996), .B2(new_n740), .ZN(new_n947));
  AOI22_X1  g522(.A1(new_n943), .A2(new_n944), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n697), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n695), .A2(new_n949), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n695), .A2(new_n949), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n945), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G1986), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n700), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT111), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(new_n954), .B2(new_n700), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n953), .B1(new_n945), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G8), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n935), .A2(KEYINPUT113), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT113), .ZN(new_n962));
  AOI211_X1 g537(.A(new_n962), .B(G1384), .C1(new_n486), .C2(new_n493), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n960), .B1(new_n964), .B2(new_n939), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1981), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n577), .A2(new_n967), .A3(new_n583), .ZN(new_n968));
  INV_X1    g543(.A(G86), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n583), .B1(new_n969), .B2(new_n504), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(G1981), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT49), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n968), .A2(KEYINPUT49), .A3(new_n971), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(new_n965), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G1976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(new_n977), .A3(new_n678), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n966), .B1(new_n978), .B2(new_n968), .ZN(new_n979));
  INV_X1    g554(.A(new_n935), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n962), .ZN(new_n981));
  INV_X1    g556(.A(new_n963), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n981), .A2(new_n982), .A3(new_n939), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n678), .A2(G1976), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(G8), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT52), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT52), .B1(G288), .B2(new_n977), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n965), .A2(new_n984), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n976), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT115), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n986), .A2(new_n988), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n991), .A2(new_n992), .A3(new_n976), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n995));
  OAI211_X1 g570(.A(G8), .B(new_n995), .C1(new_n505), .C2(new_n513), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(G303), .A2(G8), .ZN(new_n998));
  NAND2_X1  g573(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G2090), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n939), .B1(new_n935), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n981), .A2(new_n982), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n1001), .B(new_n1004), .C1(new_n1005), .C2(KEYINPUT50), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n471), .A2(new_n472), .ZN(new_n1007));
  OAI211_X1 g582(.A(G40), .B(new_n467), .C1(new_n1007), .C2(new_n469), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(KEYINPUT45), .B2(new_n935), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n935), .A2(KEYINPUT45), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1971), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI211_X1 g589(.A(new_n960), .B(new_n1000), .C1(new_n1006), .C2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n979), .B1(new_n994), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n960), .B1(new_n1006), .B2(new_n1014), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1000), .ZN(new_n1018));
  OR2_X1    g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(G168), .A2(G8), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n934), .B1(new_n961), .B2(new_n963), .ZN(new_n1022));
  AOI21_X1  g597(.A(G1966), .B1(new_n1022), .B2(new_n1009), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n961), .A2(new_n963), .A3(KEYINPUT50), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(new_n1003), .ZN(new_n1025));
  AOI22_X1  g600(.A1(new_n1021), .A2(new_n1023), .B1(new_n1025), .B2(new_n718), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1022), .A2(new_n1009), .ZN(new_n1027));
  INV_X1    g602(.A(G1966), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT116), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1020), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT63), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1019), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1034), .B1(new_n990), .B2(new_n993), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1008), .B1(new_n1002), .B2(new_n935), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(new_n964), .B2(new_n1002), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1014), .B1(new_n1037), .B2(G2090), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1018), .B1(new_n1038), .B2(G8), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n989), .A2(new_n1039), .A3(new_n1015), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT63), .B1(new_n1040), .B2(new_n1031), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1016), .B1(new_n1035), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G1384), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n494), .A2(KEYINPUT45), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n939), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1045), .A2(G2078), .A3(new_n1010), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT124), .B1(new_n1046), .B2(KEYINPUT53), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT124), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1048), .B(new_n1049), .C1(new_n1012), .C2(G2078), .ZN(new_n1050));
  INV_X1    g625(.A(G1961), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1051), .B1(new_n1024), .B2(new_n1003), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1022), .A2(KEYINPUT53), .A3(new_n771), .A4(new_n1009), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1047), .A2(new_n1050), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G171), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT125), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT125), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1054), .A2(new_n1057), .A3(G171), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1047), .A2(new_n1052), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1009), .A2(KEYINPUT53), .A3(new_n771), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1060), .A2(new_n937), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1059), .A2(G301), .A3(new_n1050), .A4(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1056), .A2(new_n1058), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1025), .A2(new_n718), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1023), .A2(new_n1021), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1030), .A2(G168), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G8), .ZN(new_n1069));
  AOI21_X1  g644(.A(G168), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT51), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1068), .A2(new_n1072), .A3(G8), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1038), .A2(G8), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n1000), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1076), .A2(new_n976), .A3(new_n991), .A4(new_n1077), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n1054), .A2(G171), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1061), .A2(new_n1047), .A3(new_n1050), .A4(new_n1052), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1064), .B1(new_n1080), .B2(G171), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1078), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1065), .A2(new_n1074), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1037), .A2(new_n778), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n1085));
  XNOR2_X1  g660(.A(G299), .B(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n559), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1088), .A2(KEYINPUT57), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(G299), .B(KEYINPUT118), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1089), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT56), .B(G2072), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1009), .A2(new_n1011), .A3(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1084), .A2(new_n1090), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT122), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1100), .A2(new_n1101), .A3(new_n1084), .A4(new_n1095), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1097), .A2(new_n1102), .A3(KEYINPUT61), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1084), .A2(new_n1095), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1090), .A2(new_n1093), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1105), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1104), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT119), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n1106), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1114), .A2(KEYINPUT120), .A3(new_n1104), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1103), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT61), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1104), .A2(new_n1112), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1096), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT121), .B1(new_n1012), .B2(G1996), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1009), .A2(new_n1011), .A3(new_n1122), .A4(new_n941), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT58), .B(G1341), .Z(new_n1124));
  NAND2_X1  g699(.A1(new_n983), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1121), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n551), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT59), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n1129), .A3(new_n551), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  XOR2_X1   g706(.A(new_n598), .B(KEYINPUT123), .Z(new_n1132));
  OAI21_X1  g707(.A(new_n788), .B1(new_n1024), .B2(new_n1003), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n964), .A2(new_n767), .A3(new_n939), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1132), .A2(new_n1133), .A3(KEYINPUT60), .A4(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n598), .A2(KEYINPUT123), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1135), .B(new_n1138), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1120), .A2(new_n1131), .A3(new_n1141), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1111), .A2(new_n1115), .B1(new_n855), .B2(new_n1136), .ZN(new_n1143));
  OAI22_X1  g718(.A1(new_n1116), .A2(new_n1142), .B1(new_n1143), .B2(new_n1119), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1042), .B1(new_n1083), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1146), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n1040), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1150), .B1(KEYINPUT62), .B2(new_n1074), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n959), .B1(new_n1145), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n948), .A2(new_n950), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(G2067), .B2(new_n761), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n945), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n945), .A2(new_n941), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT46), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n946), .A2(new_n741), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1157), .B1(new_n940), .B2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT47), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n956), .A2(new_n940), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT48), .Z(new_n1162));
  NAND3_X1  g737(.A1(new_n1162), .A2(new_n952), .A3(new_n948), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1155), .A2(new_n1160), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(KEYINPUT126), .B1(new_n1152), .B2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1039), .A2(new_n1015), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1166), .A2(new_n976), .A3(new_n991), .A4(new_n1031), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1019), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1168));
  AOI22_X1  g743(.A1(new_n1032), .A2(new_n1167), .B1(new_n1168), .B2(new_n994), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n994), .A2(new_n1015), .ZN(new_n1170));
  INV_X1    g745(.A(new_n979), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1120), .A2(new_n1131), .A3(new_n1141), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1117), .B1(new_n1119), .B2(new_n1101), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1176));
  AOI21_X1  g751(.A(KEYINPUT120), .B1(new_n1114), .B2(new_n1104), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1097), .B(new_n1175), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1136), .A2(new_n855), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1179), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1180));
  AOI22_X1  g755(.A1(new_n1174), .A2(new_n1178), .B1(new_n1180), .B2(new_n1096), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1065), .A2(new_n1074), .A3(new_n1082), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1173), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1074), .A2(KEYINPUT62), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n1184), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n958), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1164), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1165), .A2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g765(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1192));
  NOR3_X1   g766(.A1(new_n846), .A2(G229), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n1194));
  NAND3_X1  g768(.A1(new_n1193), .A2(new_n1194), .A3(new_n926), .ZN(new_n1195));
  INV_X1    g769(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g770(.A(new_n1194), .B1(new_n1193), .B2(new_n926), .ZN(new_n1197));
  NOR2_X1   g771(.A1(new_n1196), .A2(new_n1197), .ZN(G308));
  INV_X1    g772(.A(new_n1197), .ZN(new_n1199));
  NAND2_X1  g773(.A1(new_n1199), .A2(new_n1195), .ZN(G225));
endmodule


