

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U555 ( .A1(n605), .A2(n702), .ZN(n673) );
  NOR2_X1 U556 ( .A1(n975), .A2(n621), .ZN(n632) );
  INV_X1 U557 ( .A(KEYINPUT103), .ZN(n639) );
  XNOR2_X1 U558 ( .A(n640), .B(n639), .ZN(n653) );
  AND2_X1 U559 ( .A1(G40), .A2(G160), .ZN(n605) );
  NOR2_X1 U560 ( .A1(G651), .A2(n584), .ZN(n812) );
  XOR2_X1 U561 ( .A(KEYINPUT4), .B(KEYINPUT74), .Z(n524) );
  NOR2_X1 U562 ( .A1(G651), .A2(G543), .ZN(n807) );
  NAND2_X1 U563 ( .A1(G89), .A2(n807), .ZN(n523) );
  XNOR2_X1 U564 ( .A(n524), .B(n523), .ZN(n528) );
  XNOR2_X1 U565 ( .A(G543), .B(KEYINPUT0), .ZN(n525) );
  XNOR2_X1 U566 ( .A(n525), .B(KEYINPUT67), .ZN(n584) );
  INV_X1 U567 ( .A(G651), .ZN(n531) );
  NOR2_X1 U568 ( .A1(n584), .A2(n531), .ZN(n808) );
  NAND2_X1 U569 ( .A1(n808), .A2(G76), .ZN(n526) );
  XNOR2_X1 U570 ( .A(KEYINPUT75), .B(n526), .ZN(n527) );
  NOR2_X1 U571 ( .A1(n528), .A2(n527), .ZN(n530) );
  XNOR2_X1 U572 ( .A(KEYINPUT5), .B(KEYINPUT76), .ZN(n529) );
  XNOR2_X1 U573 ( .A(n530), .B(n529), .ZN(n537) );
  NOR2_X1 U574 ( .A1(G543), .A2(n531), .ZN(n532) );
  XOR2_X1 U575 ( .A(KEYINPUT1), .B(n532), .Z(n815) );
  NAND2_X1 U576 ( .A1(G63), .A2(n815), .ZN(n534) );
  NAND2_X1 U577 ( .A1(G51), .A2(n812), .ZN(n533) );
  NAND2_X1 U578 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U579 ( .A(KEYINPUT6), .B(n535), .ZN(n536) );
  NOR2_X1 U580 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U581 ( .A(KEYINPUT7), .B(n538), .Z(G168) );
  XOR2_X1 U582 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n539) );
  XOR2_X1 U584 ( .A(KEYINPUT17), .B(n539), .Z(n540) );
  XNOR2_X2 U585 ( .A(n540), .B(KEYINPUT66), .ZN(n893) );
  NAND2_X1 U586 ( .A1(G137), .A2(n893), .ZN(n549) );
  XOR2_X1 U587 ( .A(KEYINPUT23), .B(KEYINPUT65), .Z(n542) );
  INV_X1 U588 ( .A(G2105), .ZN(n543) );
  AND2_X1 U589 ( .A1(n543), .A2(G2104), .ZN(n892) );
  NAND2_X1 U590 ( .A1(G101), .A2(n892), .ZN(n541) );
  XNOR2_X1 U591 ( .A(n542), .B(n541), .ZN(n547) );
  AND2_X1 U592 ( .A1(G2104), .A2(G2105), .ZN(n896) );
  NAND2_X1 U593 ( .A1(G113), .A2(n896), .ZN(n545) );
  NOR2_X1 U594 ( .A1(G2104), .A2(n543), .ZN(n897) );
  NAND2_X1 U595 ( .A1(G125), .A2(n897), .ZN(n544) );
  NAND2_X1 U596 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U597 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U598 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X2 U599 ( .A(KEYINPUT64), .B(n550), .Z(G160) );
  XOR2_X1 U600 ( .A(G2435), .B(G2454), .Z(n552) );
  XNOR2_X1 U601 ( .A(G2430), .B(G2438), .ZN(n551) );
  XNOR2_X1 U602 ( .A(n552), .B(n551), .ZN(n559) );
  XOR2_X1 U603 ( .A(G2446), .B(KEYINPUT113), .Z(n554) );
  XNOR2_X1 U604 ( .A(G2451), .B(G2443), .ZN(n553) );
  XNOR2_X1 U605 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U606 ( .A(n555), .B(G2427), .Z(n557) );
  XNOR2_X1 U607 ( .A(G1348), .B(G1341), .ZN(n556) );
  XNOR2_X1 U608 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U609 ( .A(n559), .B(n558), .ZN(n560) );
  AND2_X1 U610 ( .A1(n560), .A2(G14), .ZN(G401) );
  NAND2_X1 U611 ( .A1(n812), .A2(G52), .ZN(n562) );
  NAND2_X1 U612 ( .A1(n815), .A2(G64), .ZN(n561) );
  NAND2_X1 U613 ( .A1(n562), .A2(n561), .ZN(n567) );
  NAND2_X1 U614 ( .A1(G90), .A2(n807), .ZN(n564) );
  NAND2_X1 U615 ( .A1(G77), .A2(n808), .ZN(n563) );
  NAND2_X1 U616 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U617 ( .A(KEYINPUT9), .B(n565), .Z(n566) );
  NOR2_X1 U618 ( .A1(n567), .A2(n566), .ZN(G171) );
  AND2_X1 U619 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U620 ( .A(G57), .ZN(G237) );
  INV_X1 U621 ( .A(G69), .ZN(G235) );
  INV_X1 U622 ( .A(G108), .ZN(G238) );
  INV_X1 U623 ( .A(G120), .ZN(G236) );
  INV_X1 U624 ( .A(G132), .ZN(G219) );
  INV_X1 U625 ( .A(G82), .ZN(G220) );
  NAND2_X1 U626 ( .A1(G102), .A2(n892), .ZN(n569) );
  NAND2_X1 U627 ( .A1(G138), .A2(n893), .ZN(n568) );
  NAND2_X1 U628 ( .A1(n569), .A2(n568), .ZN(n574) );
  NAND2_X1 U629 ( .A1(G114), .A2(n896), .ZN(n571) );
  NAND2_X1 U630 ( .A1(G126), .A2(n897), .ZN(n570) );
  NAND2_X1 U631 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U632 ( .A(KEYINPUT93), .B(n572), .Z(n573) );
  NOR2_X1 U633 ( .A1(n574), .A2(n573), .ZN(G164) );
  NAND2_X1 U634 ( .A1(G88), .A2(n807), .ZN(n575) );
  XNOR2_X1 U635 ( .A(n575), .B(KEYINPUT88), .ZN(n582) );
  NAND2_X1 U636 ( .A1(G62), .A2(n815), .ZN(n577) );
  NAND2_X1 U637 ( .A1(G50), .A2(n812), .ZN(n576) );
  NAND2_X1 U638 ( .A1(n577), .A2(n576), .ZN(n580) );
  NAND2_X1 U639 ( .A1(G75), .A2(n808), .ZN(n578) );
  XNOR2_X1 U640 ( .A(KEYINPUT89), .B(n578), .ZN(n579) );
  NOR2_X1 U641 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U642 ( .A1(n582), .A2(n581), .ZN(G303) );
  INV_X1 U643 ( .A(G303), .ZN(G166) );
  NAND2_X1 U644 ( .A1(G74), .A2(G651), .ZN(n583) );
  XNOR2_X1 U645 ( .A(n583), .B(KEYINPUT86), .ZN(n589) );
  NAND2_X1 U646 ( .A1(G49), .A2(n812), .ZN(n586) );
  NAND2_X1 U647 ( .A1(G87), .A2(n584), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U649 ( .A1(n815), .A2(n587), .ZN(n588) );
  NAND2_X1 U650 ( .A1(n589), .A2(n588), .ZN(G288) );
  NAND2_X1 U651 ( .A1(G73), .A2(n808), .ZN(n590) );
  XNOR2_X1 U652 ( .A(n590), .B(KEYINPUT2), .ZN(n597) );
  NAND2_X1 U653 ( .A1(G86), .A2(n807), .ZN(n592) );
  NAND2_X1 U654 ( .A1(G61), .A2(n815), .ZN(n591) );
  NAND2_X1 U655 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U656 ( .A1(G48), .A2(n812), .ZN(n593) );
  XNOR2_X1 U657 ( .A(KEYINPUT87), .B(n593), .ZN(n594) );
  NOR2_X1 U658 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U659 ( .A1(n597), .A2(n596), .ZN(G305) );
  NAND2_X1 U660 ( .A1(G85), .A2(n807), .ZN(n599) );
  NAND2_X1 U661 ( .A1(G60), .A2(n815), .ZN(n598) );
  NAND2_X1 U662 ( .A1(n599), .A2(n598), .ZN(n603) );
  NAND2_X1 U663 ( .A1(G72), .A2(n808), .ZN(n601) );
  NAND2_X1 U664 ( .A1(G47), .A2(n812), .ZN(n600) );
  NAND2_X1 U665 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U666 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U667 ( .A(KEYINPUT68), .B(n604), .Z(G290) );
  INV_X1 U668 ( .A(KEYINPUT40), .ZN(n775) );
  NOR2_X1 U669 ( .A1(G164), .A2(G1384), .ZN(n702) );
  XNOR2_X1 U670 ( .A(G2078), .B(KEYINPUT25), .ZN(n955) );
  NOR2_X1 U671 ( .A1(n673), .A2(n955), .ZN(n607) );
  INV_X1 U672 ( .A(n673), .ZN(n642) );
  INV_X1 U673 ( .A(G1961), .ZN(n1008) );
  NOR2_X1 U674 ( .A1(n642), .A2(n1008), .ZN(n606) );
  NOR2_X1 U675 ( .A1(n607), .A2(n606), .ZN(n666) );
  NAND2_X1 U676 ( .A1(G171), .A2(n666), .ZN(n662) );
  NAND2_X1 U677 ( .A1(G56), .A2(n815), .ZN(n608) );
  XOR2_X1 U678 ( .A(KEYINPUT14), .B(n608), .Z(n614) );
  NAND2_X1 U679 ( .A1(n807), .A2(G81), .ZN(n609) );
  XNOR2_X1 U680 ( .A(n609), .B(KEYINPUT12), .ZN(n611) );
  NAND2_X1 U681 ( .A1(G68), .A2(n808), .ZN(n610) );
  NAND2_X1 U682 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U683 ( .A(KEYINPUT13), .B(n612), .Z(n613) );
  NOR2_X1 U684 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U685 ( .A1(n812), .A2(G43), .ZN(n615) );
  NAND2_X1 U686 ( .A1(n616), .A2(n615), .ZN(n975) );
  INV_X1 U687 ( .A(n673), .ZN(n617) );
  NAND2_X1 U688 ( .A1(n617), .A2(G1996), .ZN(n618) );
  XNOR2_X1 U689 ( .A(n618), .B(KEYINPUT26), .ZN(n620) );
  NAND2_X1 U690 ( .A1(n673), .A2(G1341), .ZN(n619) );
  NAND2_X1 U691 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U692 ( .A1(G79), .A2(n808), .ZN(n623) );
  NAND2_X1 U693 ( .A1(G54), .A2(n812), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U695 ( .A(KEYINPUT72), .B(n624), .ZN(n627) );
  NAND2_X1 U696 ( .A1(G66), .A2(n815), .ZN(n625) );
  XNOR2_X1 U697 ( .A(KEYINPUT71), .B(n625), .ZN(n626) );
  NOR2_X1 U698 ( .A1(n627), .A2(n626), .ZN(n629) );
  NAND2_X1 U699 ( .A1(n807), .A2(G92), .ZN(n628) );
  NAND2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U701 ( .A(KEYINPUT15), .B(n630), .ZN(n985) );
  NOR2_X1 U702 ( .A1(n632), .A2(n985), .ZN(n631) );
  XOR2_X1 U703 ( .A(n631), .B(KEYINPUT102), .Z(n638) );
  NAND2_X1 U704 ( .A1(n632), .A2(n985), .ZN(n636) );
  NOR2_X1 U705 ( .A1(G2067), .A2(n673), .ZN(n634) );
  NOR2_X1 U706 ( .A1(n642), .A2(G1348), .ZN(n633) );
  NOR2_X1 U707 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U709 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U710 ( .A1(n642), .A2(G2072), .ZN(n641) );
  XNOR2_X1 U711 ( .A(n641), .B(KEYINPUT27), .ZN(n644) );
  INV_X1 U712 ( .A(G1956), .ZN(n999) );
  NOR2_X1 U713 ( .A1(n999), .A2(n642), .ZN(n643) );
  NOR2_X1 U714 ( .A1(n644), .A2(n643), .ZN(n654) );
  NAND2_X1 U715 ( .A1(n808), .A2(G78), .ZN(n647) );
  NAND2_X1 U716 ( .A1(G65), .A2(n815), .ZN(n645) );
  XOR2_X1 U717 ( .A(KEYINPUT69), .B(n645), .Z(n646) );
  NAND2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U719 ( .A1(G91), .A2(n807), .ZN(n649) );
  NAND2_X1 U720 ( .A1(G53), .A2(n812), .ZN(n648) );
  NAND2_X1 U721 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U722 ( .A1(n651), .A2(n650), .ZN(n980) );
  NAND2_X1 U723 ( .A1(n654), .A2(n980), .ZN(n652) );
  NAND2_X1 U724 ( .A1(n653), .A2(n652), .ZN(n658) );
  NOR2_X1 U725 ( .A1(n654), .A2(n980), .ZN(n656) );
  XNOR2_X1 U726 ( .A(KEYINPUT28), .B(KEYINPUT101), .ZN(n655) );
  XNOR2_X1 U727 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n660) );
  XOR2_X1 U729 ( .A(KEYINPUT104), .B(KEYINPUT29), .Z(n659) );
  XNOR2_X1 U730 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X1 U731 ( .A1(n662), .A2(n661), .ZN(n684) );
  NAND2_X1 U732 ( .A1(G8), .A2(n673), .ZN(n751) );
  NOR2_X1 U733 ( .A1(G1966), .A2(n751), .ZN(n686) );
  NOR2_X1 U734 ( .A1(G2084), .A2(n673), .ZN(n682) );
  NOR2_X1 U735 ( .A1(n686), .A2(n682), .ZN(n663) );
  NAND2_X1 U736 ( .A1(G8), .A2(n663), .ZN(n664) );
  XNOR2_X1 U737 ( .A(KEYINPUT30), .B(n664), .ZN(n665) );
  NOR2_X1 U738 ( .A1(G168), .A2(n665), .ZN(n668) );
  NOR2_X1 U739 ( .A1(G171), .A2(n666), .ZN(n667) );
  NOR2_X1 U740 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U741 ( .A(n669), .B(KEYINPUT105), .ZN(n670) );
  XNOR2_X1 U742 ( .A(n670), .B(KEYINPUT31), .ZN(n683) );
  NAND2_X1 U743 ( .A1(n684), .A2(n683), .ZN(n671) );
  NAND2_X1 U744 ( .A1(n671), .A2(G286), .ZN(n672) );
  XNOR2_X1 U745 ( .A(n672), .B(KEYINPUT106), .ZN(n679) );
  NOR2_X1 U746 ( .A1(G2090), .A2(n673), .ZN(n674) );
  XNOR2_X1 U747 ( .A(KEYINPUT107), .B(n674), .ZN(n677) );
  NOR2_X1 U748 ( .A1(G1971), .A2(n751), .ZN(n675) );
  NOR2_X1 U749 ( .A1(G166), .A2(n675), .ZN(n676) );
  NAND2_X1 U750 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U751 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U752 ( .A1(n680), .A2(G8), .ZN(n681) );
  XNOR2_X1 U753 ( .A(KEYINPUT32), .B(n681), .ZN(n742) );
  NAND2_X1 U754 ( .A1(G8), .A2(n682), .ZN(n688) );
  AND2_X1 U755 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U756 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U757 ( .A1(n688), .A2(n687), .ZN(n740) );
  NAND2_X1 U758 ( .A1(G1976), .A2(G288), .ZN(n978) );
  AND2_X1 U759 ( .A1(n740), .A2(n978), .ZN(n689) );
  NAND2_X1 U760 ( .A1(n742), .A2(n689), .ZN(n698) );
  INV_X1 U761 ( .A(n978), .ZN(n694) );
  NOR2_X1 U762 ( .A1(G1976), .A2(G288), .ZN(n977) );
  NOR2_X1 U763 ( .A1(G1971), .A2(G303), .ZN(n690) );
  XNOR2_X1 U764 ( .A(KEYINPUT108), .B(n690), .ZN(n691) );
  NOR2_X1 U765 ( .A1(n977), .A2(n691), .ZN(n692) );
  XOR2_X1 U766 ( .A(KEYINPUT109), .B(n692), .Z(n693) );
  OR2_X1 U767 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U768 ( .A1(n751), .A2(n695), .ZN(n696) );
  NOR2_X1 U769 ( .A1(n696), .A2(KEYINPUT33), .ZN(n697) );
  NAND2_X1 U770 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U771 ( .A(n699), .B(KEYINPUT110), .ZN(n739) );
  NAND2_X1 U772 ( .A1(n977), .A2(KEYINPUT33), .ZN(n700) );
  NOR2_X1 U773 ( .A1(n751), .A2(n700), .ZN(n737) );
  XOR2_X1 U774 ( .A(G1981), .B(G305), .Z(n972) );
  NAND2_X1 U775 ( .A1(G40), .A2(G160), .ZN(n701) );
  NOR2_X1 U776 ( .A1(n702), .A2(n701), .ZN(n767) );
  NAND2_X1 U777 ( .A1(G117), .A2(n896), .ZN(n704) );
  NAND2_X1 U778 ( .A1(G129), .A2(n897), .ZN(n703) );
  NAND2_X1 U779 ( .A1(n704), .A2(n703), .ZN(n707) );
  NAND2_X1 U780 ( .A1(n892), .A2(G105), .ZN(n705) );
  XOR2_X1 U781 ( .A(KEYINPUT38), .B(n705), .Z(n706) );
  NOR2_X1 U782 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U783 ( .A(n708), .B(KEYINPUT98), .ZN(n710) );
  NAND2_X1 U784 ( .A1(G141), .A2(n893), .ZN(n709) );
  NAND2_X1 U785 ( .A1(n710), .A2(n709), .ZN(n906) );
  NAND2_X1 U786 ( .A1(G1996), .A2(n906), .ZN(n720) );
  NAND2_X1 U787 ( .A1(G119), .A2(n897), .ZN(n711) );
  XNOR2_X1 U788 ( .A(n711), .B(KEYINPUT96), .ZN(n718) );
  NAND2_X1 U789 ( .A1(G95), .A2(n892), .ZN(n713) );
  NAND2_X1 U790 ( .A1(G131), .A2(n893), .ZN(n712) );
  NAND2_X1 U791 ( .A1(n713), .A2(n712), .ZN(n716) );
  NAND2_X1 U792 ( .A1(G107), .A2(n896), .ZN(n714) );
  XNOR2_X1 U793 ( .A(KEYINPUT97), .B(n714), .ZN(n715) );
  NOR2_X1 U794 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U795 ( .A1(n718), .A2(n717), .ZN(n879) );
  NAND2_X1 U796 ( .A1(G1991), .A2(n879), .ZN(n719) );
  NAND2_X1 U797 ( .A1(n720), .A2(n719), .ZN(n935) );
  NAND2_X1 U798 ( .A1(n767), .A2(n935), .ZN(n756) );
  NAND2_X1 U799 ( .A1(G104), .A2(n892), .ZN(n722) );
  NAND2_X1 U800 ( .A1(G140), .A2(n893), .ZN(n721) );
  NAND2_X1 U801 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U802 ( .A(KEYINPUT34), .B(n723), .ZN(n729) );
  NAND2_X1 U803 ( .A1(G116), .A2(n896), .ZN(n725) );
  NAND2_X1 U804 ( .A1(G128), .A2(n897), .ZN(n724) );
  NAND2_X1 U805 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U806 ( .A(KEYINPUT94), .B(n726), .Z(n727) );
  XNOR2_X1 U807 ( .A(KEYINPUT35), .B(n727), .ZN(n728) );
  NOR2_X1 U808 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U809 ( .A(KEYINPUT36), .B(n730), .ZN(n910) );
  XNOR2_X1 U810 ( .A(G2067), .B(KEYINPUT37), .ZN(n765) );
  NOR2_X1 U811 ( .A1(n910), .A2(n765), .ZN(n925) );
  NAND2_X1 U812 ( .A1(n925), .A2(n767), .ZN(n731) );
  XOR2_X1 U813 ( .A(KEYINPUT95), .B(n731), .Z(n763) );
  NAND2_X1 U814 ( .A1(n756), .A2(n763), .ZN(n732) );
  XNOR2_X1 U815 ( .A(n732), .B(KEYINPUT99), .ZN(n734) );
  XNOR2_X1 U816 ( .A(G1986), .B(G290), .ZN(n991) );
  NAND2_X1 U817 ( .A1(n767), .A2(n991), .ZN(n733) );
  NAND2_X1 U818 ( .A1(n734), .A2(n733), .ZN(n755) );
  INV_X1 U819 ( .A(n755), .ZN(n735) );
  NAND2_X1 U820 ( .A1(n972), .A2(n735), .ZN(n736) );
  NOR2_X1 U821 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U822 ( .A1(n739), .A2(n738), .ZN(n773) );
  AND2_X1 U823 ( .A1(n740), .A2(n751), .ZN(n741) );
  NAND2_X1 U824 ( .A1(n742), .A2(n741), .ZN(n747) );
  INV_X1 U825 ( .A(n751), .ZN(n745) );
  NOR2_X1 U826 ( .A1(G2090), .A2(G303), .ZN(n743) );
  NAND2_X1 U827 ( .A1(G8), .A2(n743), .ZN(n744) );
  OR2_X1 U828 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U829 ( .A1(n747), .A2(n746), .ZN(n753) );
  NOR2_X1 U830 ( .A1(G1981), .A2(G305), .ZN(n748) );
  XOR2_X1 U831 ( .A(n748), .B(KEYINPUT24), .Z(n749) );
  XNOR2_X1 U832 ( .A(KEYINPUT100), .B(n749), .ZN(n750) );
  NOR2_X1 U833 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U834 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U835 ( .A1(n755), .A2(n754), .ZN(n771) );
  NOR2_X1 U836 ( .A1(G1996), .A2(n906), .ZN(n929) );
  INV_X1 U837 ( .A(n756), .ZN(n759) );
  NOR2_X1 U838 ( .A1(G1986), .A2(G290), .ZN(n757) );
  NOR2_X1 U839 ( .A1(G1991), .A2(n879), .ZN(n932) );
  NOR2_X1 U840 ( .A1(n757), .A2(n932), .ZN(n758) );
  NOR2_X1 U841 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U842 ( .A1(n929), .A2(n760), .ZN(n762) );
  XOR2_X1 U843 ( .A(KEYINPUT111), .B(KEYINPUT39), .Z(n761) );
  XNOR2_X1 U844 ( .A(n762), .B(n761), .ZN(n764) );
  NAND2_X1 U845 ( .A1(n764), .A2(n763), .ZN(n766) );
  NAND2_X1 U846 ( .A1(n910), .A2(n765), .ZN(n926) );
  NAND2_X1 U847 ( .A1(n766), .A2(n926), .ZN(n768) );
  NAND2_X1 U848 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U849 ( .A(KEYINPUT112), .B(n769), .Z(n770) );
  NOR2_X1 U850 ( .A1(n771), .A2(n770), .ZN(n772) );
  AND2_X1 U851 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U852 ( .A(n775), .B(n774), .ZN(G329) );
  NAND2_X1 U853 ( .A1(G7), .A2(G661), .ZN(n776) );
  XNOR2_X1 U854 ( .A(n776), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U855 ( .A(G223), .ZN(n845) );
  NAND2_X1 U856 ( .A1(n845), .A2(G567), .ZN(n777) );
  XOR2_X1 U857 ( .A(KEYINPUT11), .B(n777), .Z(G234) );
  INV_X1 U858 ( .A(G860), .ZN(n804) );
  OR2_X1 U859 ( .A1(n975), .A2(n804), .ZN(G153) );
  INV_X1 U860 ( .A(G171), .ZN(G301) );
  NOR2_X1 U861 ( .A1(n985), .A2(G868), .ZN(n778) );
  XNOR2_X1 U862 ( .A(n778), .B(KEYINPUT73), .ZN(n780) );
  NAND2_X1 U863 ( .A1(G868), .A2(G301), .ZN(n779) );
  NAND2_X1 U864 ( .A1(n780), .A2(n779), .ZN(G284) );
  XOR2_X1 U865 ( .A(n980), .B(KEYINPUT70), .Z(G299) );
  NOR2_X1 U866 ( .A1(G299), .A2(G868), .ZN(n783) );
  INV_X1 U867 ( .A(G868), .ZN(n781) );
  NOR2_X1 U868 ( .A1(G286), .A2(n781), .ZN(n782) );
  NOR2_X1 U869 ( .A1(n783), .A2(n782), .ZN(G297) );
  NAND2_X1 U870 ( .A1(G559), .A2(n804), .ZN(n784) );
  XOR2_X1 U871 ( .A(KEYINPUT77), .B(n784), .Z(n785) );
  NAND2_X1 U872 ( .A1(n785), .A2(n985), .ZN(n786) );
  XNOR2_X1 U873 ( .A(n786), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U874 ( .A1(G868), .A2(n975), .ZN(n787) );
  XNOR2_X1 U875 ( .A(KEYINPUT78), .B(n787), .ZN(n790) );
  NAND2_X1 U876 ( .A1(G868), .A2(n985), .ZN(n788) );
  NOR2_X1 U877 ( .A1(G559), .A2(n788), .ZN(n789) );
  NOR2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U879 ( .A(KEYINPUT79), .B(n791), .Z(G282) );
  NAND2_X1 U880 ( .A1(G99), .A2(n892), .ZN(n793) );
  NAND2_X1 U881 ( .A1(G111), .A2(n896), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U883 ( .A(KEYINPUT80), .B(n794), .ZN(n799) );
  NAND2_X1 U884 ( .A1(n897), .A2(G123), .ZN(n795) );
  XNOR2_X1 U885 ( .A(n795), .B(KEYINPUT18), .ZN(n797) );
  NAND2_X1 U886 ( .A1(G135), .A2(n893), .ZN(n796) );
  NAND2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U888 ( .A1(n799), .A2(n798), .ZN(n931) );
  XNOR2_X1 U889 ( .A(G2096), .B(n931), .ZN(n801) );
  INV_X1 U890 ( .A(G2100), .ZN(n800) );
  NAND2_X1 U891 ( .A1(n801), .A2(n800), .ZN(G156) );
  XOR2_X1 U892 ( .A(KEYINPUT82), .B(KEYINPUT85), .Z(n806) );
  XNOR2_X1 U893 ( .A(n975), .B(KEYINPUT81), .ZN(n803) );
  NAND2_X1 U894 ( .A1(n985), .A2(G559), .ZN(n802) );
  XNOR2_X1 U895 ( .A(n803), .B(n802), .ZN(n826) );
  NAND2_X1 U896 ( .A1(n826), .A2(n804), .ZN(n805) );
  XNOR2_X1 U897 ( .A(n806), .B(n805), .ZN(n819) );
  NAND2_X1 U898 ( .A1(G93), .A2(n807), .ZN(n810) );
  NAND2_X1 U899 ( .A1(G80), .A2(n808), .ZN(n809) );
  NAND2_X1 U900 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U901 ( .A(n811), .B(KEYINPUT83), .ZN(n814) );
  NAND2_X1 U902 ( .A1(G55), .A2(n812), .ZN(n813) );
  NAND2_X1 U903 ( .A1(n814), .A2(n813), .ZN(n818) );
  NAND2_X1 U904 ( .A1(n815), .A2(G67), .ZN(n816) );
  XOR2_X1 U905 ( .A(KEYINPUT84), .B(n816), .Z(n817) );
  NOR2_X1 U906 ( .A1(n818), .A2(n817), .ZN(n828) );
  XOR2_X1 U907 ( .A(n819), .B(n828), .Z(G145) );
  XNOR2_X1 U908 ( .A(KEYINPUT19), .B(G303), .ZN(n820) );
  XNOR2_X1 U909 ( .A(n820), .B(G288), .ZN(n821) );
  XNOR2_X1 U910 ( .A(KEYINPUT90), .B(n821), .ZN(n823) );
  XNOR2_X1 U911 ( .A(G305), .B(G290), .ZN(n822) );
  XNOR2_X1 U912 ( .A(n823), .B(n822), .ZN(n825) );
  XOR2_X1 U913 ( .A(n828), .B(G299), .Z(n824) );
  XNOR2_X1 U914 ( .A(n825), .B(n824), .ZN(n915) );
  XNOR2_X1 U915 ( .A(n915), .B(n826), .ZN(n827) );
  NAND2_X1 U916 ( .A1(n827), .A2(G868), .ZN(n830) );
  OR2_X1 U917 ( .A1(G868), .A2(n828), .ZN(n829) );
  NAND2_X1 U918 ( .A1(n830), .A2(n829), .ZN(G295) );
  NAND2_X1 U919 ( .A1(G2078), .A2(G2084), .ZN(n831) );
  XNOR2_X1 U920 ( .A(n831), .B(KEYINPUT91), .ZN(n832) );
  XNOR2_X1 U921 ( .A(n832), .B(KEYINPUT20), .ZN(n833) );
  NAND2_X1 U922 ( .A1(n833), .A2(G2090), .ZN(n834) );
  XNOR2_X1 U923 ( .A(KEYINPUT21), .B(n834), .ZN(n835) );
  NAND2_X1 U924 ( .A1(n835), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U925 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U926 ( .A1(G220), .A2(G219), .ZN(n836) );
  XOR2_X1 U927 ( .A(KEYINPUT22), .B(n836), .Z(n837) );
  NOR2_X1 U928 ( .A1(G218), .A2(n837), .ZN(n838) );
  NAND2_X1 U929 ( .A1(G96), .A2(n838), .ZN(n849) );
  NAND2_X1 U930 ( .A1(n849), .A2(G2106), .ZN(n843) );
  NOR2_X1 U931 ( .A1(G236), .A2(G238), .ZN(n840) );
  NOR2_X1 U932 ( .A1(G235), .A2(G237), .ZN(n839) );
  NAND2_X1 U933 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U934 ( .A(KEYINPUT92), .B(n841), .ZN(n850) );
  NAND2_X1 U935 ( .A1(n850), .A2(G567), .ZN(n842) );
  NAND2_X1 U936 ( .A1(n843), .A2(n842), .ZN(n851) );
  NAND2_X1 U937 ( .A1(G661), .A2(G483), .ZN(n844) );
  NOR2_X1 U938 ( .A1(n851), .A2(n844), .ZN(n848) );
  NAND2_X1 U939 ( .A1(n848), .A2(G36), .ZN(G176) );
  NAND2_X1 U940 ( .A1(G2106), .A2(n845), .ZN(G217) );
  AND2_X1 U941 ( .A1(G15), .A2(G2), .ZN(n846) );
  NAND2_X1 U942 ( .A1(G661), .A2(n846), .ZN(G259) );
  NAND2_X1 U943 ( .A1(G3), .A2(G1), .ZN(n847) );
  NAND2_X1 U944 ( .A1(n848), .A2(n847), .ZN(G188) );
  INV_X1 U946 ( .A(G96), .ZN(G221) );
  NOR2_X1 U947 ( .A1(n850), .A2(n849), .ZN(G325) );
  INV_X1 U948 ( .A(G325), .ZN(G261) );
  INV_X1 U949 ( .A(n851), .ZN(G319) );
  XOR2_X1 U950 ( .A(G2096), .B(KEYINPUT114), .Z(n853) );
  XNOR2_X1 U951 ( .A(G2090), .B(KEYINPUT43), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U953 ( .A(n854), .B(KEYINPUT42), .Z(n856) );
  XNOR2_X1 U954 ( .A(G2072), .B(G2067), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U956 ( .A(G2678), .B(G2100), .Z(n858) );
  XNOR2_X1 U957 ( .A(G2078), .B(G2084), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(G227) );
  XOR2_X1 U960 ( .A(G1991), .B(G1976), .Z(n862) );
  XNOR2_X1 U961 ( .A(G1966), .B(G1981), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U963 ( .A(G1986), .B(G1971), .Z(n864) );
  XNOR2_X1 U964 ( .A(G1961), .B(G1956), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U966 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U967 ( .A(KEYINPUT115), .B(G2474), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U969 ( .A(KEYINPUT41), .B(n869), .ZN(n870) );
  XOR2_X1 U970 ( .A(n870), .B(G1996), .Z(G229) );
  NAND2_X1 U971 ( .A1(n893), .A2(G136), .ZN(n871) );
  XNOR2_X1 U972 ( .A(n871), .B(KEYINPUT116), .ZN(n874) );
  NAND2_X1 U973 ( .A1(G124), .A2(n897), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n872), .B(KEYINPUT44), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n878) );
  NAND2_X1 U976 ( .A1(G100), .A2(n892), .ZN(n876) );
  NAND2_X1 U977 ( .A1(G112), .A2(n896), .ZN(n875) );
  NAND2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U979 ( .A1(n878), .A2(n877), .ZN(G162) );
  XNOR2_X1 U980 ( .A(KEYINPUT48), .B(KEYINPUT118), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n879), .B(KEYINPUT46), .ZN(n880) );
  XNOR2_X1 U982 ( .A(n881), .B(n880), .ZN(n891) );
  NAND2_X1 U983 ( .A1(G118), .A2(n896), .ZN(n883) );
  NAND2_X1 U984 ( .A1(G130), .A2(n897), .ZN(n882) );
  NAND2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n889) );
  NAND2_X1 U986 ( .A1(G142), .A2(n893), .ZN(n884) );
  XOR2_X1 U987 ( .A(KEYINPUT117), .B(n884), .Z(n886) );
  NAND2_X1 U988 ( .A1(n892), .A2(G106), .ZN(n885) );
  NAND2_X1 U989 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U990 ( .A(KEYINPUT45), .B(n887), .Z(n888) );
  NOR2_X1 U991 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U992 ( .A(n891), .B(n890), .Z(n904) );
  NAND2_X1 U993 ( .A1(G103), .A2(n892), .ZN(n895) );
  NAND2_X1 U994 ( .A1(G139), .A2(n893), .ZN(n894) );
  NAND2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n902) );
  NAND2_X1 U996 ( .A1(G115), .A2(n896), .ZN(n899) );
  NAND2_X1 U997 ( .A1(G127), .A2(n897), .ZN(n898) );
  NAND2_X1 U998 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U999 ( .A(KEYINPUT47), .B(n900), .Z(n901) );
  NOR2_X1 U1000 ( .A1(n902), .A2(n901), .ZN(n938) );
  XNOR2_X1 U1001 ( .A(G164), .B(n938), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n905), .B(G160), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(G162), .B(n931), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n911) );
  XOR2_X1 U1007 ( .A(n911), .B(n910), .Z(n912) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n912), .ZN(G395) );
  XNOR2_X1 U1009 ( .A(n975), .B(G286), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(G171), .B(n985), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(n914), .B(n913), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(n916), .B(n915), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n917), .ZN(G397) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(KEYINPUT119), .B(KEYINPUT49), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(n919), .B(n918), .ZN(n922) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(n920), .B(KEYINPUT120), .ZN(n921) );
  NAND2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1020 ( .A1(G401), .A2(n923), .ZN(n924) );
  NAND2_X1 U1021 ( .A1(G319), .A2(n924), .ZN(G225) );
  INV_X1 U1022 ( .A(G225), .ZN(G308) );
  INV_X1 U1023 ( .A(n925), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n947) );
  XOR2_X1 U1025 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1027 ( .A(KEYINPUT51), .B(n930), .Z(n945) );
  XNOR2_X1 U1028 ( .A(G2084), .B(G160), .ZN(n937) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(KEYINPUT121), .B(n933), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n943) );
  XOR2_X1 U1033 ( .A(G2072), .B(n938), .Z(n940) );
  XOR2_X1 U1034 ( .A(G164), .B(G2078), .Z(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1036 ( .A(KEYINPUT50), .B(n941), .Z(n942) );
  NOR2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(KEYINPUT52), .B(n948), .ZN(n950) );
  INV_X1 U1041 ( .A(KEYINPUT55), .ZN(n949) );
  NAND2_X1 U1042 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1043 ( .A1(n951), .A2(G29), .ZN(n1030) );
  XOR2_X1 U1044 ( .A(G29), .B(KEYINPUT122), .Z(n970) );
  XNOR2_X1 U1045 ( .A(G2072), .B(G33), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(G2067), .B(G26), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n961) );
  XOR2_X1 U1048 ( .A(G1991), .B(G25), .Z(n954) );
  NAND2_X1 U1049 ( .A1(n954), .A2(G28), .ZN(n959) );
  XOR2_X1 U1050 ( .A(G1996), .B(G32), .Z(n957) );
  XNOR2_X1 U1051 ( .A(n955), .B(G27), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(n962), .B(KEYINPUT53), .ZN(n965) );
  XOR2_X1 U1056 ( .A(G2084), .B(KEYINPUT54), .Z(n963) );
  XNOR2_X1 U1057 ( .A(G34), .B(n963), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(G35), .B(G2090), .ZN(n966) );
  NOR2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(n968), .B(KEYINPUT55), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(G11), .A2(n971), .ZN(n1028) );
  XNOR2_X1 U1064 ( .A(G16), .B(KEYINPUT56), .ZN(n998) );
  XNOR2_X1 U1065 ( .A(G1966), .B(G168), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n974), .B(KEYINPUT57), .ZN(n996) );
  XNOR2_X1 U1068 ( .A(G1341), .B(KEYINPUT124), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(n976), .B(n975), .ZN(n994) );
  INV_X1 U1070 ( .A(n977), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(G166), .B(G1971), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(n980), .B(G1956), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n989) );
  XOR2_X1 U1076 ( .A(G1348), .B(n985), .Z(n987) );
  XOR2_X1 U1077 ( .A(G171), .B(G1961), .Z(n986) );
  NOR2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(n992), .B(KEYINPUT123), .ZN(n993) );
  NOR2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n1026) );
  INV_X1 U1085 ( .A(G16), .ZN(n1024) );
  XNOR2_X1 U1086 ( .A(G20), .B(n999), .ZN(n1003) );
  XNOR2_X1 U1087 ( .A(G1341), .B(G19), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(G6), .B(G1981), .ZN(n1000) );
  NOR2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1006) );
  XOR2_X1 U1091 ( .A(KEYINPUT59), .B(G1348), .Z(n1004) );
  XNOR2_X1 U1092 ( .A(G4), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(KEYINPUT60), .B(n1007), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(n1008), .B(G5), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1021) );
  XOR2_X1 U1097 ( .A(G1966), .B(G21), .Z(n1019) );
  XOR2_X1 U1098 ( .A(G1971), .B(G22), .Z(n1013) );
  XOR2_X1 U1099 ( .A(G24), .B(KEYINPUT126), .Z(n1011) );
  XNOR2_X1 U1100 ( .A(n1011), .B(G1986), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1016) );
  XOR2_X1 U1102 ( .A(KEYINPUT125), .B(G1976), .Z(n1014) );
  XNOR2_X1 U1103 ( .A(G23), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(n1017), .B(KEYINPUT58), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(KEYINPUT61), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1112 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1113 ( .A(n1031), .B(KEYINPUT127), .ZN(n1032) );
  XNOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1032), .ZN(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

