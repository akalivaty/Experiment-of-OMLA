//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1161, new_n1162, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT65), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n217), .A2(new_n218), .ZN(new_n220));
  AOI211_X1 g0020(.A(new_n219), .B(new_n220), .C1(G77), .C2(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G226), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n202), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G116), .ZN(new_n226));
  INV_X1    g0026(.A(G270), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n208), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(G50), .B1(G58), .B2(G68), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n211), .B(new_n230), .C1(new_n233), .C2(new_n235), .ZN(G361));
  XOR2_X1   g0036(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G358));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  INV_X1    g0046(.A(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(KEYINPUT67), .B(G50), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n251), .B(new_n252), .Z(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(KEYINPUT68), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G41), .A2(G45), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n255), .B1(new_n256), .B2(G1), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G1), .A3(G13), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n260), .B(KEYINPUT68), .C1(G41), .C2(G45), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n257), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(new_n262), .B(KEYINPUT69), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G226), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n259), .A2(KEYINPUT70), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT70), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n258), .A2(new_n270), .A3(G1), .A4(G13), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G223), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G1698), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n276), .B1(G222), .B2(G1698), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n273), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n205), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n268), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n265), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G169), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n231), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OR2_X1    g0091(.A1(new_n291), .A2(KEYINPUT71), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(KEYINPUT71), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n260), .A2(G20), .ZN(new_n294));
  AND3_X1   g0094(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G50), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n204), .A2(new_n232), .ZN(new_n297));
  XNOR2_X1  g0097(.A(KEYINPUT8), .B(G58), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n232), .A2(G33), .ZN(new_n299));
  INV_X1    g0099(.A(G150), .ZN(new_n300));
  NOR2_X1   g0100(.A1(G20), .A2(G33), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  OAI22_X1  g0102(.A1(new_n298), .A2(new_n299), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n288), .B1(new_n297), .B2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n296), .B(new_n304), .C1(G50), .C2(new_n290), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n286), .B(new_n305), .C1(G179), .C2(new_n284), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n284), .A2(G200), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT74), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n305), .B(KEYINPUT9), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n265), .A2(new_n283), .A3(G190), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  OR2_X1    g0112(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n307), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G1698), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n222), .A2(new_n316), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n274), .B(new_n317), .C1(G232), .C2(new_n316), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G33), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(new_n215), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n272), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n268), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n322), .B(new_n323), .C1(new_n263), .C2(new_n224), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT13), .ZN(new_n325));
  INV_X1    g0125(.A(G190), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n302), .A2(new_n202), .B1(new_n232), .B2(G68), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n299), .A2(new_n205), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n288), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT11), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n289), .A2(G68), .A3(new_n294), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT12), .ZN(new_n333));
  INV_X1    g0133(.A(new_n290), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n333), .B1(new_n334), .B2(new_n223), .ZN(new_n335));
  NOR3_X1   g0135(.A1(new_n290), .A2(KEYINPUT12), .A3(G68), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n331), .B(new_n332), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n327), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n325), .A2(G200), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT75), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n325), .A2(KEYINPUT75), .A3(G200), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n338), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT76), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n325), .A2(new_n344), .A3(KEYINPUT14), .A4(G169), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n345), .A2(new_n337), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n325), .A2(new_n344), .A3(G169), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT14), .ZN(new_n348));
  INV_X1    g0148(.A(G179), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n347), .B(new_n348), .C1(new_n349), .C2(new_n325), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n274), .A2(G232), .A3(new_n316), .ZN(new_n352));
  XOR2_X1   g0152(.A(new_n352), .B(KEYINPUT72), .Z(new_n353));
  NAND2_X1  g0153(.A1(new_n274), .A2(G1698), .ZN(new_n354));
  INV_X1    g0154(.A(G107), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n354), .A2(new_n224), .B1(new_n355), .B2(new_n274), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n272), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n264), .A2(G244), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n357), .A2(new_n358), .A3(new_n323), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G200), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XOR2_X1   g0162(.A(KEYINPUT15), .B(G87), .Z(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(new_n299), .ZN(new_n365));
  OAI22_X1  g0165(.A1(new_n298), .A2(new_n302), .B1(new_n232), .B2(new_n205), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n288), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n289), .A2(G77), .A3(new_n294), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n367), .B(new_n368), .C1(G77), .C2(new_n290), .ZN(new_n369));
  XOR2_X1   g0169(.A(new_n369), .B(KEYINPUT73), .Z(new_n370));
  NOR2_X1   g0170(.A1(new_n362), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n326), .B2(new_n359), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n315), .A2(new_n343), .A3(new_n351), .A4(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT80), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G87), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT78), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n275), .A2(new_n316), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n222), .A2(G1698), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n377), .B(new_n378), .C1(new_n279), .C2(new_n280), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n268), .B1(new_n380), .B2(new_n272), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n257), .A2(new_n259), .A3(G232), .A4(new_n261), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n382), .A2(KEYINPUT79), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(KEYINPUT79), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n381), .B(new_n326), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  XNOR2_X1  g0186(.A(new_n382), .B(KEYINPUT79), .ZN(new_n387));
  AOI21_X1  g0187(.A(G200), .B1(new_n387), .B2(new_n381), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n374), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n361), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(KEYINPUT80), .A3(new_n385), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT7), .B1(new_n281), .B2(new_n232), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  NOR4_X1   g0195(.A1(new_n279), .A2(new_n280), .A3(new_n395), .A4(G20), .ZN(new_n396));
  OAI21_X1  g0196(.A(G68), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n301), .A2(G159), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G58), .A2(G68), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT77), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n399), .B(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(G20), .B1(new_n401), .B2(new_n201), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n397), .A2(new_n398), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT16), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n397), .A2(KEYINPUT16), .A3(new_n398), .A4(new_n402), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n288), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n298), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n295), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n298), .A2(new_n334), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n407), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  XNOR2_X1  g0211(.A(KEYINPUT81), .B(KEYINPUT17), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n393), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n407), .A2(new_n409), .A3(new_n410), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n389), .B2(new_n392), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT17), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT81), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n413), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n360), .A2(new_n349), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n359), .A2(new_n285), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n370), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n390), .A2(new_n285), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n387), .A2(new_n349), .A3(new_n381), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n414), .A2(KEYINPUT18), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT18), .B1(new_n414), .B2(new_n426), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OR3_X1    g0229(.A1(new_n418), .A2(new_n422), .A3(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n373), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n334), .A2(new_n288), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n260), .A2(G33), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(new_n355), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n274), .A2(new_n232), .A3(G87), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT22), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n355), .A2(G20), .ZN(new_n438));
  OAI22_X1  g0238(.A1(KEYINPUT23), .A2(new_n438), .B1(new_n299), .B2(new_n226), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(KEYINPUT23), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n440), .A2(KEYINPUT88), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(KEYINPUT88), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT24), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT24), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n437), .A2(new_n446), .A3(new_n443), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n435), .B1(new_n448), .B2(new_n288), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n290), .A2(G107), .ZN(new_n450));
  XNOR2_X1  g0250(.A(new_n450), .B(KEYINPUT25), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n274), .A2(G257), .A3(G1698), .ZN(new_n452));
  INV_X1    g0252(.A(G294), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n274), .A2(new_n316), .ZN(new_n454));
  OAI221_X1 g0254(.A(new_n452), .B1(new_n320), .B2(new_n453), .C1(new_n454), .C2(new_n214), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n272), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT83), .ZN(new_n457));
  INV_X1    g0257(.A(G41), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(KEYINPUT5), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n260), .A2(G45), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(KEYINPUT5), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT5), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G41), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n464), .A2(KEYINPUT83), .A3(new_n260), .A4(G45), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n461), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(G264), .A3(new_n259), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n461), .A2(new_n465), .A3(G274), .A4(new_n462), .ZN(new_n468));
  INV_X1    g0268(.A(new_n259), .ZN(new_n469));
  OR2_X1    g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n456), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n471), .A2(new_n326), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(G200), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n449), .A2(new_n451), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n437), .A2(new_n446), .A3(new_n443), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n446), .B1(new_n437), .B2(new_n443), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n288), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n435), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n477), .A2(new_n478), .A3(new_n451), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT89), .B1(new_n471), .B2(G169), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n456), .A2(new_n467), .A3(G179), .A4(new_n470), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n481), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT89), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n479), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n474), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n434), .A2(new_n215), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n290), .A2(G97), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(G107), .B1(new_n394), .B2(new_n396), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT6), .ZN(new_n491));
  AND2_X1   g0291(.A1(G97), .A2(G107), .ZN(new_n492));
  NOR2_X1   g0292(.A1(G97), .A2(G107), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n355), .A2(KEYINPUT6), .A3(G97), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n496), .A2(G20), .B1(G77), .B2(new_n301), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n289), .B1(new_n490), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(KEYINPUT82), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT82), .ZN(new_n500));
  AOI211_X1 g0300(.A(new_n500), .B(new_n289), .C1(new_n490), .C2(new_n497), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n489), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(G244), .B(new_n316), .C1(new_n279), .C2(new_n280), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT4), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n274), .A2(KEYINPUT4), .A3(G244), .A4(new_n316), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G283), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n354), .B2(new_n214), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n272), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n466), .A2(G257), .A3(new_n259), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n470), .A3(new_n511), .ZN(new_n512));
  OR2_X1    g0312(.A1(new_n512), .A2(G179), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n502), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT84), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n505), .A2(new_n506), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n281), .A2(new_n316), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n517), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n273), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n511), .B1(new_n469), .B2(new_n468), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n510), .A2(new_n470), .A3(KEYINPUT84), .A4(new_n511), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n521), .A2(new_n285), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n512), .A2(G200), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n524), .B(new_n489), .C1(new_n499), .C2(new_n501), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n326), .B1(new_n521), .B2(new_n522), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n514), .A2(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT85), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n521), .A2(new_n522), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G190), .ZN(new_n530));
  INV_X1    g0330(.A(new_n502), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n531), .A3(new_n524), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT85), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n502), .B(new_n513), .C1(new_n529), .C2(G169), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g0336(.A(KEYINPUT86), .B(G87), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n493), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n538), .B(KEYINPUT19), .C1(G20), .C2(new_n321), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n274), .A2(new_n232), .A3(G68), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n299), .A2(new_n215), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n539), .B(new_n540), .C1(KEYINPUT19), .C2(new_n541), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n542), .A2(new_n288), .B1(new_n334), .B2(new_n364), .ZN(new_n543));
  INV_X1    g0343(.A(new_n434), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n363), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n224), .A2(new_n316), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n274), .B(new_n547), .C1(G244), .C2(new_n316), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G116), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n272), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n259), .A2(G250), .A3(new_n460), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n267), .B2(new_n460), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n285), .ZN(new_n556));
  INV_X1    g0356(.A(new_n555), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n349), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n546), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n555), .A2(G200), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n551), .A2(G190), .A3(new_n554), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n544), .A2(G87), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n543), .A2(new_n560), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n508), .B(new_n232), .C1(G33), .C2(new_n215), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n565), .B(new_n288), .C1(new_n232), .C2(G116), .ZN(new_n566));
  XOR2_X1   g0366(.A(new_n566), .B(KEYINPUT20), .Z(new_n567));
  NAND2_X1  g0367(.A1(new_n334), .A2(new_n226), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT87), .B1(new_n434), .B2(new_n226), .ZN(new_n569));
  OR3_X1    g0369(.A1(new_n434), .A2(KEYINPUT87), .A3(new_n226), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n567), .A2(new_n568), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n274), .A2(G264), .A3(G1698), .ZN(new_n572));
  INV_X1    g0372(.A(G303), .ZN(new_n573));
  OAI221_X1 g0373(.A(new_n572), .B1(new_n573), .B2(new_n274), .C1(new_n454), .C2(new_n216), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n272), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n466), .A2(new_n259), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n575), .B(new_n470), .C1(new_n227), .C2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n571), .A2(new_n577), .A3(G169), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT21), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT21), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n571), .A2(new_n577), .A3(new_n580), .A4(G169), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n571), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n583), .A2(new_n349), .ZN(new_n584));
  INV_X1    g0384(.A(new_n577), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n577), .A2(G200), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n587), .B(new_n583), .C1(new_n326), .C2(new_n577), .ZN(new_n588));
  AND4_X1   g0388(.A1(new_n564), .A2(new_n582), .A3(new_n586), .A4(new_n588), .ZN(new_n589));
  AND4_X1   g0389(.A1(new_n431), .A2(new_n486), .A3(new_n536), .A4(new_n589), .ZN(G372));
  AOI22_X1  g0390(.A1(new_n579), .A2(new_n581), .B1(new_n584), .B2(new_n585), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n485), .ZN(new_n592));
  INV_X1    g0392(.A(new_n527), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n543), .A2(new_n562), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n550), .A2(KEYINPUT90), .A3(new_n272), .ZN(new_n596));
  AOI21_X1  g0396(.A(KEYINPUT90), .B1(new_n550), .B2(new_n272), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n554), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n595), .B(new_n561), .C1(new_n361), .C2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n592), .A2(new_n474), .A3(new_n593), .A4(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n546), .B(new_n558), .C1(new_n599), .C2(G169), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  OR3_X1    g0403(.A1(new_n603), .A2(KEYINPUT26), .A3(new_n534), .ZN(new_n604));
  INV_X1    g0404(.A(new_n534), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n564), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT26), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n601), .A2(new_n604), .A3(new_n602), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n431), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n429), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n343), .A2(new_n422), .B1(new_n346), .B2(new_n350), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n610), .B1(new_n611), .B2(new_n418), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n313), .A2(new_n314), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n609), .A2(new_n306), .A3(new_n614), .ZN(G369));
  INV_X1    g0415(.A(G13), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n616), .A2(G20), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  OR3_X1    g0418(.A1(new_n618), .A2(KEYINPUT27), .A3(G1), .ZN(new_n619));
  OAI21_X1  g0419(.A(KEYINPUT27), .B1(new_n618), .B2(G1), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(G213), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(G343), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n479), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n486), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT91), .ZN(new_n626));
  XNOR2_X1  g0426(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n623), .ZN(new_n628));
  OR2_X1    g0428(.A1(new_n485), .A2(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n591), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n583), .A2(new_n628), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n591), .A2(new_n588), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n633), .B1(new_n634), .B2(new_n632), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(G330), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n591), .A2(new_n623), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n627), .A2(new_n639), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n485), .A2(new_n623), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n637), .A2(new_n642), .ZN(G399));
  INV_X1    g0443(.A(KEYINPUT92), .ZN(new_n644));
  INV_X1    g0444(.A(new_n209), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(G41), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n209), .A2(KEYINPUT92), .A3(new_n458), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n537), .A2(new_n226), .A3(new_n493), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n648), .A2(G1), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n234), .B2(new_n648), .ZN(new_n652));
  XOR2_X1   g0452(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n653));
  XNOR2_X1  g0453(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n601), .A2(new_n602), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT26), .B1(new_n603), .B2(new_n534), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(KEYINPUT26), .B2(new_n606), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n628), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT29), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n608), .A2(new_n628), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(KEYINPUT29), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G330), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n576), .A2(new_n227), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n272), .B2(new_n574), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n529), .A2(new_n483), .A3(new_n557), .A4(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT30), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n555), .B1(new_n521), .B2(new_n522), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n668), .A2(KEYINPUT30), .A3(new_n483), .A4(new_n664), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n577), .A2(new_n512), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n670), .A2(new_n349), .A3(new_n598), .A4(new_n471), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n667), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n672), .A2(KEYINPUT31), .A3(new_n623), .ZN(new_n673));
  AOI21_X1  g0473(.A(KEYINPUT31), .B1(new_n672), .B2(new_n623), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n536), .A2(new_n589), .A3(new_n486), .A4(new_n628), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n662), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n661), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n654), .B1(new_n678), .B2(G1), .ZN(new_n679));
  XOR2_X1   g0479(.A(new_n679), .B(KEYINPUT94), .Z(G364));
  NOR2_X1   g0480(.A1(new_n645), .A2(new_n274), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n250), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n682), .B1(new_n683), .B2(G45), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(G45), .B2(new_n234), .ZN(new_n685));
  INV_X1    g0485(.A(G355), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n645), .A2(new_n281), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT95), .ZN(new_n688));
  OAI221_X1 g0488(.A(new_n685), .B1(G116), .B2(new_n209), .C1(new_n686), .C2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(G13), .A2(G33), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT96), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G20), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n231), .B1(G20), .B2(new_n285), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n232), .A2(G190), .ZN(new_n697));
  NOR2_X1   g0497(.A1(G179), .A2(G200), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G159), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n349), .A2(G200), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n697), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n702), .A2(KEYINPUT32), .B1(G77), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT32), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n232), .B1(new_n698), .B2(G190), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n701), .A2(new_n707), .B1(new_n709), .B2(G97), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n232), .A2(new_n326), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n703), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G58), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n706), .A2(new_n274), .A3(new_n710), .A4(new_n714), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n232), .A2(new_n349), .A3(new_n361), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT97), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(new_n717), .A3(new_n326), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n717), .B1(new_n716), .B2(new_n326), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n361), .A2(G179), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n697), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n721), .A2(G68), .B1(G107), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n711), .A2(new_n722), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n537), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n716), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n326), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n715), .B(new_n727), .C1(G50), .C2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n699), .ZN(new_n731));
  AOI22_X1  g0531(.A1(G311), .A2(new_n705), .B1(new_n731), .B2(G329), .ZN(new_n732));
  INV_X1    g0532(.A(new_n726), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n733), .A2(G303), .B1(new_n709), .B2(G294), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n732), .A2(new_n734), .A3(new_n281), .ZN(new_n735));
  INV_X1    g0535(.A(G283), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n723), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g0537(.A(KEYINPUT33), .B(G317), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n737), .B1(new_n721), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G326), .ZN(new_n740));
  INV_X1    g0540(.A(new_n729), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI211_X1 g0542(.A(new_n735), .B(new_n742), .C1(G322), .C2(new_n713), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n694), .B1(new_n730), .B2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n648), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n260), .B1(new_n617), .B2(G45), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n696), .A2(new_n744), .A3(new_n748), .ZN(new_n749));
  XOR2_X1   g0549(.A(new_n749), .B(KEYINPUT98), .Z(new_n750));
  INV_X1    g0550(.A(new_n693), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n750), .B1(new_n635), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n748), .B1(new_n635), .B2(G330), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G330), .B2(new_n635), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(G396));
  INV_X1    g0556(.A(G311), .ZN(new_n757));
  INV_X1    g0557(.A(new_n721), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n281), .B1(new_n757), .B2(new_n699), .C1(new_n758), .C2(new_n736), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n713), .A2(G294), .B1(new_n709), .B2(G97), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(new_n355), .B2(new_n726), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n761), .B1(G116), .B2(new_n705), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(new_n573), .B2(new_n741), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n759), .B(new_n763), .C1(G87), .C2(new_n724), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT99), .Z(new_n765));
  AOI22_X1  g0565(.A1(new_n721), .A2(G150), .B1(G137), .B2(new_n729), .ZN(new_n766));
  XNOR2_X1  g0566(.A(KEYINPUT100), .B(G143), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n713), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n766), .B(new_n768), .C1(new_n700), .C2(new_n704), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT34), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n724), .A2(G68), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n202), .B2(new_n726), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n281), .B1(new_n731), .B2(G132), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n774), .B(new_n775), .C1(new_n247), .C2(new_n708), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(new_n770), .B2(new_n769), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n694), .B1(new_n765), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n694), .A2(new_n690), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n205), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n778), .A2(new_n748), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n370), .A2(new_n623), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n422), .B1(new_n372), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n421), .A2(new_n623), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n781), .B1(new_n691), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n660), .B(new_n785), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n677), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT101), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n748), .B1(new_n788), .B2(new_n677), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n787), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(G384));
  NAND2_X1  g0593(.A1(new_n337), .A2(new_n623), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n351), .A2(new_n343), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(KEYINPUT102), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n346), .A2(new_n350), .A3(new_n623), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT102), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n351), .A2(new_n798), .A3(new_n343), .A4(new_n794), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n796), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT106), .ZN(new_n801));
  INV_X1    g0601(.A(new_n674), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n672), .A2(KEYINPUT31), .A3(new_n623), .ZN(new_n803));
  AND4_X1   g0603(.A1(new_n801), .A2(new_n676), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n801), .B1(new_n675), .B2(new_n676), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n785), .B(new_n800), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT37), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n393), .A2(new_n411), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT103), .ZN(new_n809));
  INV_X1    g0609(.A(new_n621), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n414), .B1(new_n426), .B2(new_n810), .ZN(new_n811));
  AND3_X1   g0611(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n809), .B1(new_n808), .B2(new_n811), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n807), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n411), .A2(new_n621), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n418), .B2(new_n429), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n407), .A2(new_n410), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n817), .A2(new_n409), .B1(new_n425), .B2(new_n621), .ZN(new_n818));
  OAI21_X1  g0618(.A(KEYINPUT103), .B1(new_n818), .B2(new_n415), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n819), .A2(KEYINPUT37), .A3(new_n820), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n814), .A2(new_n816), .A3(new_n821), .A4(KEYINPUT38), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n818), .A2(new_n415), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n807), .B1(new_n811), .B2(KEYINPUT105), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  AND3_X1   g0626(.A1(new_n825), .A2(new_n816), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n822), .B1(new_n827), .B2(KEYINPUT38), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(KEYINPUT40), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n806), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n676), .A2(new_n802), .A3(new_n803), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(KEYINPUT106), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n675), .A2(new_n801), .A3(new_n676), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n786), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n814), .A2(new_n821), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n836), .A2(KEYINPUT104), .A3(KEYINPUT38), .A4(new_n816), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n814), .A2(new_n816), .A3(new_n821), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT38), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT104), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n840), .A2(new_n841), .A3(new_n822), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n835), .A2(new_n800), .A3(new_n837), .A4(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT40), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT107), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n842), .A2(new_n837), .ZN(new_n846));
  OAI211_X1 g0646(.A(KEYINPUT107), .B(new_n844), .C1(new_n806), .C2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(G330), .B(new_n831), .C1(new_n845), .C2(new_n848), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n430), .B(new_n373), .C1(new_n833), .C2(new_n834), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(G330), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n844), .B1(new_n806), .B2(new_n846), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT107), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n830), .B1(new_n854), .B2(new_n847), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n849), .A2(new_n851), .B1(new_n855), .B2(new_n850), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n660), .A2(new_n783), .B1(new_n421), .B2(new_n623), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n800), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n858), .A2(new_n846), .B1(new_n610), .B2(new_n810), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n351), .A2(new_n623), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OR2_X1    g0661(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n842), .A2(KEYINPUT39), .A3(new_n837), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n856), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n614), .A2(new_n306), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(new_n661), .B2(new_n431), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n867), .A2(new_n869), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n870), .B(new_n871), .C1(new_n260), .C2(new_n617), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n226), .B1(new_n496), .B2(KEYINPUT35), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n873), .B(new_n233), .C1(KEYINPUT35), .C2(new_n496), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(KEYINPUT36), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n401), .A2(new_n205), .A3(new_n234), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n223), .A2(G50), .ZN(new_n877));
  OAI211_X1 g0677(.A(G1), .B(new_n616), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n872), .A2(new_n875), .A3(new_n878), .ZN(G367));
  INV_X1    g0679(.A(new_n678), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n532), .B1(new_n531), .B2(new_n628), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n534), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n534), .A2(new_n623), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n640), .A2(new_n641), .A3(new_n886), .ZN(new_n887));
  XOR2_X1   g0687(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n888));
  XNOR2_X1  g0688(.A(new_n887), .B(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT44), .B1(new_n642), .B2(new_n885), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n642), .A2(KEYINPUT44), .A3(new_n885), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n630), .A2(new_n639), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n640), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n637), .B1(new_n895), .B2(new_n636), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n678), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT109), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT109), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n892), .A2(new_n899), .A3(new_n678), .A4(new_n896), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n880), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  XOR2_X1   g0701(.A(new_n648), .B(KEYINPUT41), .Z(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n746), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n641), .A2(KEYINPUT42), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n642), .A2(new_n886), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n627), .A2(new_n639), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n882), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n883), .B1(new_n908), .B2(KEYINPUT42), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n595), .A2(new_n628), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(new_n602), .A3(new_n600), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n602), .B2(new_n911), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n906), .A2(new_n909), .B1(KEYINPUT43), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n913), .A2(KEYINPUT43), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n914), .B(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n637), .A2(new_n886), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n916), .B(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n904), .A2(new_n918), .ZN(new_n919));
  OAI221_X1 g0719(.A(new_n695), .B1(new_n209), .B2(new_n364), .C1(new_n244), .C2(new_n682), .ZN(new_n920));
  AOI22_X1  g0720(.A1(G50), .A2(new_n705), .B1(new_n731), .B2(G137), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n300), .B2(new_n712), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n721), .A2(G159), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n733), .A2(G58), .B1(new_n709), .B2(G68), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n724), .A2(G77), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n923), .A2(new_n274), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  AOI211_X1 g0726(.A(new_n922), .B(new_n926), .C1(new_n729), .C2(new_n767), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n724), .A2(G97), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n712), .A2(new_n573), .B1(new_n704), .B2(new_n736), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n733), .A2(KEYINPUT46), .A3(G116), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n281), .ZN(new_n931));
  AOI211_X1 g0731(.A(new_n929), .B(new_n931), .C1(G107), .C2(new_n709), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n729), .A2(G311), .B1(G317), .B2(new_n731), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT46), .B1(new_n733), .B2(G116), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(new_n721), .B2(G294), .ZN(new_n935));
  AND3_X1   g0735(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n927), .B1(new_n928), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT47), .ZN(new_n938));
  INV_X1    g0738(.A(new_n694), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n748), .B(new_n920), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n913), .A2(new_n751), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n919), .A2(new_n943), .ZN(G387));
  AOI21_X1  g0744(.A(new_n281), .B1(new_n721), .B2(new_n408), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n945), .B1(new_n202), .B2(new_n712), .C1(new_n364), .C2(new_n708), .ZN(new_n946));
  XOR2_X1   g0746(.A(KEYINPUT112), .B(G150), .Z(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(new_n699), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n726), .A2(new_n205), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n928), .B1(new_n223), .B2(new_n704), .C1(new_n741), .C2(new_n700), .ZN(new_n950));
  NOR4_X1   g0750(.A1(new_n946), .A2(new_n948), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT113), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n721), .A2(G311), .B1(G322), .B2(new_n729), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n573), .B2(new_n704), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(G317), .B2(new_n713), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT115), .Z(new_n956));
  INV_X1    g0756(.A(KEYINPUT48), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n726), .A2(new_n453), .B1(new_n708), .B2(new_n736), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT114), .Z(new_n961));
  NAND3_X1  g0761(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT49), .Z(new_n963));
  OAI221_X1 g0763(.A(new_n281), .B1(new_n699), .B2(new_n740), .C1(new_n226), .C2(new_n723), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT116), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n952), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n694), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n630), .A2(new_n693), .ZN(new_n968));
  INV_X1    g0768(.A(new_n748), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n241), .A2(G45), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT110), .Z(new_n971));
  NOR2_X1   g0771(.A1(new_n298), .A2(G50), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT50), .ZN(new_n973));
  AOI21_X1  g0773(.A(G45), .B1(G68), .B2(G77), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n973), .A2(new_n650), .A3(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n971), .A2(new_n681), .A3(new_n975), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n976), .B1(G107), .B2(new_n209), .C1(new_n650), .C2(new_n688), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n969), .B1(new_n977), .B2(new_n695), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT111), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n967), .A2(new_n968), .A3(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT117), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n896), .A2(new_n747), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n896), .A2(new_n678), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n983), .A2(new_n745), .A3(new_n897), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n981), .A2(new_n982), .A3(new_n984), .ZN(G393));
  NAND2_X1  g0785(.A1(new_n892), .A2(new_n637), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n889), .B1(new_n636), .B2(new_n630), .C1(new_n890), .C2(new_n891), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n648), .B1(new_n988), .B2(new_n897), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n898), .A2(new_n900), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT119), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n969), .B1(new_n885), .B2(new_n693), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n729), .A2(G150), .B1(G159), .B2(new_n713), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT51), .Z(new_n996));
  NAND2_X1  g0796(.A1(new_n731), .A2(new_n767), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n708), .A2(new_n205), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n726), .A2(new_n223), .B1(new_n704), .B2(new_n298), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n721), .B2(G50), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n996), .A2(new_n997), .A3(new_n999), .A4(new_n1001), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n281), .B(new_n1002), .C1(G87), .C2(new_n724), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n281), .B1(new_n453), .B2(new_n704), .C1(new_n758), .C2(new_n573), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n729), .A2(G317), .B1(G311), .B2(new_n713), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT52), .Z(new_n1006));
  NAND2_X1  g0806(.A1(new_n731), .A2(G322), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G283), .A2(new_n733), .B1(new_n724), .B2(G107), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1004), .B(new_n1009), .C1(G116), .C2(new_n709), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n694), .B1(new_n1003), .B2(new_n1010), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n695), .B1(new_n215), .B2(new_n209), .C1(new_n253), .C2(new_n682), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n994), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n989), .A2(KEYINPUT119), .A3(new_n990), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT118), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n988), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n986), .A2(new_n987), .A3(KEYINPUT118), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1016), .A2(new_n747), .A3(new_n1017), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n993), .A2(new_n1013), .A3(new_n1014), .A4(new_n1018), .ZN(G390));
  NOR2_X1   g0819(.A1(new_n658), .A2(new_n783), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1020), .A2(new_n784), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n800), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n828), .B(new_n861), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n862), .A2(new_n863), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n860), .B1(new_n857), .B2(new_n800), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n806), .A2(new_n662), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n800), .A2(new_n677), .A3(new_n785), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1023), .B(new_n1029), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n747), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n862), .A2(new_n691), .A3(new_n863), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n779), .A2(new_n298), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n999), .B1(new_n213), .B2(new_n726), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n274), .B(new_n1036), .C1(G283), .C2(new_n729), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n772), .B1(new_n226), .B2(new_n712), .C1(new_n453), .C2(new_n699), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G97), .B2(new_n705), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1037), .B(new_n1039), .C1(new_n355), .C2(new_n758), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n947), .A2(new_n726), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT53), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  XOR2_X1   g0843(.A(KEYINPUT54), .B(G143), .Z(new_n1044));
  AOI22_X1  g0844(.A1(new_n721), .A2(G137), .B1(new_n705), .B2(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n729), .A2(G128), .B1(G132), .B2(new_n713), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G50), .A2(new_n724), .B1(new_n731), .B2(G125), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n281), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n709), .A2(G159), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1045), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1040), .B1(new_n1043), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n694), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1034), .A2(new_n748), .A3(new_n1035), .A4(new_n1053), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n851), .A2(new_n869), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n835), .A2(G330), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1029), .B(new_n1021), .C1(new_n1056), .C2(new_n800), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n800), .B1(new_n677), .B2(new_n785), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n857), .B1(new_n1027), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1055), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n1031), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1055), .A2(new_n1028), .A3(new_n1030), .A4(new_n1060), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n745), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1033), .B(new_n1054), .C1(new_n1063), .C2(new_n1065), .ZN(G378));
  NAND2_X1  g0866(.A1(new_n854), .A2(new_n847), .ZN(new_n1067));
  XOR2_X1   g0867(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n315), .A2(KEYINPUT55), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n315), .A2(KEYINPUT55), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n305), .A2(new_n810), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n1071), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n315), .A2(KEYINPUT55), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1073), .B1(new_n1076), .B2(new_n1070), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1069), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1074), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1076), .A2(new_n1073), .A3(new_n1070), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1079), .A2(new_n1068), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  AND4_X1   g0882(.A1(G330), .A2(new_n1067), .A3(new_n831), .A4(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1082), .B1(new_n855), .B2(G330), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n866), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1064), .A2(new_n1055), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1082), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n849), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n855), .A2(G330), .A3(new_n1082), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1088), .A2(new_n865), .A3(new_n1089), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1085), .A2(new_n1086), .A3(KEYINPUT57), .A4(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n745), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1086), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT123), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n1088), .A2(new_n865), .A3(new_n1089), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n865), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1095), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1085), .A2(KEYINPUT123), .A3(new_n1090), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1094), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1093), .B1(new_n1100), .B2(KEYINPUT57), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1082), .A2(new_n691), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n721), .A2(G97), .B1(G68), .B2(new_n709), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n226), .B2(new_n741), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n723), .A2(new_n247), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n1104), .A2(new_n274), .A3(new_n1105), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n458), .B1(new_n699), .B2(new_n736), .C1(new_n205), .C2(new_n726), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n363), .B2(new_n705), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1106), .B(new_n1108), .C1(new_n355), .C2(new_n712), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT58), .Z(new_n1110));
  OAI21_X1  g0910(.A(new_n202), .B1(new_n279), .B2(G41), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n721), .A2(G132), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n729), .A2(G125), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n733), .A2(new_n1044), .B1(new_n709), .B2(G150), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G128), .A2(new_n713), .B1(new_n705), .B2(G137), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1116), .B(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(G41), .B1(new_n731), .B2(G124), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1119), .B(new_n320), .C1(new_n700), .C2(new_n723), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT121), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1111), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n694), .B1(new_n1110), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n779), .A2(new_n202), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1102), .A2(new_n748), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1126), .B1(new_n1127), .B2(new_n747), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1101), .A2(new_n1128), .ZN(G375));
  INV_X1    g0929(.A(new_n1060), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n851), .A2(new_n869), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1132), .A2(new_n902), .A3(new_n1061), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n969), .B1(new_n1022), .B2(new_n690), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n721), .A2(new_n1044), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n700), .B2(new_n726), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G137), .B2(new_n713), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n729), .A2(G132), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT124), .Z(new_n1139));
  NAND2_X1  g0939(.A1(new_n709), .A2(G50), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n731), .A2(G128), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n704), .A2(new_n300), .ZN(new_n1143));
  NOR4_X1   g0943(.A1(new_n1142), .A2(new_n281), .A3(new_n1105), .A4(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n274), .B1(new_n733), .B2(G97), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1145), .B(new_n925), .C1(new_n355), .C2(new_n704), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G303), .A2(new_n731), .B1(new_n709), .B2(new_n363), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1147), .B1(new_n736), .B2(new_n712), .C1(new_n741), .C2(new_n453), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1146), .B(new_n1148), .C1(G116), .C2(new_n721), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n694), .B1(new_n1144), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1134), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n223), .B2(new_n779), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n1060), .B2(new_n747), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1133), .A2(new_n1153), .ZN(G381));
  AND3_X1   g0954(.A1(new_n993), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1155), .A2(new_n919), .A3(new_n943), .A4(new_n1018), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1156), .A2(G396), .A3(G393), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(G375), .A2(G378), .ZN(new_n1158));
  INV_X1    g0958(.A(G381), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1157), .A2(new_n1158), .A3(new_n792), .A4(new_n1159), .ZN(G407));
  INV_X1    g0960(.A(G213), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n1158), .B2(new_n622), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(G407), .A2(new_n1162), .ZN(G409));
  INV_X1    g0963(.A(KEYINPUT126), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n1085), .A2(KEYINPUT123), .A3(new_n1090), .ZN(new_n1165));
  AOI21_X1  g0965(.A(KEYINPUT123), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1086), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT57), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1092), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n747), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n1125), .ZN(new_n1171));
  OAI21_X1  g0971(.A(G378), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT60), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1132), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1130), .A2(KEYINPUT60), .A3(new_n1131), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1174), .A2(new_n745), .A3(new_n1061), .A4(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n1153), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n792), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(G384), .A3(new_n1153), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1161), .A2(G343), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n902), .B(new_n1086), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1184));
  INV_X1    g0984(.A(G378), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1085), .A2(new_n747), .A3(new_n1090), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1125), .A4(new_n1186), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1172), .A2(new_n1181), .A3(new_n1183), .A4(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT62), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1182), .B1(G375), .B2(G378), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT62), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1190), .A2(new_n1191), .A3(new_n1181), .A4(new_n1187), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT61), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1185), .B1(new_n1101), .B2(new_n1128), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1187), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1195), .A2(new_n1196), .A3(new_n1182), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1182), .A2(G2897), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT125), .Z(new_n1199));
  XNOR2_X1  g0999(.A(new_n1180), .B(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1194), .B1(new_n1197), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1164), .B1(new_n1193), .B2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(G393), .B(new_n755), .ZN(new_n1204));
  AND2_X1   g1004(.A1(G387), .A2(G390), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(G387), .A2(G390), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1204), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(G387), .A2(G390), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1156), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1207), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1172), .A2(new_n1183), .A3(new_n1187), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT61), .B1(new_n1212), .B2(new_n1200), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1213), .A2(new_n1189), .A3(KEYINPUT126), .A4(new_n1192), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1203), .A2(new_n1211), .A3(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(KEYINPUT63), .B1(new_n1197), .B2(new_n1201), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT61), .B1(new_n1216), .B2(new_n1188), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1197), .A2(KEYINPUT63), .A3(new_n1181), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1217), .A2(new_n1218), .A3(new_n1207), .A4(new_n1210), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1215), .A2(new_n1219), .ZN(G405));
  OR2_X1    g1020(.A1(new_n1181), .A2(KEYINPUT127), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1181), .A2(KEYINPUT127), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1205), .A2(new_n1206), .A3(new_n1204), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1208), .B1(new_n1156), .B2(new_n1209), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1221), .B(new_n1222), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(new_n1207), .A3(new_n1210), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1158), .A2(new_n1195), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1228), .B(new_n1229), .Z(G402));
endmodule


