//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n451, new_n452, new_n454, new_n455,
    new_n456, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n586, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G234));
  INV_X1    g025(.A(G2106), .ZN(new_n451));
  NOR2_X1   g026(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR4_X1   g030(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  OAI22_X1  g033(.A1(new_n455), .A2(new_n451), .B1(new_n448), .B2(new_n456), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT68), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(G101), .A3(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n462), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n472), .A2(new_n465), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n474), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n473), .A2(new_n470), .A3(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n469), .B(new_n471), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NAND4_X1  g054(.A1(new_n475), .A2(new_n472), .A3(G2105), .A4(new_n465), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n470), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n476), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(G136), .B2(new_n486), .ZN(new_n487));
  XOR2_X1   g062(.A(new_n487), .B(KEYINPUT70), .Z(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n490), .A2(new_n463), .A3(new_n465), .A4(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n475), .A2(new_n472), .A3(new_n490), .A4(new_n465), .ZN(new_n493));
  AND3_X1   g068(.A1(new_n493), .A2(KEYINPUT72), .A3(KEYINPUT4), .ZN(new_n494));
  AOI21_X1  g069(.A(KEYINPUT72), .B1(new_n493), .B2(KEYINPUT4), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(G2104), .C1(G114), .C2(new_n470), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n480), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT71), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n498), .B(new_n502), .C1(new_n480), .C2(new_n499), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n496), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(KEYINPUT73), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT5), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n514), .A2(new_n520), .ZN(G166));
  AND2_X1   g096(.A1(new_n511), .A2(new_n515), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n522), .A2(G89), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(G51), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n524), .B(new_n526), .C1(new_n527), .C2(new_n518), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n523), .A2(new_n528), .ZN(G168));
  AOI22_X1  g104(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(KEYINPUT74), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(KEYINPUT74), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n531), .A2(G651), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n518), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n522), .A2(G90), .B1(new_n534), .B2(G52), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT75), .ZN(G171));
  AOI22_X1  g112(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(new_n513), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n522), .A2(G81), .B1(new_n534), .B2(G43), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XOR2_X1   g116(.A(new_n541), .B(KEYINPUT76), .Z(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  INV_X1    g122(.A(G53), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT77), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n548), .B1(new_n549), .B2(KEYINPUT9), .ZN(new_n550));
  OAI211_X1 g125(.A(new_n534), .B(new_n550), .C1(new_n549), .C2(KEYINPUT9), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n522), .A2(G91), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n553));
  OAI211_X1 g128(.A(KEYINPUT77), .B(new_n553), .C1(new_n518), .C2(new_n548), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n513), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  INV_X1    g135(.A(G168), .ZN(G286));
  INV_X1    g136(.A(G166), .ZN(G303));
  OAI21_X1  g137(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT78), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n522), .A2(G87), .B1(new_n534), .B2(G49), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(G288));
  AOI22_X1  g141(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n567), .A2(new_n513), .ZN(new_n568));
  INV_X1    g143(.A(G86), .ZN(new_n569));
  INV_X1    g144(.A(G48), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n516), .A2(new_n569), .B1(new_n518), .B2(new_n570), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n568), .A2(new_n571), .ZN(G305));
  AOI22_X1  g147(.A1(new_n522), .A2(G85), .B1(new_n534), .B2(G47), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n513), .B2(new_n574), .ZN(G290));
  NAND2_X1  g150(.A1(new_n522), .A2(G92), .ZN(new_n576));
  XOR2_X1   g151(.A(new_n576), .B(KEYINPUT10), .Z(new_n577));
  NAND2_X1  g152(.A1(new_n511), .A2(G66), .ZN(new_n578));
  INV_X1    g153(.A(G79), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n579), .B2(new_n507), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(G54), .B2(new_n534), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(G868), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g159(.A(new_n583), .B1(G171), .B2(G868), .ZN(G321));
  NAND2_X1  g160(.A1(G286), .A2(G868), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n586), .B1(G868), .B2(new_n558), .ZN(G297));
  OAI21_X1  g162(.A(new_n586), .B1(G868), .B2(new_n558), .ZN(G280));
  AND2_X1   g163(.A1(new_n577), .A2(new_n581), .ZN(new_n589));
  INV_X1    g164(.A(G559), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n590), .B2(G860), .ZN(G148));
  NOR2_X1   g166(.A1(new_n582), .A2(G559), .ZN(new_n592));
  INV_X1    g167(.A(G868), .ZN(new_n593));
  NOR3_X1   g168(.A1(new_n592), .A2(KEYINPUT79), .A3(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n595));
  INV_X1    g170(.A(new_n592), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(new_n597));
  INV_X1    g172(.A(new_n542), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(new_n593), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n594), .B1(new_n597), .B2(new_n599), .ZN(G323));
  XOR2_X1   g175(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n601));
  XNOR2_X1  g176(.A(G323), .B(new_n601), .ZN(G282));
  NAND2_X1  g177(.A1(new_n481), .A2(G123), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n470), .A2(G111), .ZN(new_n604));
  OAI21_X1  g179(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(G135), .B2(new_n486), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT81), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(G2096), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(G2096), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n470), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2100), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n609), .A2(new_n610), .A3(new_n614), .ZN(G156));
  INV_X1    g190(.A(KEYINPUT14), .ZN(new_n616));
  XNOR2_X1  g191(.A(G2427), .B(G2438), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2430), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT15), .B(G2435), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n619), .B2(new_n618), .ZN(new_n621));
  XNOR2_X1  g196(.A(G2451), .B(G2454), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT16), .ZN(new_n623));
  XOR2_X1   g198(.A(G1341), .B(G1348), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n621), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2443), .B(G2446), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n626), .A2(new_n629), .A3(new_n627), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n631), .A2(new_n632), .A3(G14), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT82), .ZN(G401));
  XNOR2_X1  g209(.A(G2067), .B(G2678), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT84), .Z(new_n636));
  XOR2_X1   g211(.A(G2084), .B(G2090), .Z(new_n637));
  OAI21_X1  g212(.A(KEYINPUT17), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2072), .B(G2078), .Z(new_n639));
  AOI22_X1  g214(.A1(new_n638), .A2(new_n639), .B1(new_n637), .B2(new_n636), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n639), .B2(new_n638), .ZN(new_n641));
  INV_X1    g216(.A(new_n639), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n642), .A2(new_n637), .A3(new_n635), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT83), .B(KEYINPUT18), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2096), .B(G2100), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(G227));
  XOR2_X1   g223(.A(KEYINPUT85), .B(KEYINPUT19), .Z(new_n649));
  XNOR2_X1  g224(.A(G1971), .B(G1976), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1956), .B(G2474), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1961), .B(G1966), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT20), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(new_n653), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n654), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n656), .B(new_n659), .C1(new_n651), .C2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1991), .B(G1996), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1981), .B(G1986), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT86), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n663), .B(new_n667), .Z(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(G229));
  INV_X1    g244(.A(KEYINPUT99), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n486), .A2(G141), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT94), .Z(new_n672));
  INV_X1    g247(.A(G105), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n673), .A2(new_n464), .A3(G2105), .ZN(new_n674));
  NAND3_X1  g249(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT26), .ZN(new_n676));
  AOI211_X1 g251(.A(new_n674), .B(new_n676), .C1(new_n481), .C2(G129), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(KEYINPUT95), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT95), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n672), .A2(new_n680), .A3(new_n677), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G29), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(G29), .B2(G32), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT27), .B(G1996), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT96), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n685), .A2(new_n686), .ZN(new_n689));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G26), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT28), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n481), .A2(G128), .ZN(new_n693));
  INV_X1    g268(.A(G140), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n470), .A2(G116), .ZN(new_n695));
  OAI21_X1  g270(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n696));
  OAI221_X1 g271(.A(new_n693), .B1(new_n476), .B2(new_n694), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT91), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n692), .B1(new_n698), .B2(G29), .ZN(new_n699));
  INV_X1    g274(.A(G2067), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G19), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n542), .B2(new_n702), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(G1341), .ZN(new_n705));
  INV_X1    g280(.A(G34), .ZN(new_n706));
  AOI21_X1  g281(.A(G29), .B1(new_n706), .B2(KEYINPUT24), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(KEYINPUT24), .B2(new_n706), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n478), .B2(new_n690), .ZN(new_n709));
  INV_X1    g284(.A(G2084), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT30), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n713), .A2(G28), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n690), .B1(new_n713), .B2(G28), .ZN(new_n715));
  AND2_X1   g290(.A1(KEYINPUT31), .A2(G11), .ZN(new_n716));
  NOR2_X1   g291(.A1(KEYINPUT31), .A2(G11), .ZN(new_n717));
  OAI22_X1  g292(.A1(new_n714), .A2(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR3_X1   g293(.A1(new_n711), .A2(new_n712), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n704), .A2(G1341), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT98), .B(KEYINPUT23), .Z(new_n721));
  NAND2_X1  g296(.A1(new_n702), .A2(G20), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(new_n558), .B2(new_n702), .ZN(new_n724));
  INV_X1    g299(.A(G1956), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n705), .A2(new_n719), .A3(new_n720), .A4(new_n726), .ZN(new_n727));
  NOR3_X1   g302(.A1(new_n689), .A2(new_n701), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G29), .A2(G35), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G162), .B2(G29), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT29), .ZN(new_n731));
  INV_X1    g306(.A(G2090), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n688), .A2(new_n728), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n702), .A2(G4), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n589), .B2(new_n702), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT90), .ZN(new_n737));
  INV_X1    g312(.A(G1348), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(G168), .A2(G16), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT97), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n740), .B(new_n741), .C1(G16), .C2(G21), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n741), .B2(new_n740), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n743), .A2(G1966), .ZN(new_n744));
  OAI22_X1  g319(.A1(new_n743), .A2(G1966), .B1(new_n608), .B2(new_n690), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n739), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(G5), .A2(G16), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G171), .B2(G16), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(G1961), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n690), .A2(G33), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT25), .Z(new_n752));
  INV_X1    g327(.A(G139), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n476), .B2(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT92), .Z(new_n755));
  NAND2_X1  g330(.A1(G115), .A2(G2104), .ZN(new_n756));
  INV_X1    g331(.A(G127), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n466), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n470), .B1(new_n758), .B2(KEYINPUT93), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(KEYINPUT93), .B2(new_n758), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n750), .B1(new_n762), .B2(new_n690), .ZN(new_n763));
  INV_X1    g338(.A(G2078), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n690), .A2(G27), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G164), .B2(new_n690), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  OAI22_X1  g342(.A1(new_n763), .A2(G2072), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n764), .B2(new_n767), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n737), .A2(new_n738), .B1(new_n763), .B2(G2072), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n746), .A2(new_n749), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n670), .B1(new_n734), .B2(new_n771), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n728), .A2(new_n733), .ZN(new_n773));
  INV_X1    g348(.A(new_n771), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n773), .A2(KEYINPUT99), .A3(new_n774), .A4(new_n688), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  MUX2_X1   g351(.A(G6), .B(G305), .S(G16), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT32), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1981), .ZN(new_n779));
  NOR2_X1   g354(.A1(G16), .A2(G23), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT87), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G288), .B2(new_n702), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT33), .B(G1976), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n702), .A2(G22), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G166), .B2(new_n702), .ZN(new_n786));
  INV_X1    g361(.A(G1971), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n782), .A2(new_n783), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n784), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  OR3_X1    g365(.A1(new_n779), .A2(KEYINPUT34), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(KEYINPUT34), .B1(new_n779), .B2(new_n790), .ZN(new_n792));
  MUX2_X1   g367(.A(G24), .B(G290), .S(G16), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1986), .ZN(new_n794));
  NOR2_X1   g369(.A1(G25), .A2(G29), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n486), .A2(G131), .ZN(new_n796));
  INV_X1    g371(.A(G119), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n470), .A2(G107), .ZN(new_n798));
  OAI21_X1  g373(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n799));
  OAI22_X1  g374(.A1(new_n480), .A2(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n795), .B1(new_n801), .B2(G29), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT35), .B(G1991), .Z(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n802), .A2(new_n804), .ZN(new_n806));
  NOR3_X1   g381(.A1(new_n794), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n791), .A2(new_n792), .A3(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(KEYINPUT88), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(KEYINPUT88), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n809), .A2(KEYINPUT36), .A3(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n808), .A2(KEYINPUT36), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n811), .A2(KEYINPUT89), .A3(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT89), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n809), .A2(new_n814), .A3(KEYINPUT36), .A4(new_n810), .ZN(new_n815));
  AND3_X1   g390(.A1(new_n776), .A2(new_n813), .A3(new_n815), .ZN(G311));
  NAND3_X1  g391(.A1(new_n776), .A2(new_n813), .A3(new_n815), .ZN(G150));
  AOI22_X1  g392(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(new_n513), .ZN(new_n819));
  INV_X1    g394(.A(G93), .ZN(new_n820));
  INV_X1    g395(.A(G55), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n516), .A2(new_n820), .B1(new_n518), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n823), .A2(new_n539), .A3(new_n540), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n542), .B2(new_n823), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT38), .Z(new_n826));
  NAND2_X1  g401(.A1(new_n589), .A2(G559), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n829));
  INV_X1    g404(.A(G860), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n823), .A2(new_n830), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT37), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(G145));
  XNOR2_X1  g410(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n478), .B(KEYINPUT100), .ZN(new_n838));
  XNOR2_X1  g413(.A(G162), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n608), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n481), .A2(G130), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n470), .A2(G118), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(G142), .B2(new_n486), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n612), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n801), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT101), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n500), .B1(new_n496), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g424(.A(KEYINPUT101), .B(new_n492), .C1(new_n494), .C2(new_n495), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n698), .B(new_n851), .Z(new_n852));
  INV_X1    g427(.A(KEYINPUT102), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n682), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n679), .A2(KEYINPUT102), .A3(new_n681), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n761), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n678), .A2(new_n761), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n852), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n855), .ZN(new_n860));
  AOI21_X1  g435(.A(KEYINPUT102), .B1(new_n679), .B2(new_n681), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n762), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n852), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n863), .A3(new_n857), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n847), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n859), .A2(new_n864), .A3(new_n847), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n840), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n865), .A2(new_n866), .ZN(new_n872));
  AOI211_X1 g447(.A(KEYINPUT103), .B(new_n847), .C1(new_n859), .C2(new_n864), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n840), .B(new_n868), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(G37), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n837), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n840), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n872), .A2(new_n873), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n868), .B(KEYINPUT104), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n881), .A2(new_n875), .A3(new_n874), .A4(new_n836), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n877), .A2(new_n882), .ZN(G395));
  XNOR2_X1  g458(.A(G288), .B(G305), .ZN(new_n884));
  XNOR2_X1  g459(.A(G290), .B(G166), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT108), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n887), .B1(new_n888), .B2(KEYINPUT42), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n589), .A2(G299), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n582), .A2(new_n558), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(KEYINPUT106), .A3(new_n892), .ZN(new_n893));
  OR3_X1    g468(.A1(new_n582), .A2(KEYINPUT106), .A3(new_n558), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT107), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n825), .B(new_n596), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n888), .A2(KEYINPUT42), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n898), .ZN(new_n902));
  INV_X1    g477(.A(new_n895), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT41), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n891), .A2(new_n892), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n902), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n899), .A2(new_n901), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n901), .B1(new_n899), .B2(new_n908), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n890), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n899), .A2(new_n908), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n900), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n899), .A2(new_n901), .A3(new_n908), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n914), .A3(new_n889), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(G868), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n823), .A2(G868), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(G295));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n917), .A2(new_n921), .A3(new_n919), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n593), .B1(new_n911), .B2(new_n915), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT109), .B1(new_n923), .B2(new_n918), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(G331));
  XNOR2_X1  g500(.A(G171), .B(G168), .ZN(new_n926));
  INV_X1    g501(.A(new_n825), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n926), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n904), .A2(new_n907), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n926), .A2(new_n825), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n926), .A2(new_n825), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n903), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n887), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n933), .B(new_n887), .C1(new_n928), .C2(new_n929), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n875), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT43), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n895), .B(KEYINPUT107), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n887), .B1(new_n928), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n905), .A2(KEYINPUT41), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n940), .B(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(KEYINPUT41), .B2(new_n895), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n939), .B1(new_n943), .B2(new_n928), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n944), .A2(new_n945), .A3(new_n875), .A4(new_n935), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n937), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n945), .B1(new_n934), .B2(new_n936), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n944), .A2(KEYINPUT43), .A3(new_n875), .A4(new_n935), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  MUX2_X1   g525(.A(new_n947), .B(new_n950), .S(KEYINPUT44), .Z(G397));
  INV_X1    g526(.A(G1384), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n851), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n954));
  INV_X1    g529(.A(G40), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n478), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT111), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT111), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n953), .A2(new_n959), .A3(new_n954), .A4(new_n956), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT112), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n958), .A2(KEYINPUT112), .A3(new_n960), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n698), .A2(G2067), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n698), .A2(G2067), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n678), .A2(G1996), .ZN(new_n968));
  AOI22_X1  g543(.A1(new_n963), .A2(new_n964), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n801), .A2(new_n803), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n796), .A2(new_n800), .A3(new_n804), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n972), .B1(new_n963), .B2(new_n964), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n961), .A2(new_n682), .A3(G1996), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n969), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(G290), .B(G1986), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n958), .A2(new_n960), .A3(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n481), .A2(G126), .ZN(new_n980));
  INV_X1    g555(.A(new_n492), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT72), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n493), .A2(KEYINPUT72), .A3(KEYINPUT4), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n981), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n980), .B(new_n498), .C1(new_n986), .C2(KEYINPUT101), .ZN(new_n987));
  INV_X1    g562(.A(new_n850), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n979), .B(new_n952), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT114), .ZN(new_n990));
  AOI211_X1 g565(.A(new_n990), .B(new_n979), .C1(new_n504), .C2(new_n952), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n501), .A2(new_n503), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n952), .B1(new_n986), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT114), .B1(new_n993), .B2(KEYINPUT50), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n956), .B(new_n989), .C1(new_n991), .C2(new_n994), .ZN(new_n995));
  XOR2_X1   g570(.A(KEYINPUT121), .B(G1961), .Z(new_n996));
  INV_X1    g571(.A(new_n956), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(new_n953), .B2(new_n954), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(G2078), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(G1384), .B1(new_n849), .B2(new_n850), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1001), .B1(new_n1002), .B2(KEYINPUT45), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n995), .A2(new_n996), .B1(new_n998), .B2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(KEYINPUT45), .B(new_n952), .C1(new_n987), .C2(new_n988), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n1006));
  AOI211_X1 g581(.A(new_n1006), .B(KEYINPUT45), .C1(new_n504), .C2(new_n952), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT113), .B1(new_n993), .B2(new_n954), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n956), .B(new_n1005), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n999), .B1(new_n1009), .B2(G2078), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1004), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(G171), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n995), .A2(new_n996), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n952), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n998), .A2(new_n1000), .A3(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1010), .A2(G301), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1012), .A2(KEYINPUT54), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT123), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1012), .A2(KEYINPUT123), .A3(KEYINPUT54), .A4(new_n1016), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT122), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G303), .A2(G8), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT55), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G8), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1009), .A2(new_n787), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n956), .B1(new_n993), .B2(KEYINPUT50), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1028), .B1(KEYINPUT50), .B2(new_n953), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n732), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1026), .B1(new_n1031), .B2(KEYINPUT116), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n787), .A2(new_n1009), .B1(new_n1029), .B2(new_n732), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1025), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n564), .A2(G1976), .A3(new_n565), .ZN(new_n1037));
  XOR2_X1   g612(.A(new_n1037), .B(KEYINPUT115), .Z(new_n1038));
  NAND2_X1  g613(.A1(new_n1002), .A2(new_n956), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(G8), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT52), .ZN(new_n1041));
  INV_X1    g616(.A(G1976), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(G288), .B2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1038), .A2(G8), .A3(new_n1039), .A4(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(G305), .A2(G1981), .ZN(new_n1045));
  OR3_X1    g620(.A1(new_n568), .A2(new_n571), .A3(G1981), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(KEYINPUT49), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(G8), .A3(new_n1039), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1041), .A2(new_n1044), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n501), .A2(new_n503), .ZN(new_n1052));
  AOI21_X1  g627(.A(G1384), .B1(new_n1052), .B2(new_n496), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n990), .B1(new_n1053), .B2(new_n979), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n993), .A2(KEYINPUT114), .A3(KEYINPUT50), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n997), .B1(new_n1002), .B2(new_n979), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n732), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1026), .B1(new_n1027), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n1025), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1051), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1022), .B1(new_n1036), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(G8), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1031), .A2(KEYINPUT116), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1024), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1050), .B1(new_n1025), .B2(new_n1059), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(KEYINPUT122), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1010), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G171), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1004), .A2(new_n1010), .A3(G301), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT54), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1056), .A2(new_n710), .A3(new_n1057), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n956), .B(new_n1014), .C1(new_n1002), .C2(KEYINPUT45), .ZN(new_n1073));
  INV_X1    g648(.A(G1966), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G8), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1026), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1080));
  NAND2_X1  g655(.A1(G286), .A2(G8), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n1081), .B(KEYINPUT120), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT51), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  AOI211_X1 g658(.A(new_n1026), .B(G168), .C1(new_n1072), .C2(new_n1075), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1079), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1071), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1021), .A2(new_n1062), .A3(new_n1067), .A4(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1002), .A2(new_n979), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n725), .B1(new_n1088), .B2(new_n1028), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT56), .B(G2072), .Z(new_n1090));
  OAI21_X1  g665(.A(new_n1089), .B1(new_n1009), .B2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n558), .B(KEYINPUT57), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1039), .A2(G2067), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1095), .B1(new_n995), .B2(new_n738), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1094), .B1(new_n582), .B2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1089), .B(new_n1092), .C1(new_n1009), .C2(new_n1090), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1096), .A2(KEYINPUT60), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1100), .A2(KEYINPUT119), .A3(new_n582), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n582), .B1(new_n1100), .B2(KEYINPUT119), .ZN(new_n1102));
  OAI22_X1  g677(.A1(new_n1101), .A2(new_n1102), .B1(KEYINPUT119), .B2(new_n1100), .ZN(new_n1103));
  OR2_X1    g678(.A1(new_n1096), .A2(KEYINPUT60), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT58), .B(G1341), .Z(new_n1106));
  NAND2_X1  g681(.A1(new_n1039), .A2(new_n1106), .ZN(new_n1107));
  XOR2_X1   g682(.A(KEYINPUT117), .B(G1996), .Z(new_n1108));
  OAI21_X1  g683(.A(new_n1107), .B1(new_n1009), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n542), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT59), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1109), .A2(new_n1112), .A3(new_n542), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT61), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1094), .A2(new_n1115), .A3(new_n1098), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1115), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1114), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1120), .B(new_n1114), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1105), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1087), .B1(new_n1099), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1077), .A2(G286), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1065), .A2(new_n1066), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT63), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n1059), .A2(new_n1025), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1066), .A2(KEYINPUT63), .A3(new_n1128), .A4(new_n1124), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1039), .A2(G8), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1049), .A2(new_n1042), .A3(new_n564), .A4(new_n565), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1131), .B1(new_n1132), .B2(new_n1046), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1060), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1133), .B1(new_n1134), .B2(new_n1051), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1069), .B1(new_n1085), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1137), .A2(new_n1062), .A3(new_n1067), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT124), .B1(new_n1085), .B2(new_n1136), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1080), .A2(G286), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1140), .B(KEYINPUT51), .C1(new_n1080), .C2(new_n1082), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1141), .A2(new_n1142), .A3(KEYINPUT62), .A4(new_n1079), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1130), .B(new_n1135), .C1(new_n1138), .C2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n978), .B1(new_n1123), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n967), .A2(new_n968), .ZN(new_n1147));
  INV_X1    g722(.A(new_n964), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT112), .B1(new_n958), .B2(new_n960), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n974), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1150), .A2(new_n1151), .A3(new_n971), .ZN(new_n1152));
  INV_X1    g727(.A(new_n966), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n963), .A2(new_n964), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n961), .A2(G1986), .A3(G290), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT48), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1154), .A2(new_n1155), .B1(new_n975), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT47), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n965), .A2(new_n966), .A3(new_n678), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1161), .B1(new_n963), .B2(new_n964), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT125), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n961), .A2(G1996), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT46), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1164), .B(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1160), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1162), .A2(KEYINPUT125), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n1169));
  AOI211_X1 g744(.A(new_n1169), .B(new_n1161), .C1(new_n963), .C2(new_n964), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1166), .B(new_n1160), .C1(new_n1168), .C2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1159), .B1(new_n1167), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(KEYINPUT126), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n1175));
  OAI211_X1 g750(.A(new_n1159), .B(new_n1175), .C1(new_n1167), .C2(new_n1172), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1146), .A2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g753(.A(G319), .ZN(new_n1180));
  NOR3_X1   g754(.A1(G401), .A2(new_n1180), .A3(G227), .ZN(new_n1181));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n1182));
  XNOR2_X1  g756(.A(new_n1181), .B(new_n1182), .ZN(new_n1183));
  NAND2_X1  g757(.A1(new_n1183), .A2(new_n668), .ZN(new_n1184));
  AOI21_X1  g758(.A(new_n1184), .B1(new_n937), .B2(new_n946), .ZN(new_n1185));
  OAI21_X1  g759(.A(new_n1185), .B1(new_n871), .B2(new_n876), .ZN(G225));
  INV_X1    g760(.A(G225), .ZN(G308));
endmodule


