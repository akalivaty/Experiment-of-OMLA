//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT3), .B1(new_n187), .B2(G107), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G104), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n187), .A2(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G101), .ZN(new_n194));
  INV_X1    g008(.A(G101), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n188), .A2(new_n191), .A3(new_n195), .A4(new_n192), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(KEYINPUT4), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT4), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n193), .A2(new_n198), .A3(G101), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n203), .A2(KEYINPUT64), .A3(G146), .ZN(new_n204));
  AOI21_X1  g018(.A(KEYINPUT64), .B1(new_n203), .B2(G146), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n202), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(KEYINPUT65), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n203), .A2(G146), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n213), .B1(new_n201), .B2(G143), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n203), .A2(KEYINPUT64), .A3(G146), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n212), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  OR2_X1    g030(.A1(new_n207), .A2(new_n208), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n211), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n203), .A2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n202), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n207), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n210), .A2(new_n218), .A3(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n187), .A2(G107), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n190), .A2(G104), .ZN(new_n225));
  OAI21_X1  g039(.A(G101), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n196), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G128), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n230), .B1(G143), .B2(new_n201), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT76), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n229), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT76), .B1(new_n212), .B2(new_n230), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n221), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n202), .A2(new_n219), .A3(new_n230), .A4(G128), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n228), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT10), .ZN(new_n239));
  AOI22_X1  g053(.A1(new_n200), .A2(new_n223), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n229), .B1(new_n202), .B2(KEYINPUT1), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n236), .B1(new_n216), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT77), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n196), .A2(new_n226), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n243), .B1(new_n196), .B2(new_n226), .ZN(new_n245));
  OAI211_X1 g059(.A(KEYINPUT10), .B(new_n242), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT11), .ZN(new_n247));
  INV_X1    g061(.A(G134), .ZN(new_n248));
  OAI211_X1 g062(.A(KEYINPUT66), .B(new_n247), .C1(new_n248), .C2(G137), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G137), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G134), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT66), .B1(new_n252), .B2(new_n247), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT67), .B1(new_n251), .B2(G134), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n255), .B1(new_n247), .B2(new_n252), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n251), .A2(KEYINPUT67), .A3(KEYINPUT11), .A4(G134), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(G131), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT66), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n248), .A2(G137), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n260), .B1(new_n261), .B2(KEYINPUT11), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n249), .ZN(new_n263));
  INV_X1    g077(.A(G131), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n263), .A2(new_n264), .A3(new_n256), .A4(new_n257), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT78), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT78), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n259), .A2(new_n268), .A3(new_n265), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n240), .A2(new_n246), .A3(new_n267), .A4(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n202), .A2(new_n232), .A3(KEYINPUT1), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n234), .A2(G128), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n237), .B1(new_n272), .B2(new_n220), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n239), .B1(new_n273), .B2(new_n227), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n210), .A2(new_n218), .A3(new_n222), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n197), .A2(new_n199), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n274), .B(new_n246), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n266), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n270), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(G110), .B(G140), .ZN(new_n280));
  INV_X1    g094(.A(G953), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n281), .A2(G227), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n280), .B(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n283), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT80), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n286), .B1(new_n228), .B2(new_n242), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n206), .B1(new_n229), .B2(new_n231), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n288), .A2(KEYINPUT80), .A3(new_n236), .A4(new_n227), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n238), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(KEYINPUT79), .A2(KEYINPUT12), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT12), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT79), .B1(new_n259), .B2(new_n265), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n290), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n293), .B1(new_n290), .B2(new_n294), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n270), .B(new_n285), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n284), .B2(new_n297), .ZN(new_n298));
  XOR2_X1   g112(.A(KEYINPUT82), .B(G469), .Z(new_n299));
  AND2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n270), .B1(new_n295), .B2(new_n296), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT81), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT81), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n270), .B(new_n304), .C1(new_n295), .C2(new_n296), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n285), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n270), .A2(new_n285), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n307), .B1(new_n266), .B2(new_n277), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n301), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n300), .B1(new_n309), .B2(G469), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT9), .B(G234), .ZN(new_n311));
  OAI21_X1  g125(.A(G221), .B1(new_n311), .B2(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G125), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n315), .B(new_n236), .C1(new_n216), .C2(new_n241), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n317), .B1(new_n275), .B2(G125), .ZN(new_n318));
  INV_X1    g132(.A(G224), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(G953), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n318), .B(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G119), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G116), .ZN(new_n324));
  OAI21_X1  g138(.A(G113), .B1(new_n324), .B2(KEYINPUT5), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(G116), .B(G119), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT5), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT2), .B(G113), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  AOI22_X1  g144(.A1(new_n326), .A2(new_n328), .B1(new_n330), .B2(new_n327), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n244), .B2(new_n245), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n327), .ZN(new_n333));
  INV_X1    g147(.A(G116), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G119), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n324), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n329), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n197), .A2(new_n338), .A3(new_n199), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT6), .ZN(new_n341));
  XNOR2_X1  g155(.A(G110), .B(G122), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n340), .A2(new_n343), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n332), .A2(new_n339), .A3(new_n342), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(KEYINPUT6), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n322), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n328), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n333), .B1(new_n349), .B2(new_n325), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n228), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n331), .A2(new_n227), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT83), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n342), .B(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT8), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n342), .B(KEYINPUT83), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT8), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n351), .A2(new_n352), .A3(new_n356), .A4(new_n358), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n359), .A2(new_n346), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n275), .A2(G125), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n361), .A2(KEYINPUT7), .A3(new_n321), .A4(new_n316), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT84), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT84), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n318), .A2(new_n364), .A3(KEYINPUT7), .A4(new_n321), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n321), .A2(KEYINPUT7), .ZN(new_n366));
  OR2_X1    g180(.A1(new_n318), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n360), .A2(new_n363), .A3(new_n365), .A4(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n348), .A2(new_n368), .A3(new_n301), .ZN(new_n369));
  OAI21_X1  g183(.A(G210), .B1(G237), .B2(G902), .ZN(new_n370));
  XOR2_X1   g184(.A(new_n370), .B(KEYINPUT85), .Z(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(G214), .B1(G237), .B2(G902), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n348), .A2(new_n368), .A3(new_n301), .A4(new_n371), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G475), .ZN(new_n377));
  INV_X1    g191(.A(G237), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT68), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT68), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G237), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(G214), .A3(new_n281), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n203), .ZN(new_n384));
  AOI21_X1  g198(.A(G953), .B1(new_n379), .B2(new_n381), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(G143), .A3(G214), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT86), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT18), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n384), .B(new_n386), .C1(new_n264), .C2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(G125), .B(G140), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n201), .ZN(new_n391));
  INV_X1    g205(.A(G140), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n315), .B2(KEYINPUT72), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT72), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(G125), .A3(G140), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n391), .B1(new_n396), .B2(new_n201), .ZN(new_n397));
  AND4_X1   g211(.A1(G143), .A2(new_n382), .A3(G214), .A4(new_n281), .ZN(new_n398));
  AOI21_X1  g212(.A(G143), .B1(new_n385), .B2(G214), .ZN(new_n399));
  OAI21_X1  g213(.A(G131), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n389), .B(new_n397), .C1(new_n400), .C2(new_n388), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT17), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n384), .A2(new_n264), .A3(new_n386), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT16), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n392), .A3(G125), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT73), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n406), .A2(new_n392), .A3(KEYINPUT73), .A4(G125), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n406), .B1(new_n393), .B2(new_n395), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n201), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n396), .A2(KEYINPUT16), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n414), .A2(G146), .A3(new_n409), .A4(new_n410), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n413), .B(new_n415), .C1(new_n400), .C2(new_n402), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n401), .B1(new_n405), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G113), .B(G122), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(new_n187), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT89), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n419), .B(new_n401), .C1(new_n405), .C2(new_n416), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n264), .B1(new_n384), .B2(new_n386), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT17), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n404), .A2(new_n426), .A3(new_n413), .A4(new_n415), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n419), .B1(new_n427), .B2(new_n401), .ZN(new_n428));
  AOI21_X1  g242(.A(G902), .B1(new_n428), .B2(KEYINPUT89), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n377), .B1(new_n424), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(G475), .A2(G902), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n400), .A2(new_n403), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT87), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n400), .A2(KEYINPUT87), .A3(new_n403), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n411), .A2(new_n412), .A3(new_n201), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT19), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n396), .A2(new_n437), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n390), .A2(new_n437), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n436), .B1(new_n201), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n434), .A2(new_n435), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n419), .B1(new_n442), .B2(new_n401), .ZN(new_n443));
  INV_X1    g257(.A(new_n423), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n431), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT88), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n435), .A2(new_n441), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT87), .B1(new_n400), .B2(new_n403), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n401), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n420), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n446), .B1(new_n450), .B2(new_n423), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n445), .B1(new_n451), .B2(KEYINPUT20), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n423), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n453), .A2(new_n446), .A3(new_n454), .A4(new_n431), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n430), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G217), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n311), .A2(new_n457), .A3(G953), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n334), .A2(G122), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n334), .A2(G122), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n459), .B1(new_n460), .B2(KEYINPUT14), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT90), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT90), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n463), .B(new_n459), .C1(new_n460), .C2(KEYINPUT14), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n462), .B(new_n464), .C1(KEYINPUT14), .C2(new_n459), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G107), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n203), .A2(G128), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n229), .A2(G143), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G134), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n467), .A2(new_n468), .A3(new_n248), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n334), .A2(G122), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n473), .A2(new_n460), .A3(G107), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n466), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n460), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n190), .B1(new_n479), .B2(new_n459), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n471), .B1(new_n480), .B2(new_n474), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT13), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n467), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n203), .A2(KEYINPUT13), .A3(G128), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n484), .A3(new_n468), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n485), .A2(G134), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n458), .B1(new_n478), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n476), .B1(new_n465), .B2(G107), .ZN(new_n490));
  INV_X1    g304(.A(new_n458), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n490), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n301), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT91), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G478), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(KEYINPUT15), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n478), .A2(new_n488), .A3(new_n458), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n491), .B1(new_n490), .B2(new_n487), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(KEYINPUT91), .A3(new_n301), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n495), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n493), .A2(new_n497), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(G234), .A2(G237), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n505), .A2(G952), .A3(new_n281), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n505), .A2(G902), .A3(G953), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT21), .B(G898), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n376), .A2(new_n456), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n314), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT92), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n314), .A2(KEYINPUT92), .A3(new_n511), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n385), .A2(G210), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT26), .B(G101), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n338), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n275), .B1(new_n265), .B2(new_n259), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n251), .A2(G134), .ZN(new_n525));
  OAI21_X1  g339(.A(G131), .B1(new_n261), .B2(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n265), .A2(new_n242), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT30), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n266), .A2(new_n223), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n265), .A2(new_n242), .A3(new_n526), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n523), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n524), .A2(new_n338), .A3(new_n527), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n522), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n523), .B1(new_n529), .B2(new_n531), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT28), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n529), .A2(new_n523), .A3(new_n531), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT28), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n537), .A2(new_n521), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT29), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n535), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n301), .B1(new_n541), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g358(.A(G472), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n338), .B1(new_n524), .B2(new_n527), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n539), .B1(new_n546), .B2(new_n538), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n534), .A2(KEYINPUT28), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n522), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n538), .A2(new_n521), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT31), .B1(new_n533), .B2(new_n550), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n524), .A2(KEYINPUT30), .A3(new_n527), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n530), .B1(new_n529), .B2(new_n531), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n338), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT31), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n538), .A2(new_n521), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n549), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT32), .ZN(new_n559));
  NOR2_X1   g373(.A1(G472), .A2(G902), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n559), .B1(new_n558), .B2(new_n560), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n545), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT70), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT70), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n545), .B(new_n565), .C1(new_n561), .C2(new_n562), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n415), .A2(new_n413), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT71), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(G119), .B2(new_n229), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT23), .B1(new_n229), .B2(G119), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n323), .A2(G128), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT23), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT71), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n569), .A2(new_n570), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(G119), .B(G128), .ZN(new_n576));
  XOR2_X1   g390(.A(KEYINPUT24), .B(G110), .Z(new_n577));
  AOI22_X1  g391(.A1(new_n575), .A2(G110), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n567), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G110), .ZN(new_n580));
  OAI211_X1 g394(.A(G119), .B(new_n229), .C1(new_n568), .C2(KEYINPUT23), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n572), .B1(new_n323), .B2(G128), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT71), .B1(new_n323), .B2(G128), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n580), .B(new_n581), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  OAI22_X1  g398(.A1(new_n584), .A2(KEYINPUT74), .B1(new_n576), .B2(new_n577), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT74), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(new_n574), .B2(new_n580), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n415), .B(new_n391), .C1(new_n585), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n579), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT22), .B(G137), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n281), .A2(G221), .A3(G234), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n579), .A2(new_n588), .A3(new_n592), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n457), .B1(G234), .B2(new_n301), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(G902), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(new_n599), .B(KEYINPUT75), .Z(new_n600));
  NAND3_X1  g414(.A1(new_n594), .A2(new_n301), .A3(new_n595), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT25), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT25), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n594), .A2(new_n603), .A3(new_n301), .A4(new_n595), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(new_n604), .A3(new_n597), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n564), .A2(new_n566), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n516), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G101), .ZN(G3));
  INV_X1    g424(.A(G472), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n558), .B2(new_n301), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n558), .A2(new_n560), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR4_X1   g429(.A1(new_n615), .A2(new_n310), .A3(new_n606), .A4(new_n313), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n301), .A2(G478), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n498), .A2(KEYINPUT93), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n500), .A2(new_n618), .A3(KEYINPUT33), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n498), .B(new_n499), .C1(KEYINPUT93), .C2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n617), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n495), .A2(new_n501), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n622), .B1(new_n623), .B2(new_n496), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n456), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n509), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n373), .A2(new_n626), .A3(new_n374), .A4(new_n375), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n616), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT94), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT34), .B(G104), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  NAND2_X1  g446(.A1(new_n424), .A2(new_n429), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(G475), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT95), .B(KEYINPUT20), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n445), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n453), .A2(new_n431), .A3(new_n635), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n634), .A2(new_n504), .A3(new_n637), .A4(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n627), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n616), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  NOR2_X1   g457(.A1(new_n593), .A2(KEYINPUT36), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n589), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n598), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n605), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT96), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n605), .A2(KEYINPUT96), .A3(new_n646), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n615), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n516), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT37), .B(G110), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  NAND2_X1  g471(.A1(new_n614), .A2(KEYINPUT32), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n565), .B1(new_n660), .B2(new_n545), .ZN(new_n661));
  INV_X1    g475(.A(new_n566), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n651), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n506), .B(KEYINPUT99), .Z(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(G900), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n666), .B1(new_n667), .B2(new_n507), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n639), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n376), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n310), .A2(new_n670), .A3(new_n313), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n663), .A2(new_n664), .A3(new_n669), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  XOR2_X1   g487(.A(new_n668), .B(KEYINPUT39), .Z(new_n674));
  NAND2_X1  g488(.A1(new_n314), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n676));
  INV_X1    g490(.A(new_n504), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n533), .A2(new_n534), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n522), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n546), .A2(new_n538), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n301), .B1(new_n680), .B2(new_n521), .ZN(new_n681));
  OAI21_X1  g495(.A(G472), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  AOI211_X1 g496(.A(new_n456), .B(new_n677), .C1(new_n660), .C2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n373), .A2(new_n375), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT38), .ZN(new_n685));
  INV_X1    g499(.A(new_n374), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n685), .A2(new_n686), .A3(new_n647), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n676), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT100), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT100), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n676), .A2(new_n688), .A3(new_n692), .A4(new_n689), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n203), .ZN(G45));
  NOR3_X1   g509(.A1(new_n456), .A2(new_n624), .A3(new_n668), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n663), .A2(new_n664), .A3(new_n671), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G146), .ZN(G48));
  NAND2_X1  g512(.A1(new_n298), .A2(new_n299), .ZN(new_n699));
  INV_X1    g513(.A(G469), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n699), .B(new_n312), .C1(new_n298), .C2(new_n700), .ZN(new_n701));
  NOR4_X1   g515(.A1(new_n701), .A2(new_n456), .A3(new_n627), .A4(new_n624), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n702), .A2(new_n564), .A3(new_n566), .A4(new_n607), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT41), .B(G113), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  NOR3_X1   g519(.A1(new_n701), .A2(new_n639), .A3(new_n627), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n564), .A2(new_n706), .A3(new_n566), .A4(new_n607), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G116), .ZN(G18));
  OR2_X1    g522(.A1(new_n298), .A2(new_n700), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n376), .A2(new_n312), .A3(new_n709), .A4(new_n699), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n456), .A2(new_n510), .A3(new_n649), .A4(new_n650), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n564), .A3(new_n566), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT101), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n712), .A2(new_n564), .A3(KEYINPUT101), .A4(new_n566), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  NOR3_X1   g532(.A1(new_n701), .A2(new_n456), .A3(new_n677), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n521), .B1(new_n537), .B2(new_n540), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n555), .B1(new_n554), .B2(new_n556), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT103), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT103), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n549), .A2(new_n551), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n722), .A2(new_n557), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n560), .B(KEYINPUT102), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n612), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n719), .A2(new_n727), .A3(new_n607), .A4(new_n628), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  NAND3_X1  g543(.A1(new_n727), .A2(new_n696), .A3(new_n647), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n710), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n315), .ZN(G27));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n684), .A2(new_n374), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n310), .A2(new_n313), .A3(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n735), .A2(new_n564), .A3(new_n566), .A4(new_n607), .ZN(new_n736));
  INV_X1    g550(.A(new_n696), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n733), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n733), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n606), .B1(new_n660), .B2(new_n545), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n735), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G131), .ZN(G33));
  NAND3_X1  g557(.A1(new_n608), .A2(new_n669), .A3(new_n735), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G134), .ZN(G36));
  INV_X1    g559(.A(new_n624), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n456), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n615), .A3(new_n647), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n734), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n752), .B1(new_n751), .B2(new_n750), .ZN(new_n753));
  INV_X1    g567(.A(new_n305), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n290), .A2(new_n294), .ZN(new_n755));
  INV_X1    g569(.A(new_n293), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n290), .A2(new_n293), .A3(new_n294), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n304), .B1(new_n759), .B2(new_n270), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n283), .B1(new_n754), .B2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n308), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(KEYINPUT45), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n764), .B1(new_n306), .B2(new_n308), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n765), .A3(G469), .ZN(new_n766));
  NAND2_X1  g580(.A1(G469), .A2(G902), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT46), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n300), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n766), .A2(KEYINPUT46), .A3(new_n767), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n312), .A3(new_n674), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n772), .A2(KEYINPUT104), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(KEYINPUT104), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n753), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n251), .ZN(G39));
  NOR4_X1   g590(.A1(new_n663), .A2(new_n607), .A3(new_n737), .A4(new_n734), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n771), .A2(KEYINPUT47), .A3(new_n312), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT47), .B1(new_n771), .B2(new_n312), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT105), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G140), .ZN(G42));
  NOR4_X1   g596(.A1(new_n747), .A2(new_n606), .A3(new_n313), .A4(new_n686), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT106), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n660), .A2(new_n682), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n709), .A2(new_n699), .ZN(new_n786));
  XOR2_X1   g600(.A(new_n786), .B(KEYINPUT49), .Z(new_n787));
  NAND4_X1  g601(.A1(new_n784), .A2(new_n785), .A3(new_n685), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT107), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n701), .A2(new_n734), .ZN(new_n790));
  AND4_X1   g604(.A1(new_n607), .A2(new_n785), .A3(new_n506), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n625), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(G952), .A3(new_n281), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n749), .A2(new_n666), .A3(new_n790), .ZN(new_n794));
  INV_X1    g608(.A(new_n740), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT48), .ZN(new_n797));
  INV_X1    g611(.A(new_n710), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n727), .A2(new_n607), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n749), .A2(new_n799), .A3(new_n666), .ZN(new_n800));
  AOI211_X1 g614(.A(new_n793), .B(new_n797), .C1(new_n798), .C2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n734), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n778), .A2(new_n779), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n786), .A2(new_n312), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT112), .Z(new_n806));
  OAI21_X1  g620(.A(new_n803), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n701), .A2(new_n374), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n685), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n800), .A2(KEYINPUT50), .A3(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n749), .A2(new_n809), .A3(new_n799), .A4(new_n666), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n814), .B1(KEYINPUT113), .B2(KEYINPUT51), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n814), .A2(KEYINPUT113), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n456), .A2(new_n624), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n791), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n727), .A2(new_n647), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n794), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n791), .A2(KEYINPUT114), .A3(new_n817), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n820), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n816), .A2(new_n824), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n807), .A2(new_n815), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n824), .B1(new_n813), .B2(new_n810), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n801), .B1(new_n826), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT115), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g647(.A(KEYINPUT115), .B(new_n801), .C1(new_n826), .C2(new_n830), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n564), .A2(new_n566), .A3(new_n607), .ZN(new_n836));
  INV_X1    g650(.A(new_n735), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n634), .A2(new_n637), .A3(new_n638), .ZN(new_n839));
  NOR4_X1   g653(.A1(new_n651), .A2(new_n839), .A3(new_n504), .A4(new_n668), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n564), .A2(new_n840), .A3(new_n566), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n730), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n838), .A2(new_n669), .B1(new_n842), .B2(new_n735), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n742), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n514), .B(new_n515), .C1(new_n608), .C2(new_n652), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n703), .A2(new_n707), .A3(new_n728), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n456), .A2(new_n504), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(KEYINPUT108), .A3(new_n628), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n625), .A2(new_n628), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT108), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n851), .B1(new_n847), .B2(new_n627), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n849), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n616), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n845), .A2(new_n846), .A3(new_n717), .A4(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n844), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n731), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n647), .A2(new_n668), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n683), .A2(new_n671), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n672), .A2(new_n697), .A3(new_n858), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT52), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n564), .A2(new_n566), .A3(new_n664), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n314), .A2(new_n376), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n731), .B1(new_n865), .B2(new_n669), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n866), .A2(new_n867), .A3(new_n697), .A4(new_n860), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n862), .A2(KEYINPUT110), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT110), .B1(new_n862), .B2(new_n868), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n857), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n862), .A2(new_n868), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n717), .A2(new_n845), .A3(new_n846), .A4(new_n854), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n739), .A2(new_n735), .A3(new_n740), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n663), .A2(new_n607), .A3(new_n696), .A4(new_n735), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n875), .B1(new_n876), .B2(new_n733), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n842), .A2(new_n735), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n744), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT109), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n874), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT109), .B1(new_n844), .B2(new_n855), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n873), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n871), .B(new_n872), .C1(KEYINPUT53), .C2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n881), .B1(new_n874), .B2(new_n880), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n844), .A2(new_n855), .A3(KEYINPUT109), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n856), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n869), .A2(new_n870), .ZN(new_n889));
  OAI22_X1  g703(.A1(new_n888), .A2(new_n889), .B1(new_n884), .B2(new_n856), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n885), .B(KEYINPUT111), .C1(new_n890), .C2(new_n872), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n882), .A2(new_n883), .ZN(new_n892));
  INV_X1    g706(.A(new_n873), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT53), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT111), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n892), .B(new_n856), .C1(new_n869), .C2(new_n870), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .A4(KEYINPUT54), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n835), .B1(new_n891), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(G952), .A2(G953), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n789), .B1(new_n899), .B2(new_n900), .ZN(G75));
  NOR2_X1   g715(.A1(new_n281), .A2(G952), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n347), .A2(new_n344), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n322), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n871), .B1(new_n884), .B2(KEYINPUT53), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(G902), .A3(new_n371), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n908), .A3(new_n905), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT116), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT116), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n907), .A2(new_n912), .A3(new_n908), .A4(new_n905), .ZN(new_n913));
  AOI211_X1 g727(.A(new_n902), .B(new_n909), .C1(new_n911), .C2(new_n913), .ZN(G51));
  XOR2_X1   g728(.A(new_n767), .B(KEYINPUT57), .Z(new_n915));
  NAND2_X1  g729(.A1(new_n894), .A2(new_n856), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n872), .B1(new_n916), .B2(new_n871), .ZN(new_n917));
  INV_X1    g731(.A(new_n885), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n284), .A2(new_n297), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n906), .A2(G902), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n922), .A2(new_n766), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n902), .B1(new_n921), .B2(new_n923), .ZN(G54));
  NAND2_X1  g738(.A1(KEYINPUT58), .A2(G475), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT117), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n906), .A2(G902), .A3(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n453), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT118), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n902), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n927), .B2(new_n928), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n931), .A2(new_n933), .ZN(G60));
  NAND2_X1  g748(.A1(G478), .A2(G902), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT59), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n891), .A2(new_n898), .A3(new_n936), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n619), .A2(new_n621), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT119), .ZN(new_n940));
  INV_X1    g754(.A(new_n938), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n936), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n906), .A2(KEYINPUT54), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(new_n885), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n940), .B1(new_n944), .B2(new_n902), .ZN(new_n945));
  INV_X1    g759(.A(new_n942), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n917), .B2(new_n918), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n947), .A2(KEYINPUT119), .A3(new_n932), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n939), .A2(new_n945), .A3(new_n948), .ZN(G63));
  NAND2_X1  g763(.A1(G217), .A2(G902), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT60), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n645), .B(KEYINPUT121), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n906), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n932), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n596), .B1(new_n906), .B2(new_n952), .ZN(new_n956));
  OAI211_X1 g770(.A(KEYINPUT120), .B(KEYINPUT61), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n951), .B1(new_n916), .B2(new_n871), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n932), .B(new_n954), .C1(new_n959), .C2(new_n596), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT61), .B1(new_n960), .B2(KEYINPUT120), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n958), .A2(new_n961), .ZN(G66));
  NAND2_X1  g776(.A1(new_n855), .A2(new_n281), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT122), .Z(new_n964));
  OAI21_X1  g778(.A(G953), .B1(new_n508), .B2(new_n319), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n903), .B1(G898), .B2(new_n281), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(G69));
  AOI21_X1  g782(.A(new_n281), .B1(G227), .B2(G900), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n969), .A2(KEYINPUT125), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT126), .Z(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n528), .A2(new_n532), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(new_n440), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT62), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n866), .A2(new_n697), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n975), .B1(new_n694), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n976), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n978), .A2(KEYINPUT62), .A3(new_n693), .A4(new_n691), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n802), .B1(new_n848), .B2(new_n625), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n836), .A2(new_n675), .A3(new_n981), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT123), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n775), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n980), .A2(new_n781), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n974), .B1(new_n985), .B2(new_n281), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT124), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n978), .A2(new_n742), .A3(new_n744), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n990), .A2(new_n775), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n773), .A2(new_n774), .ZN(new_n992));
  NOR4_X1   g806(.A1(new_n795), .A2(new_n456), .A3(new_n677), .A4(new_n670), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n991), .A2(new_n781), .A3(new_n281), .A4(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n974), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n996), .B1(G900), .B2(G953), .ZN(new_n997));
  AOI22_X1  g811(.A1(new_n995), .A2(new_n997), .B1(KEYINPUT125), .B2(new_n969), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n998), .B1(new_n986), .B2(new_n987), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n972), .B1(new_n989), .B2(new_n999), .ZN(new_n1000));
  OR2_X1    g814(.A1(new_n986), .A2(new_n987), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n1001), .A2(new_n971), .A3(new_n988), .A4(new_n998), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n1000), .A2(new_n1002), .ZN(G72));
  INV_X1    g817(.A(new_n679), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n678), .A2(new_n522), .ZN(new_n1005));
  XNOR2_X1  g819(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1006));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1004), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n890), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1008), .B1(new_n985), .B2(new_n855), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n679), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n932), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1005), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n991), .A2(new_n781), .A3(new_n994), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1008), .B1(new_n1015), .B2(new_n855), .ZN(new_n1016));
  AOI211_X1 g830(.A(new_n1010), .B(new_n1013), .C1(new_n1014), .C2(new_n1016), .ZN(G57));
endmodule


