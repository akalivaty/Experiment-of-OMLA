//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n540, new_n541, new_n542, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT67), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT68), .Z(G217));
  NOR4_X1   g026(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  OR2_X1    g030(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT69), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  NAND2_X1  g033(.A1(new_n453), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n455), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n463), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n467), .A2(new_n463), .A3(new_n468), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n465), .A2(new_n466), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI211_X1 g049(.A(new_n469), .B(new_n470), .C1(G2105), .C2(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n472), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n472), .A2(new_n464), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  OAI211_X1 g058(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n484));
  OR2_X1    g059(.A1(G102), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n485), .A2(new_n487), .A3(G2104), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT71), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n484), .A2(KEYINPUT71), .A3(new_n488), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n494), .B1(new_n465), .B2(new_n466), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT3), .B(G2104), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(new_n498), .A3(new_n494), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n491), .A2(new_n492), .B1(new_n496), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  OR2_X1    g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G62), .ZN(new_n505));
  NAND2_X1  g080(.A1(G75), .A2(G543), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n501), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT72), .B(G88), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n504), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n508), .A2(G50), .A3(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n507), .A2(new_n512), .ZN(G166));
  INV_X1    g088(.A(new_n504), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n508), .A2(G89), .ZN(new_n515));
  NAND2_X1  g090(.A1(G63), .A2(G651), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n508), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G51), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n517), .A2(new_n522), .ZN(G168));
  AOI22_X1  g098(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n524), .A2(new_n501), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n504), .A2(new_n508), .ZN(new_n526));
  INV_X1    g101(.A(G90), .ZN(new_n527));
  INV_X1    g102(.A(G52), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n526), .A2(new_n527), .B1(new_n520), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n525), .A2(new_n529), .ZN(G171));
  AOI22_X1  g105(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n501), .ZN(new_n532));
  INV_X1    g107(.A(G81), .ZN(new_n533));
  XOR2_X1   g108(.A(KEYINPUT73), .B(G43), .Z(new_n534));
  OAI22_X1  g109(.A1(new_n526), .A2(new_n533), .B1(new_n520), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G860), .ZN(G153));
  NAND4_X1  g112(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n538));
  XOR2_X1   g113(.A(new_n538), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g114(.A1(G1), .A2(G3), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT75), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT8), .ZN(new_n542));
  NAND4_X1  g117(.A1(G319), .A2(G483), .A3(G661), .A4(new_n542), .ZN(G188));
  NAND2_X1  g118(.A1(G78), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G65), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n514), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT76), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n546), .A2(new_n547), .A3(G651), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n549));
  OAI21_X1  g124(.A(KEYINPUT76), .B1(new_n549), .B2(new_n501), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G53), .ZN(new_n552));
  OAI21_X1  g127(.A(KEYINPUT9), .B1(new_n520), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n508), .A2(new_n554), .A3(G53), .A4(G543), .ZN(new_n555));
  INV_X1    g130(.A(new_n526), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n553), .A2(new_n555), .B1(G91), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n551), .A2(new_n557), .ZN(G299));
  OR2_X1    g133(.A1(new_n525), .A2(new_n529), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(G171), .A2(KEYINPUT77), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(G301));
  INV_X1    g139(.A(G168), .ZN(G286));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n566), .B1(new_n507), .B2(new_n512), .ZN(new_n567));
  INV_X1    g142(.A(G62), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n568), .B1(new_n502), .B2(new_n503), .ZN(new_n569));
  INV_X1    g144(.A(new_n506), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n571), .A2(KEYINPUT78), .A3(new_n511), .A4(new_n510), .ZN(new_n572));
  AND2_X1   g147(.A1(new_n567), .A2(new_n572), .ZN(G303));
  AND2_X1   g148(.A1(new_n556), .A2(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n575));
  INV_X1    g150(.A(G49), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n576), .B2(new_n520), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(KEYINPUT79), .ZN(new_n580));
  OR3_X1    g155(.A1(new_n574), .A2(new_n577), .A3(KEYINPUT79), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G288));
  AOI22_X1  g158(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n501), .ZN(new_n585));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  INV_X1    g161(.A(G48), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n526), .A2(new_n586), .B1(new_n520), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT80), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n501), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n526), .A2(new_n594), .B1(new_n520), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n563), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT81), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n556), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n526), .B2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n520), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n602), .A2(new_n605), .B1(G54), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n501), .B1(new_n608), .B2(KEYINPUT82), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(KEYINPUT82), .B2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n601), .B1(G868), .B2(new_n613), .ZN(G284));
  OAI21_X1  g189(.A(new_n601), .B1(G868), .B2(new_n613), .ZN(G321));
  NAND2_X1  g190(.A1(G299), .A2(new_n599), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(new_n599), .B2(G168), .ZN(G297));
  OAI21_X1  g192(.A(new_n616), .B1(new_n599), .B2(G168), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n613), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n613), .A2(new_n619), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  OR3_X1    g197(.A1(new_n622), .A2(KEYINPUT84), .A3(new_n599), .ZN(new_n623));
  OAI21_X1  g198(.A(KEYINPUT84), .B1(new_n622), .B2(new_n599), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n623), .B(new_n624), .C1(G868), .C2(new_n536), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n476), .A2(G135), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n478), .A2(G123), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n464), .A2(G111), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G2096), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  INV_X1    g211(.A(G2100), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n633), .A2(new_n638), .A3(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT86), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2430), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G1341), .B(G1348), .Z(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n651), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(G14), .A3(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G401));
  INV_X1    g233(.A(KEYINPUT18), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n659), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(new_n637), .ZN(new_n666));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n662), .B2(KEYINPUT18), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(new_n632), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(new_n669), .ZN(G227));
  XOR2_X1   g245(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1956), .B(G2474), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1961), .B(G1966), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT20), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n674), .A2(new_n675), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n673), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n676), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n678), .B(new_n680), .C1(new_n673), .C2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT88), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n682), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1991), .B(G1996), .Z(new_n686));
  XOR2_X1   g261(.A(new_n685), .B(new_n686), .Z(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n685), .B(new_n686), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(new_n688), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n690), .A2(new_n692), .ZN(G229));
  NAND2_X1  g268(.A1(G305), .A2(G16), .ZN(new_n694));
  INV_X1    g269(.A(G6), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n694), .B1(new_n695), .B2(G16), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT32), .B(G1981), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n697), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n694), .B(new_n699), .C1(new_n695), .C2(G16), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G22), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G166), .B2(new_n701), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(G1971), .Z(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(G23), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n578), .B2(new_n701), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT33), .B(G1976), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  AND4_X1   g283(.A1(new_n698), .A2(new_n700), .A3(new_n704), .A4(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT34), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g286(.A1(new_n698), .A2(new_n700), .A3(new_n704), .A4(new_n708), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(KEYINPUT34), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT89), .B(G29), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n714), .A2(G25), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n476), .A2(G131), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n478), .A2(G119), .ZN(new_n717));
  OR2_X1    g292(.A1(G95), .A2(G2105), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n718), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n719));
  AND3_X1   g294(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n715), .B1(new_n720), .B2(new_n714), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT90), .Z(new_n722));
  XOR2_X1   g297(.A(KEYINPUT35), .B(G1991), .Z(new_n723));
  OR2_X1    g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n701), .A2(G24), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n597), .B2(new_n701), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(G1986), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(G1986), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n724), .A2(new_n725), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n711), .A2(new_n713), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(KEYINPUT36), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n730), .B1(new_n709), .B2(new_n710), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT36), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n734), .A2(new_n735), .A3(new_n713), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(G171), .A2(new_n701), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G5), .B2(new_n701), .ZN(new_n739));
  INV_X1    g314(.A(G1961), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT96), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n714), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G26), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT28), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n476), .A2(G140), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n478), .A2(G128), .ZN(new_n748));
  OR2_X1    g323(.A1(G104), .A2(G2105), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n749), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n750));
  AND3_X1   g325(.A1(new_n747), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G29), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n746), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G2067), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n741), .A2(new_n742), .ZN(new_n756));
  AND3_X1   g331(.A1(new_n743), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n482), .A2(new_n714), .ZN(new_n758));
  INV_X1    g333(.A(G35), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n714), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT99), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT29), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G2090), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n701), .A2(G20), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G299), .B2(G16), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1956), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n497), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(new_n464), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n476), .A2(G139), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT25), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n777), .A2(KEYINPUT92), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(KEYINPUT92), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n772), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  MUX2_X1   g355(.A(G33), .B(new_n780), .S(G29), .Z(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(G2072), .Z(new_n782));
  NAND4_X1  g357(.A1(new_n757), .A2(new_n765), .A3(new_n770), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n536), .A2(new_n701), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n701), .B2(G19), .ZN(new_n785));
  INV_X1    g360(.A(G1341), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT31), .B(G11), .Z(new_n788));
  NOR2_X1   g363(.A1(new_n631), .A2(new_n744), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT30), .B(G28), .ZN(new_n790));
  AOI211_X1 g365(.A(new_n788), .B(new_n789), .C1(new_n752), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n701), .A2(G21), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G168), .B2(new_n701), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT95), .B(G1966), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n786), .B2(new_n785), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n752), .A2(G32), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n478), .A2(G129), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT94), .ZN(new_n800));
  AND3_X1   g375(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n801));
  NAND3_X1  g376(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT26), .ZN(new_n803));
  AOI211_X1 g378(.A(new_n801), .B(new_n803), .C1(G141), .C2(new_n476), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n798), .B1(new_n805), .B2(G29), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT27), .B(G1996), .ZN(new_n807));
  AOI211_X1 g382(.A(new_n792), .B(new_n797), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(G160), .A2(G29), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT24), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(G34), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(G34), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n744), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(G2084), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(KEYINPUT93), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(KEYINPUT93), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n814), .A2(new_n815), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n739), .A2(new_n740), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n819), .B(new_n820), .C1(new_n806), .C2(new_n807), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT97), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n817), .A2(new_n818), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n744), .A2(G27), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT98), .Z(new_n826));
  NAND2_X1  g401(.A1(new_n496), .A2(new_n499), .ZN(new_n827));
  AND3_X1   g402(.A1(new_n484), .A2(KEYINPUT71), .A3(new_n488), .ZN(new_n828));
  AOI21_X1  g403(.A(KEYINPUT71), .B1(new_n484), .B2(new_n488), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n826), .B1(new_n830), .B2(new_n714), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G2078), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n808), .A2(new_n823), .A3(new_n824), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(G4), .A2(G16), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n613), .B2(G16), .ZN(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT91), .B(G1348), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n783), .A2(new_n833), .A3(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n737), .A2(new_n838), .ZN(G311));
  AOI21_X1  g414(.A(new_n735), .B1(new_n734), .B2(new_n713), .ZN(new_n840));
  AND4_X1   g415(.A1(new_n735), .A2(new_n711), .A3(new_n713), .A4(new_n731), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n838), .B(KEYINPUT101), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(KEYINPUT101), .B1(new_n737), .B2(new_n838), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(G150));
  AOI22_X1  g420(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(new_n501), .ZN(new_n847));
  INV_X1    g422(.A(G93), .ZN(new_n848));
  INV_X1    g423(.A(G55), .ZN(new_n849));
  OAI22_X1  g424(.A1(new_n526), .A2(new_n848), .B1(new_n520), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(G860), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT37), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n611), .B(KEYINPUT83), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n855), .A2(new_n619), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT38), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n847), .A2(new_n850), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(KEYINPUT102), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT102), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n851), .A2(new_n860), .ZN(new_n861));
  AND3_X1   g436(.A1(new_n859), .A2(new_n536), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n536), .B1(new_n859), .B2(new_n861), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n857), .B(new_n864), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n865), .A2(KEYINPUT39), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n852), .B1(new_n865), .B2(KEYINPUT39), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n854), .B1(new_n866), .B2(new_n867), .ZN(G145));
  INV_X1    g443(.A(KEYINPUT40), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n478), .A2(G130), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n464), .A2(G118), .ZN(new_n871));
  OAI21_X1  g446(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(G142), .B2(new_n476), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n635), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(new_n720), .Z(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n489), .B1(new_n496), .B2(new_n499), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n780), .A2(KEYINPUT104), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n880), .B(new_n772), .C1(new_n778), .C2(new_n779), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n879), .A2(new_n751), .A3(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n751), .B1(new_n879), .B2(new_n881), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n878), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n884), .ZN(new_n886));
  INV_X1    g461(.A(new_n489), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n827), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n888), .A3(new_n882), .ZN(new_n889));
  INV_X1    g464(.A(new_n805), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n885), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n890), .B1(new_n885), .B2(new_n889), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n877), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n888), .B1(new_n886), .B2(new_n882), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n883), .A2(new_n884), .A3(new_n878), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n805), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n885), .A2(new_n889), .A3(new_n890), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n897), .A3(new_n876), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n631), .B(KEYINPUT103), .Z(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(G160), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(G162), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n893), .A2(new_n898), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n876), .A2(KEYINPUT105), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n891), .B2(new_n892), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n876), .A2(KEYINPUT105), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(new_n896), .A3(new_n897), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n902), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n869), .B1(new_n905), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n907), .A2(new_n909), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n901), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n913), .A2(KEYINPUT40), .A3(new_n904), .A4(new_n903), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n911), .A2(new_n914), .ZN(G395));
  NOR2_X1   g490(.A1(new_n858), .A2(G868), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n578), .B(G166), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT107), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n597), .B(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(G305), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n589), .B(KEYINPUT80), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n597), .B(KEYINPUT107), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n917), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n920), .A2(new_n923), .A3(new_n917), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(KEYINPUT108), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n928));
  INV_X1    g503(.A(new_n926), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n928), .B1(new_n929), .B2(new_n924), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n931), .A2(KEYINPUT42), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n929), .A2(new_n924), .A3(KEYINPUT42), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n621), .B(new_n864), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n611), .A2(G299), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n611), .A2(G299), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT106), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT41), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n936), .A2(KEYINPUT41), .A3(new_n937), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n940), .B1(new_n945), .B2(new_n935), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT109), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n940), .B(KEYINPUT109), .C1(new_n945), .C2(new_n935), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n934), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n946), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n951), .B(KEYINPUT109), .C1(new_n933), .C2(new_n932), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n916), .B1(new_n953), .B2(G868), .ZN(G295));
  AOI21_X1  g529(.A(new_n916), .B1(new_n953), .B2(G868), .ZN(G331));
  NAND2_X1  g530(.A1(new_n859), .A2(new_n861), .ZN(new_n956));
  INV_X1    g531(.A(new_n536), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n859), .A2(new_n536), .A3(new_n861), .ZN(new_n959));
  AOI21_X1  g534(.A(G286), .B1(new_n561), .B2(new_n562), .ZN(new_n960));
  NOR2_X1   g535(.A1(G171), .A2(G168), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n958), .B(new_n959), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n563), .A2(G168), .ZN(new_n963));
  INV_X1    g538(.A(new_n961), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n963), .B(new_n964), .C1(new_n862), .C2(new_n863), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n962), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n960), .A2(new_n961), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n968), .B(KEYINPUT110), .C1(new_n862), .C2(new_n863), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n938), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n962), .A2(new_n965), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n945), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n972), .A2(KEYINPUT111), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n938), .B1(new_n967), .B2(new_n969), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n944), .B1(new_n962), .B2(new_n965), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n927), .A2(new_n930), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n975), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n970), .A2(new_n971), .B1(new_n945), .B2(new_n973), .ZN(new_n982));
  AOI21_X1  g557(.A(G37), .B1(new_n982), .B2(new_n931), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT43), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  OAI22_X1  g559(.A1(new_n970), .A2(new_n944), .B1(new_n939), .B2(new_n973), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n980), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n983), .A2(KEYINPUT43), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT44), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n990), .B1(new_n981), .B2(new_n983), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n972), .A2(new_n931), .A3(new_n974), .ZN(new_n992));
  AND4_X1   g567(.A1(new_n990), .A2(new_n986), .A3(new_n904), .A4(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n989), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n988), .A2(new_n994), .ZN(G397));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(new_n878), .B2(G1384), .ZN(new_n997));
  INV_X1    g572(.A(G40), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n998), .B1(new_n474), .B2(G2105), .ZN(new_n999));
  INV_X1    g574(.A(new_n469), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n467), .A2(new_n463), .A3(new_n468), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  OR2_X1    g578(.A1(new_n1003), .A2(KEYINPUT112), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(KEYINPUT112), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1996), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n805), .B(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n751), .B(G2067), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n720), .A2(new_n723), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n720), .A2(new_n723), .ZN(new_n1013));
  OR3_X1    g588(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  XOR2_X1   g589(.A(new_n597), .B(G1986), .Z(new_n1015));
  OAI21_X1  g590(.A(new_n1007), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n996), .A2(G1384), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n830), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n471), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1019), .B1(new_n497), .B2(G125), .ZN(new_n1020));
  OAI21_X1  g595(.A(G40), .B1(new_n1020), .B2(new_n464), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n1021), .A2(new_n469), .A3(new_n470), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1018), .A2(new_n997), .A3(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1023), .A2(KEYINPUT119), .A3(new_n795), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1384), .B1(new_n827), .B2(new_n887), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1002), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1384), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n830), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT50), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1027), .A2(new_n1030), .A3(new_n815), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1024), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT119), .B1(new_n1023), .B2(new_n795), .ZN(new_n1033));
  OAI21_X1  g608(.A(G286), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1023), .A2(new_n795), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1037), .A2(G168), .A3(new_n1031), .A4(new_n1024), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1034), .A2(G8), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT51), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT62), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1038), .A2(new_n1042), .A3(G8), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n567), .A2(G8), .A3(new_n572), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(KEYINPUT55), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n567), .A2(G8), .A3(new_n572), .A4(new_n1051), .ZN(new_n1052));
  XOR2_X1   g627(.A(KEYINPUT113), .B(G1971), .Z(new_n1053));
  OAI21_X1  g628(.A(new_n996), .B1(G164), .B2(G1384), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1017), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n827), .B2(new_n887), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1002), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1053), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n830), .A2(new_n1025), .A3(new_n1028), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT50), .B1(new_n878), .B2(G1384), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(new_n1022), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(G2090), .B1(new_n1061), .B2(KEYINPUT118), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1059), .A2(new_n1063), .A3(new_n1060), .A4(new_n1022), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1058), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G8), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1048), .B(new_n1052), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1048), .A2(new_n1052), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n888), .A2(new_n1025), .A3(new_n1028), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n1022), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1025), .B1(new_n830), .B2(new_n1028), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1070), .A2(new_n1071), .A3(G2090), .ZN(new_n1072));
  OAI211_X1 g647(.A(G8), .B(new_n1068), .C1(new_n1072), .C2(new_n1058), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1053), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT45), .B1(new_n830), .B2(new_n1028), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n470), .A2(new_n469), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1078), .B(new_n999), .C1(new_n878), .C2(new_n1055), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1076), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(G2090), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1082), .A2(KEYINPUT115), .A3(G8), .A4(new_n1068), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1075), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G1976), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n580), .A2(new_n1085), .A3(new_n581), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1066), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n578), .A2(G1976), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT52), .ZN(new_n1092));
  XOR2_X1   g667(.A(KEYINPUT116), .B(G1981), .Z(new_n1093));
  NAND2_X1  g668(.A1(new_n589), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(G1981), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1094), .B1(new_n1095), .B2(new_n589), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT49), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1094), .B(KEYINPUT49), .C1(new_n1095), .C2(new_n589), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(new_n1087), .A3(new_n1099), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1090), .A2(new_n1092), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(G2078), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT53), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1023), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n740), .B2(new_n1081), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1054), .A2(new_n1057), .A3(new_n1102), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(G301), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  AND4_X1   g684(.A1(new_n1067), .A2(new_n1084), .A3(new_n1101), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1044), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1111), .B1(new_n1044), .B2(new_n1110), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1041), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1084), .A2(new_n1067), .A3(new_n1101), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1104), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n740), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1108), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n563), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1081), .A2(new_n1122), .A3(new_n740), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1118), .A2(KEYINPUT122), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AND2_X1   g700(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1126));
  NOR2_X1   g701(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1127));
  OAI211_X1 g702(.A(KEYINPUT53), .B(G40), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1056), .A2(new_n1128), .ZN(new_n1129));
  AND3_X1   g704(.A1(G160), .A2(new_n1129), .A3(new_n997), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1130), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1125), .A2(G301), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT54), .B1(new_n1121), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n559), .B1(new_n1125), .B2(new_n1131), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1117), .A2(new_n1108), .A3(G301), .A4(new_n1118), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(KEYINPUT54), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1116), .A2(new_n1133), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(G1348), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1022), .A2(new_n1026), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1140), .B1(G2067), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n855), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(G1348), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1141), .A2(G2067), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1147), .A2(KEYINPUT60), .A3(new_n613), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1144), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT56), .B(G2072), .ZN(new_n1152));
  INV_X1    g727(.A(G1956), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1151), .A2(new_n1152), .B1(new_n1061), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT57), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n551), .A2(new_n1155), .A3(new_n557), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1155), .B1(new_n551), .B2(new_n557), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(KEYINPUT121), .B1(new_n1154), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1061), .A2(new_n1153), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1159), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT121), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT61), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1167), .B1(new_n1154), .B2(new_n1159), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1160), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1159), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1159), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1167), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1054), .A2(new_n1057), .A3(new_n1008), .ZN(new_n1173));
  XOR2_X1   g748(.A(KEYINPUT58), .B(G1341), .Z(new_n1174));
  NAND2_X1  g749(.A1(new_n1141), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n957), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT59), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1176), .B(new_n1177), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1150), .A2(new_n1169), .A3(new_n1172), .A4(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1166), .A2(new_n1160), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1147), .A2(new_n855), .ZN(new_n1181));
  OAI22_X1  g756(.A1(new_n1180), .A2(new_n1181), .B1(new_n1164), .B2(new_n1163), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1138), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT63), .ZN(new_n1186));
  NOR2_X1   g761(.A1(G286), .A2(new_n1066), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1187), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1186), .B1(new_n1116), .B2(new_n1188), .ZN(new_n1189));
  OAI211_X1 g764(.A(KEYINPUT63), .B(new_n1187), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1068), .B1(new_n1082), .B2(G8), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1192), .A2(new_n1084), .A3(new_n1101), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT120), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1192), .A2(new_n1084), .A3(KEYINPUT120), .A4(new_n1101), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1189), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1084), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1100), .A2(new_n1085), .A3(new_n582), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n1094), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1087), .B(KEYINPUT117), .ZN(new_n1201));
  AOI22_X1  g776(.A1(new_n1198), .A2(new_n1101), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1185), .A2(new_n1197), .A3(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1016), .B1(new_n1115), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1006), .B1(new_n890), .B2(new_n1010), .ZN(new_n1205));
  OR3_X1    g780(.A1(new_n1006), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1206));
  OAI21_X1  g781(.A(KEYINPUT46), .B1(new_n1006), .B2(G1996), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1205), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(KEYINPUT47), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1210));
  AOI22_X1  g785(.A1(new_n1210), .A2(new_n1013), .B1(new_n754), .B2(new_n751), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1007), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1213), .B1(new_n1212), .B2(new_n1211), .ZN(new_n1214));
  OR3_X1    g789(.A1(new_n1006), .A2(G1986), .A3(G290), .ZN(new_n1215));
  XNOR2_X1  g790(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1216));
  OR2_X1    g791(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  AOI22_X1  g792(.A1(new_n1014), .A2(new_n1007), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1218));
  AOI211_X1 g793(.A(new_n1209), .B(new_n1214), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1204), .A2(new_n1219), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g795(.A1(new_n991), .A2(new_n993), .ZN(new_n1222));
  OR2_X1    g796(.A1(G227), .A2(new_n461), .ZN(new_n1223));
  INV_X1    g797(.A(KEYINPUT127), .ZN(new_n1224));
  OR2_X1    g798(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g799(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1226));
  NAND3_X1  g800(.A1(new_n1225), .A2(new_n657), .A3(new_n1226), .ZN(new_n1227));
  AOI21_X1  g801(.A(new_n1227), .B1(new_n690), .B2(new_n692), .ZN(new_n1228));
  OAI21_X1  g802(.A(new_n1228), .B1(new_n905), .B2(new_n910), .ZN(new_n1229));
  NOR2_X1   g803(.A1(new_n1222), .A2(new_n1229), .ZN(G308));
  OAI221_X1 g804(.A(new_n1228), .B1(new_n905), .B2(new_n910), .C1(new_n991), .C2(new_n993), .ZN(G225));
endmodule


