//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1214, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  OR2_X1    g0003(.A1(new_n203), .A2(KEYINPUT64), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(KEYINPUT64), .ZN(new_n205));
  NAND3_X1  g0005(.A1(new_n204), .A2(G50), .A3(new_n205), .ZN(new_n206));
  NAND3_X1  g0006(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n208), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n213), .B1(new_n209), .B2(new_n212), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT65), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G87), .A2(G250), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI211_X1 g0022(.A(new_n218), .B(new_n222), .C1(G107), .C2(G264), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G50), .A2(G226), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G77), .A2(G244), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G116), .A2(G270), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G58), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n210), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n215), .A2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G264), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(KEYINPUT66), .B(G107), .ZN(new_n242));
  INV_X1    g0042(.A(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XOR2_X1   g0047(.A(G50), .B(G58), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(new_n203), .ZN(new_n251));
  OAI21_X1  g0051(.A(G20), .B1(new_n251), .B2(G50), .ZN(new_n252));
  INV_X1    g0052(.A(G150), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT8), .A2(G58), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT68), .B(G58), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n256), .B1(new_n257), .B2(KEYINPUT8), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G20), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G33), .ZN(new_n261));
  OAI221_X1 g0061(.A(new_n252), .B1(new_n253), .B2(new_n255), .C1(new_n259), .C2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G1), .A2(G13), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G50), .ZN(new_n266));
  INV_X1    g0066(.A(G13), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G1), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G20), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n262), .A2(new_n265), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G1), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n265), .B1(new_n272), .B2(G20), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G50), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT9), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  OAI211_X1 g0078(.A(G1), .B(G13), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT3), .B(G33), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(G222), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT67), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n281), .A2(G1698), .ZN(new_n286));
  INV_X1    g0086(.A(G223), .ZN(new_n287));
  INV_X1    g0087(.A(G77), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n286), .A2(new_n287), .B1(new_n288), .B2(new_n281), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n280), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n272), .B1(G41), .B2(G45), .ZN(new_n291));
  INV_X1    g0091(.A(G274), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n279), .A2(new_n291), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G226), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n290), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n275), .A2(new_n276), .B1(G200), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n271), .A2(KEYINPUT9), .A3(new_n274), .ZN(new_n299));
  INV_X1    g0099(.A(new_n297), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G190), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n298), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n298), .A2(new_n299), .A3(new_n304), .A4(new_n301), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n279), .A2(G238), .A3(new_n291), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n293), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT70), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n307), .A2(new_n293), .A3(KEYINPUT70), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n281), .A2(G226), .A3(new_n282), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G97), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n312), .B(new_n313), .C1(new_n286), .C2(new_n229), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n310), .A2(new_n311), .B1(new_n314), .B2(new_n280), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT13), .ZN(new_n316));
  INV_X1    g0116(.A(G200), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n268), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n216), .A2(G20), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n321), .B(KEYINPUT12), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n322), .B1(G68), .B2(new_n273), .ZN(new_n323));
  OAI221_X1 g0123(.A(new_n320), .B1(new_n261), .B2(new_n288), .C1(new_n255), .C2(new_n266), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n265), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT11), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n310), .A2(new_n311), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n314), .A2(new_n280), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT13), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n315), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G190), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n328), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n318), .A2(new_n337), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n316), .A2(G179), .B1(KEYINPUT71), .B2(KEYINPUT14), .ZN(new_n339));
  NOR2_X1   g0139(.A1(KEYINPUT71), .A2(KEYINPUT14), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G169), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n341), .B1(new_n316), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n335), .A2(G169), .A3(new_n340), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n339), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n338), .B1(new_n345), .B2(new_n327), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n297), .A2(new_n342), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n347), .B(new_n275), .C1(G179), .C2(new_n297), .ZN(new_n348));
  XNOR2_X1  g0148(.A(KEYINPUT8), .B(G58), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n349), .A2(new_n255), .B1(new_n260), .B2(new_n288), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT15), .B(G87), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n261), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(new_n265), .B1(new_n288), .B2(new_n270), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n273), .A2(G77), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n356), .A2(KEYINPUT69), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(KEYINPUT69), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n281), .A2(G232), .A3(new_n282), .ZN(new_n359));
  INV_X1    g0159(.A(G107), .ZN(new_n360));
  OAI221_X1 g0160(.A(new_n359), .B1(new_n360), .B2(new_n281), .C1(new_n286), .C2(new_n217), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n280), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n295), .A2(G244), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(new_n293), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n357), .A2(new_n358), .B1(G190), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(G200), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n306), .A2(new_n346), .A3(new_n348), .A4(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT72), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n228), .A2(KEYINPUT68), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT68), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G58), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n373), .A3(G68), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n260), .B1(new_n374), .B2(new_n251), .ZN(new_n375));
  INV_X1    g0175(.A(G159), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n255), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n370), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n377), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n203), .B1(new_n257), .B2(G68), .ZN(new_n380));
  OAI211_X1 g0180(.A(KEYINPUT72), .B(new_n379), .C1(new_n380), .C2(new_n260), .ZN(new_n381));
  AND2_X1   g0181(.A1(KEYINPUT3), .A2(G33), .ZN(new_n382));
  NOR2_X1   g0182(.A1(KEYINPUT3), .A2(G33), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT7), .B1(new_n384), .B2(new_n260), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  NOR4_X1   g0186(.A1(new_n382), .A2(new_n383), .A3(new_n386), .A4(G20), .ZN(new_n387));
  OAI21_X1  g0187(.A(G68), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n378), .A2(new_n381), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT16), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n378), .A2(new_n381), .A3(KEYINPUT16), .A4(new_n388), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(new_n265), .A3(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n258), .A2(new_n269), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n258), .B1(G1), .B2(new_n260), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n395), .B(KEYINPUT73), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n270), .A2(new_n265), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n287), .A2(new_n282), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n281), .B(new_n399), .C1(G226), .C2(new_n282), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G33), .A2(G87), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n279), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n293), .B1(new_n294), .B2(new_n229), .ZN(new_n403));
  OAI21_X1  g0203(.A(G200), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n402), .A2(new_n403), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G190), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n393), .A2(new_n398), .A3(new_n404), .A4(new_n406), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT17), .ZN(new_n408));
  INV_X1    g0208(.A(G179), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(G169), .B2(new_n405), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(new_n393), .B2(new_n398), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n412), .B(KEYINPUT18), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n365), .A2(new_n409), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n364), .A2(new_n342), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n356), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n408), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n369), .A2(new_n417), .ZN(new_n418));
  AND2_X1   g0218(.A1(KEYINPUT5), .A2(G41), .ZN(new_n419));
  NOR2_X1   g0219(.A1(KEYINPUT5), .A2(G41), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n272), .B(G45), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  OR2_X1    g0221(.A1(new_n421), .A2(new_n292), .ZN(new_n422));
  OAI211_X1 g0222(.A(G257), .B(G1698), .C1(new_n382), .C2(new_n383), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT82), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT82), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n281), .A2(new_n425), .A3(G257), .A4(G1698), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n281), .A2(G250), .A3(new_n282), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G294), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n280), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n421), .A2(G264), .A3(new_n279), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT84), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT84), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n421), .A2(new_n434), .A3(G264), .A4(new_n279), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n431), .A2(KEYINPUT85), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT85), .B1(new_n431), .B2(new_n436), .ZN(new_n438));
  OAI211_X1 g0238(.A(G179), .B(new_n422), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT86), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n431), .A2(new_n436), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT85), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n431), .A2(KEYINPUT85), .A3(new_n436), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n446), .A2(KEYINPUT86), .A3(G179), .A4(new_n422), .ZN(new_n447));
  INV_X1    g0247(.A(new_n422), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(new_n431), .B2(KEYINPUT83), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n449), .B(new_n436), .C1(KEYINPUT83), .C2(new_n431), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G169), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n441), .A2(new_n447), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT24), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n260), .B(G87), .C1(new_n382), .C2(new_n383), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT22), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT22), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n281), .A2(new_n456), .A3(new_n260), .A4(G87), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G33), .A2(G116), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(G20), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n360), .A2(G20), .ZN(new_n462));
  XOR2_X1   g0262(.A(new_n462), .B(KEYINPUT23), .Z(new_n463));
  AND4_X1   g0263(.A1(new_n453), .A2(new_n458), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n460), .B1(new_n455), .B2(new_n457), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n453), .B1(new_n465), .B2(new_n463), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n265), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT80), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT80), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n469), .B(new_n265), .C1(new_n464), .C2(new_n466), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n277), .A2(G1), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n270), .A2(new_n265), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G107), .ZN(new_n473));
  INV_X1    g0273(.A(new_n462), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT81), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n474), .B(new_n268), .C1(new_n475), .C2(KEYINPUT25), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(KEYINPUT25), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n476), .B(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n468), .A2(new_n470), .A3(new_n473), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n452), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT74), .ZN(new_n481));
  XNOR2_X1  g0281(.A(G97), .B(G107), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT6), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n483), .A2(new_n220), .A3(G107), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n260), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n255), .A2(new_n288), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n481), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(G107), .B1(new_n385), .B2(new_n387), .ZN(new_n490));
  INV_X1    g0290(.A(new_n488), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n485), .B1(new_n483), .B2(new_n482), .ZN(new_n492));
  OAI211_X1 g0292(.A(KEYINPUT74), .B(new_n491), .C1(new_n492), .C2(new_n260), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n489), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n265), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n472), .A2(G97), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n269), .A2(G97), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n497), .B(KEYINPUT75), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n495), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n281), .A2(G244), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G283), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n281), .A2(KEYINPUT4), .A3(G244), .A4(new_n282), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n281), .A2(G250), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n282), .B1(new_n506), .B2(KEYINPUT4), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n280), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n421), .A2(new_n279), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G257), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n422), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n342), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n500), .A2(new_n501), .B1(G33), .B2(G283), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n501), .B1(new_n281), .B2(G250), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n513), .B(new_n504), .C1(new_n282), .C2(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n515), .A2(new_n280), .B1(G257), .B2(new_n509), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(new_n409), .A3(new_n422), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n499), .A2(new_n512), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n511), .A2(G200), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n494), .A2(new_n265), .B1(G97), .B2(new_n472), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n508), .A2(G190), .A3(new_n422), .A4(new_n510), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n498), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n479), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n448), .B1(new_n444), .B2(new_n445), .ZN(new_n525));
  OAI22_X1  g0325(.A1(new_n525), .A2(G200), .B1(new_n450), .B2(G190), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n523), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT21), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n503), .B(new_n260), .C1(G33), .C2(new_n220), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n243), .A2(G20), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(new_n265), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT20), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n529), .A2(KEYINPUT20), .A3(new_n265), .A4(new_n530), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n472), .A2(G116), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(G116), .B2(new_n269), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G303), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n384), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G264), .A2(G1698), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n221), .B2(G1698), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n539), .B(new_n280), .C1(new_n384), .C2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n421), .A2(G270), .A3(new_n279), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(new_n422), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G169), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n528), .B1(new_n537), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(G200), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n537), .B(new_n547), .C1(new_n336), .C2(new_n544), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n542), .A2(new_n422), .A3(G179), .A4(new_n543), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n545), .B2(new_n528), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT79), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n550), .A2(new_n551), .A3(new_n536), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n551), .B1(new_n550), .B2(new_n536), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n546), .B(new_n548), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n217), .A2(new_n282), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n281), .B(new_n555), .C1(G244), .C2(new_n282), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n279), .B1(new_n556), .B2(new_n459), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n272), .A2(G45), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n279), .A2(G250), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT77), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n279), .A2(KEYINPUT77), .A3(G250), .A4(new_n558), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n272), .A2(G45), .A3(G274), .ZN(new_n563));
  XNOR2_X1  g0363(.A(new_n563), .B(KEYINPUT76), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT78), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT78), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n561), .A2(new_n567), .A3(new_n564), .A4(new_n562), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n557), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n409), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n281), .A2(new_n260), .A3(G68), .ZN(new_n571));
  INV_X1    g0371(.A(G87), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n572), .A2(new_n220), .A3(new_n360), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n313), .A2(new_n260), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n574), .A3(KEYINPUT19), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n313), .A2(G20), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n571), .B(new_n575), .C1(KEYINPUT19), .C2(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(new_n265), .B1(new_n270), .B2(new_n351), .ZN(new_n578));
  INV_X1    g0378(.A(new_n351), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n472), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n570), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n569), .A2(G169), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n569), .A2(G190), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n472), .A2(G87), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n578), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n569), .B2(new_n317), .ZN(new_n589));
  OAI22_X1  g0389(.A1(new_n582), .A2(new_n583), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n554), .A2(new_n590), .ZN(new_n591));
  AND4_X1   g0391(.A1(new_n418), .A2(new_n480), .A3(new_n527), .A4(new_n591), .ZN(G372));
  INV_X1    g0392(.A(new_n413), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n345), .A2(new_n327), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n338), .B2(new_n416), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n593), .B1(new_n595), .B2(new_n408), .ZN(new_n596));
  INV_X1    g0396(.A(new_n306), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n348), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n583), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(new_n570), .A3(new_n581), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n518), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n566), .A2(new_n568), .ZN(new_n603));
  INV_X1    g0403(.A(new_n557), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n587), .B1(new_n605), .B2(G200), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n584), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n602), .A2(new_n607), .A3(new_n600), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n601), .B1(new_n608), .B2(KEYINPUT26), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n589), .A2(KEYINPUT87), .B1(G190), .B2(new_n569), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT87), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n582), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n610), .A2(new_n612), .B1(new_n613), .B2(new_n599), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT26), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(new_n615), .A3(new_n602), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n524), .A2(new_n526), .ZN(new_n617));
  INV_X1    g0417(.A(new_n523), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n614), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n550), .A2(new_n536), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n546), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n452), .B2(new_n479), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n609), .B(new_n616), .C1(new_n619), .C2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n598), .B1(new_n418), .B2(new_n623), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n624), .B(KEYINPUT88), .ZN(G369));
  OAI21_X1  g0425(.A(new_n546), .B1(new_n552), .B2(new_n553), .ZN(new_n626));
  OR3_X1    g0426(.A1(new_n319), .A2(KEYINPUT27), .A3(G20), .ZN(new_n627));
  OAI21_X1  g0427(.A(KEYINPUT27), .B1(new_n319), .B2(G20), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(G213), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(G343), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n441), .A2(new_n447), .A3(new_n451), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n479), .A2(new_n631), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT90), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n479), .A2(new_n631), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT90), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(new_n638), .A3(new_n452), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n480), .A2(new_n617), .A3(new_n635), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n633), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n480), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n642), .B1(new_n643), .B2(new_n632), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n634), .A2(KEYINPUT90), .A3(new_n635), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n638), .B1(new_n637), .B2(new_n452), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n641), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n537), .A2(new_n632), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n621), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n554), .B2(new_n648), .ZN(new_n650));
  XNOR2_X1  g0450(.A(KEYINPUT89), .B(G330), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n644), .A2(new_n654), .ZN(G399));
  NAND2_X1  g0455(.A1(new_n211), .A2(new_n278), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(G1), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n573), .A2(G116), .ZN(new_n658));
  OAI22_X1  g0458(.A1(new_n206), .A2(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT28), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT93), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n614), .A2(new_n602), .A3(new_n661), .A4(KEYINPUT26), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n626), .B1(new_n452), .B2(new_n479), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n662), .B(new_n600), .C1(new_n619), .C2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n614), .A2(KEYINPUT26), .A3(new_n602), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n608), .A2(new_n615), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n665), .A2(KEYINPUT93), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n632), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT29), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n623), .A2(new_n632), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT29), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT30), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n516), .B1(new_n437), .B2(new_n438), .ZN(new_n673));
  INV_X1    g0473(.A(new_n549), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n569), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n672), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  AOI211_X1 g0476(.A(new_n557), .B(new_n549), .C1(new_n566), .C2(new_n568), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n677), .A2(new_n446), .A3(KEYINPUT30), .A4(new_n516), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n422), .B1(new_n437), .B2(new_n438), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n569), .A2(KEYINPUT91), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(new_n544), .A3(new_n680), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n409), .B(new_n511), .C1(new_n569), .C2(KEYINPUT91), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n676), .B(new_n678), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n683), .A2(KEYINPUT31), .A3(new_n631), .ZN(new_n684));
  AOI21_X1  g0484(.A(KEYINPUT31), .B1(new_n683), .B2(new_n631), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT92), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(new_n631), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT31), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT92), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n683), .A2(KEYINPUT31), .A3(new_n631), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n527), .A2(new_n591), .A3(new_n480), .A4(new_n632), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n686), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n651), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n669), .A2(new_n671), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n660), .B1(new_n697), .B2(G1), .ZN(G364));
  AOI21_X1  g0498(.A(new_n264), .B1(G20), .B2(new_n342), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n260), .A2(G190), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(G179), .A3(new_n317), .ZN(new_n701));
  INV_X1    g0501(.A(G311), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g0503(.A(KEYINPUT99), .B(G317), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT33), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n409), .A2(new_n317), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n700), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n260), .A2(new_n336), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n709), .A2(G179), .A3(new_n317), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n705), .A2(new_n708), .B1(G322), .B2(new_n711), .ZN(new_n712));
  XOR2_X1   g0512(.A(new_n712), .B(KEYINPUT100), .Z(new_n713));
  NAND2_X1  g0513(.A1(new_n709), .A2(new_n706), .ZN(new_n714));
  INV_X1    g0514(.A(G326), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n384), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(G179), .A2(G200), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n260), .B1(new_n717), .B2(G190), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n716), .B1(G294), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n317), .A2(G179), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n709), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n700), .A2(new_n717), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI22_X1  g0525(.A1(G303), .A2(new_n723), .B1(new_n725), .B2(G329), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n713), .A2(new_n720), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n700), .A2(new_n721), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n703), .B(new_n727), .C1(G283), .C2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n701), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n731), .A2(KEYINPUT96), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(KEYINPUT96), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI22_X1  g0534(.A1(new_n734), .A2(new_n288), .B1(new_n220), .B2(new_n718), .ZN(new_n735));
  AOI22_X1  g0535(.A1(G68), .A2(new_n708), .B1(new_n723), .B2(G87), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n728), .A2(new_n360), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n384), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n736), .B(new_n738), .C1(new_n266), .C2(new_n714), .ZN(new_n739));
  INV_X1    g0539(.A(new_n257), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n710), .ZN(new_n741));
  XOR2_X1   g0541(.A(KEYINPUT97), .B(G159), .Z(new_n742));
  NAND2_X1  g0542(.A1(new_n725), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g0543(.A(KEYINPUT98), .B(KEYINPUT32), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NOR4_X1   g0545(.A1(new_n735), .A2(new_n739), .A3(new_n741), .A4(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n699), .B1(new_n730), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n267), .A2(G20), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G45), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n656), .A2(G1), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT94), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n281), .A2(G355), .A3(new_n211), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n384), .A2(new_n211), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT95), .Z(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(G45), .B2(new_n206), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n249), .A2(G45), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n753), .B1(G116), .B2(new_n211), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G13), .A2(G33), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G20), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n699), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n752), .B1(new_n758), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n761), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n747), .B(new_n763), .C1(new_n650), .C2(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT101), .Z(new_n766));
  NOR2_X1   g0566(.A1(new_n653), .A2(new_n751), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(new_n651), .B2(new_n650), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n766), .A2(new_n768), .ZN(G396));
  INV_X1    g0569(.A(new_n699), .ZN(new_n770));
  XOR2_X1   g0570(.A(KEYINPUT102), .B(G143), .Z(new_n771));
  AOI22_X1  g0571(.A1(new_n711), .A2(new_n771), .B1(new_n708), .B2(G150), .ZN(new_n772));
  INV_X1    g0572(.A(new_n742), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n772), .B1(new_n734), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n714), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n774), .B1(G137), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT34), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(G50), .B2(new_n723), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n384), .B1(new_n725), .B2(G132), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n719), .A2(new_n257), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n729), .A2(G68), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n778), .A2(new_n779), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n734), .A2(new_n243), .B1(new_n220), .B2(new_n718), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n728), .A2(new_n572), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(new_n702), .B2(new_n724), .ZN(new_n786));
  INV_X1    g0586(.A(G294), .ZN(new_n787));
  INV_X1    g0587(.A(G283), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n710), .A2(new_n787), .B1(new_n707), .B2(new_n788), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n786), .A2(new_n281), .A3(new_n789), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n790), .B1(new_n360), .B2(new_n722), .C1(new_n538), .C2(new_n714), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n770), .B1(new_n782), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n699), .A2(new_n759), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n752), .B(new_n792), .C1(new_n288), .C2(new_n793), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n414), .A2(new_n415), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n795), .A2(KEYINPUT103), .A3(new_n356), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT103), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n416), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n632), .B1(new_n355), .B2(new_n354), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n799), .A2(new_n368), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n795), .A2(new_n800), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT104), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n795), .A2(KEYINPUT104), .A3(new_n800), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n794), .B1(new_n760), .B2(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n796), .A2(new_n798), .B1(new_n367), .B2(new_n366), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n810), .A2(new_n801), .B1(new_n805), .B2(new_n806), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n670), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n623), .A2(new_n632), .A3(new_n808), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(new_n695), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n809), .B1(new_n815), .B2(new_n751), .ZN(G384));
  INV_X1    g0616(.A(KEYINPUT37), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n393), .A2(new_n398), .ZN(new_n818));
  INV_X1    g0618(.A(new_n629), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(KEYINPUT106), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT106), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n818), .A2(new_n822), .A3(new_n819), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n411), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n818), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n407), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n817), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n826), .A2(new_n820), .A3(new_n817), .A4(new_n407), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(KEYINPUT107), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT17), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n407), .A2(new_n833), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n393), .A2(new_n398), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n835), .A2(KEYINPUT17), .A3(new_n404), .A4(new_n406), .ZN(new_n836));
  AND3_X1   g0636(.A1(new_n818), .A2(KEYINPUT18), .A3(new_n825), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n412), .A2(KEYINPUT18), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n834), .B(new_n836), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n839), .A2(new_n821), .A3(new_n823), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT107), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n827), .B1(new_n821), .B2(new_n823), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n841), .B(new_n830), .C1(new_n842), .C2(new_n817), .ZN(new_n843));
  AND4_X1   g0643(.A1(KEYINPUT38), .A2(new_n832), .A3(new_n840), .A4(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n820), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n826), .A2(new_n820), .A3(new_n407), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(KEYINPUT37), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n839), .A2(new_n845), .B1(new_n847), .B2(new_n830), .ZN(new_n848));
  OAI21_X1  g0648(.A(KEYINPUT108), .B1(new_n848), .B2(KEYINPUT38), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT108), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n847), .A2(new_n830), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n820), .B1(new_n408), .B2(new_n413), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n850), .B(new_n851), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n844), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n345), .A2(new_n327), .A3(new_n631), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT105), .ZN(new_n858));
  INV_X1    g0658(.A(new_n338), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n327), .A2(new_n631), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n594), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n346), .A2(KEYINPUT105), .A3(new_n860), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n811), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n693), .A2(new_n689), .A3(new_n691), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT40), .B1(new_n856), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n832), .A2(new_n840), .A3(new_n843), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n851), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n832), .A2(KEYINPUT38), .A3(new_n840), .A4(new_n843), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n866), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT40), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n418), .A2(new_n865), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n875), .B(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n651), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT39), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n844), .B2(new_n855), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n869), .A2(KEYINPUT39), .A3(new_n870), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n594), .A2(new_n631), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n413), .A2(new_n819), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n862), .A2(new_n863), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n796), .A2(new_n632), .A3(new_n798), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n885), .B1(new_n813), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n884), .B1(new_n871), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n878), .B(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n418), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n669), .B2(new_n671), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n892), .A2(new_n598), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n890), .B(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n272), .B2(new_n748), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT35), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n207), .B1(new_n492), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n897), .B(G116), .C1(new_n896), .C2(new_n492), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT36), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n374), .A2(G77), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n206), .A2(new_n900), .B1(G50), .B2(new_n216), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(G1), .A3(new_n267), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n895), .A2(new_n899), .A3(new_n902), .ZN(G367));
  INV_X1    g0703(.A(new_n654), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n499), .A2(new_n631), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n618), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n518), .B2(new_n632), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT110), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT42), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n642), .B2(new_n907), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n618), .A2(new_n479), .A3(new_n452), .A4(new_n905), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n631), .B1(new_n913), .B2(new_n518), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT109), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n633), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n647), .A2(new_n916), .A3(new_n907), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT42), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT109), .ZN(new_n919));
  INV_X1    g0719(.A(new_n914), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n915), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n917), .A2(KEYINPUT42), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n910), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  AOI211_X1 g0725(.A(KEYINPUT110), .B(new_n923), .C1(new_n915), .C2(new_n921), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT111), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n588), .A2(new_n632), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n601), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n614), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n929), .B1(new_n930), .B2(new_n928), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n927), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n919), .B1(new_n918), .B2(new_n920), .ZN(new_n934));
  AOI211_X1 g0734(.A(KEYINPUT109), .B(new_n914), .C1(new_n917), .C2(KEYINPUT42), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n924), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT110), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n922), .A2(new_n910), .A3(new_n924), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n939), .A2(KEYINPUT111), .A3(new_n931), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n933), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT43), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n933), .B2(new_n941), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n909), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n644), .A2(new_n907), .ZN(new_n946));
  XOR2_X1   g0746(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n644), .A2(new_n907), .A3(new_n947), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT44), .B1(new_n644), .B2(new_n907), .ZN(new_n952));
  OR3_X1    g0752(.A1(new_n644), .A2(KEYINPUT44), .A3(new_n907), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n951), .A2(new_n654), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n647), .B(new_n916), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(new_n652), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(new_n696), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n953), .A2(new_n949), .A3(new_n952), .A4(new_n950), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n904), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n954), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n697), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n656), .B(KEYINPUT41), .Z(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n749), .A2(G1), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n931), .B1(new_n939), .B2(KEYINPUT111), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT111), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n968), .B(new_n932), .C1(new_n937), .C2(new_n938), .ZN(new_n969));
  OAI21_X1  g0769(.A(KEYINPUT43), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n933), .A2(new_n940), .A3(new_n941), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n970), .A2(new_n908), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n945), .A2(new_n966), .A3(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n722), .A2(new_n243), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n974), .A2(KEYINPUT46), .B1(new_n538), .B2(new_n710), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n729), .A2(G97), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n976), .B1(new_n787), .B2(new_n707), .C1(new_n702), .C2(new_n714), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(G107), .B2(new_n719), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n974), .A2(KEYINPUT46), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n978), .A2(new_n384), .A3(new_n979), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n975), .B(new_n980), .C1(G317), .C2(new_n725), .ZN(new_n981));
  INV_X1    g0781(.A(new_n734), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(G283), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n281), .B1(new_n718), .B2(new_n216), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n773), .A2(new_n707), .B1(new_n728), .B2(new_n288), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n984), .B(new_n985), .C1(new_n775), .C2(new_n771), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n253), .B2(new_n710), .C1(new_n740), .C2(new_n722), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G137), .B2(new_n725), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n982), .A2(G50), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n981), .A2(new_n983), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT47), .Z(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n699), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n932), .A2(new_n761), .ZN(new_n993));
  INV_X1    g0793(.A(new_n755), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n762), .B1(new_n211), .B2(new_n351), .C1(new_n236), .C2(new_n994), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n992), .A2(new_n751), .A3(new_n993), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n973), .A2(new_n996), .ZN(G387));
  INV_X1    g0797(.A(new_n957), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n656), .B1(new_n956), .B2(new_n696), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n384), .B1(new_n724), .B2(new_n715), .ZN(new_n1001));
  XOR2_X1   g0801(.A(KEYINPUT114), .B(G322), .Z(new_n1002));
  AOI22_X1  g0802(.A1(G317), .A2(new_n711), .B1(new_n775), .B2(new_n1002), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n702), .B2(new_n707), .C1(new_n734), .C2(new_n538), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT48), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n788), .B2(new_n718), .C1(new_n787), .C2(new_n722), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT49), .Z(new_n1007));
  AOI211_X1 g0807(.A(new_n1001), .B(new_n1007), .C1(G116), .C2(new_n729), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n258), .A2(new_n708), .B1(new_n731), .B2(G68), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT113), .Z(new_n1010));
  AOI22_X1  g0810(.A1(new_n775), .A2(G159), .B1(new_n725), .B2(G150), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n266), .B2(new_n710), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n722), .A2(new_n288), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n718), .A2(new_n351), .ZN(new_n1014));
  NOR3_X1   g0814(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  AND4_X1   g0815(.A1(new_n281), .A2(new_n1010), .A3(new_n1015), .A4(new_n976), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n699), .B1(new_n1008), .B2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n640), .A2(new_n641), .A3(new_n761), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n349), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n266), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT50), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n216), .A2(new_n288), .ZN(new_n1022));
  NOR4_X1   g0822(.A1(new_n1021), .A2(G45), .A3(new_n1022), .A4(new_n658), .ZN(new_n1023));
  INV_X1    g0823(.A(G45), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n755), .B1(new_n240), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n658), .A2(new_n211), .A3(new_n281), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n211), .A2(G107), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n762), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1017), .A2(new_n751), .A3(new_n1018), .A4(new_n1029), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1000), .B(new_n1030), .C1(new_n965), .C2(new_n956), .ZN(G393));
  NAND3_X1  g0831(.A1(new_n954), .A2(KEYINPUT115), .A3(new_n959), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1032), .B(new_n998), .C1(KEYINPUT115), .C2(new_n954), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n656), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n1034), .A3(new_n960), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n246), .A2(new_n755), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1036), .B(new_n762), .C1(new_n220), .C2(new_n211), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n751), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n907), .A2(new_n764), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n982), .A2(new_n1019), .B1(G68), .B2(new_n723), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n718), .A2(new_n288), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n707), .A2(new_n266), .B1(new_n728), .B2(new_n572), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n384), .B(new_n1043), .C1(new_n725), .C2(new_n771), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n710), .A2(new_n376), .B1(new_n714), .B2(new_n253), .ZN(new_n1045));
  XOR2_X1   g0845(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n1046));
  XNOR2_X1  g0846(.A(new_n1045), .B(new_n1046), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1040), .A2(new_n1042), .A3(new_n1044), .A4(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n711), .A2(G311), .B1(new_n775), .B2(G317), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT52), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n281), .B(new_n1050), .C1(G283), .C2(new_n723), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n731), .A2(G294), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n725), .A2(new_n1002), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n708), .A2(G303), .B1(new_n719), .B2(G116), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n737), .B1(new_n1054), .B2(KEYINPUT117), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1054), .A2(KEYINPUT117), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1048), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1038), .B(new_n1039), .C1(new_n699), .C2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1032), .B1(KEYINPUT115), .B2(new_n954), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1059), .B1(new_n1060), .B2(new_n964), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1035), .A2(new_n1061), .ZN(G390));
  INV_X1    g0862(.A(G330), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n876), .A2(new_n1063), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n892), .A2(new_n1064), .A3(new_n598), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n872), .A2(G330), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n885), .B1(new_n695), .B2(new_n811), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n813), .A2(new_n886), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n864), .A2(new_n694), .A3(new_n651), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n865), .A2(G330), .A3(new_n808), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n885), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n632), .B(new_n808), .C1(new_n664), .C2(new_n667), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1071), .A2(new_n1073), .A3(new_n886), .A4(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT118), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1074), .A2(new_n886), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1078), .A2(KEYINPUT118), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1070), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1066), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n880), .A2(new_n881), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n862), .A2(new_n863), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1069), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n882), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1082), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1085), .B1(new_n844), .B2(new_n855), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n885), .B1(new_n1074), .B2(new_n886), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1081), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n880), .A2(new_n881), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1093));
  NOR3_X1   g0893(.A1(new_n1092), .A2(new_n1093), .A3(new_n1071), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1065), .B(new_n1080), .C1(new_n1091), .C2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1066), .A2(new_n1067), .B1(new_n813), .B2(new_n886), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1065), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1066), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1071), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1087), .A2(new_n1090), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1098), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1095), .A2(new_n1102), .A3(new_n1034), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1042), .B1(new_n734), .B2(new_n220), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n722), .A2(new_n572), .B1(new_n724), .B2(new_n787), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n781), .B(new_n384), .C1(new_n243), .C2(new_n710), .ZN(new_n1106));
  NOR3_X1   g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1107), .B1(new_n360), .B2(new_n707), .C1(new_n788), .C2(new_n714), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n711), .A2(G132), .B1(new_n775), .B2(G128), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1109), .B(new_n281), .C1(new_n266), .C2(new_n728), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G125), .B2(new_n725), .ZN(new_n1111));
  XOR2_X1   g0911(.A(KEYINPUT54), .B(G143), .Z(new_n1112));
  AOI22_X1  g0912(.A1(new_n982), .A2(new_n1112), .B1(G137), .B2(new_n708), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n719), .A2(G159), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n722), .A2(new_n253), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT53), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1111), .A2(new_n1113), .A3(new_n1114), .A4(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n770), .B1(new_n1108), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n793), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n751), .B1(new_n258), .B2(new_n1119), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1118), .B(new_n1120), .C1(new_n1082), .C2(new_n759), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1101), .A2(new_n1099), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1121), .B1(new_n1122), .B2(new_n964), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1103), .A2(new_n1123), .ZN(G378));
  NAND2_X1  g0924(.A1(new_n1095), .A2(new_n1065), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n875), .A2(G330), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n306), .A2(new_n348), .ZN(new_n1127));
  XOR2_X1   g0927(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1128));
  XOR2_X1   g0928(.A(new_n1127), .B(new_n1128), .Z(new_n1129));
  NAND2_X1  g0929(.A1(new_n275), .A2(new_n819), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1129), .B(new_n1131), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n883), .A2(new_n888), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1132), .B1(new_n883), .B2(new_n888), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1126), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1129), .B(new_n1130), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n889), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1063), .B1(new_n867), .B2(new_n874), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n883), .A2(new_n888), .A3(new_n1132), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1135), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1125), .A2(new_n1141), .A3(KEYINPUT57), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT57), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1065), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n1122), .B2(new_n1080), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1135), .A2(new_n1140), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1143), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1142), .A2(new_n1147), .A3(new_n1034), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1135), .A2(new_n1140), .A3(new_n964), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n751), .B1(G50), .B2(new_n1119), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n382), .ZN(new_n1151));
  AOI21_X1  g0951(.A(G50), .B1(new_n1151), .B2(new_n278), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n278), .B1(new_n724), .B2(new_n788), .C1(new_n710), .C2(new_n360), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n714), .A2(new_n243), .B1(new_n718), .B2(new_n216), .ZN(new_n1154));
  OR2_X1    g0954(.A1(new_n1154), .A2(KEYINPUT119), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(KEYINPUT119), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1013), .B(new_n1153), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n729), .A2(new_n257), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n384), .B1(new_n707), .B2(new_n220), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n579), .B2(new_n731), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1157), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT120), .Z(new_n1162));
  INV_X1    g0962(.A(KEYINPUT58), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1152), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT121), .Z(new_n1165));
  AOI22_X1  g0965(.A1(G128), .A2(new_n711), .B1(new_n731), .B2(G137), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n708), .A2(G132), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n723), .A2(new_n1112), .B1(new_n719), .B2(G150), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n775), .A2(G125), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1171), .A2(G33), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n729), .A2(new_n742), .ZN(new_n1174));
  AOI21_X1  g0974(.A(G41), .B1(new_n725), .B2(G124), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1165), .B(new_n1176), .C1(new_n1163), .C2(new_n1162), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1150), .B1(new_n1177), .B2(new_n699), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n1136), .B2(new_n760), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT122), .Z(new_n1180));
  AND2_X1   g0980(.A1(new_n1149), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1148), .A2(new_n1181), .ZN(G375));
  NAND4_X1  g0982(.A1(new_n1144), .A2(new_n1070), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1183), .A2(new_n962), .A3(new_n1098), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n885), .A2(new_n759), .ZN(new_n1185));
  INV_X1    g0985(.A(G128), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1158), .B1(new_n1186), .B2(new_n724), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n384), .B(new_n1187), .C1(G50), .C2(new_n719), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(new_n253), .B2(new_n701), .C1(new_n376), .C2(new_n722), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1189), .A2(KEYINPUT123), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1189), .A2(KEYINPUT123), .B1(G137), .B2(new_n711), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n775), .A2(G132), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n708), .A2(new_n1112), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1014), .B1(G97), .B2(new_n723), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n288), .B2(new_n728), .C1(new_n734), .C2(new_n360), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n384), .B1(new_n707), .B2(new_n243), .C1(new_n788), .C2(new_n710), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1198), .B1(new_n787), .B2(new_n714), .C1(new_n538), .C2(new_n724), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n770), .B1(new_n1194), .B2(new_n1199), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n752), .B(new_n1200), .C1(new_n216), .C2(new_n793), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1080), .A2(new_n964), .B1(new_n1185), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1184), .A2(new_n1202), .ZN(G381));
  AND2_X1   g1003(.A1(new_n1035), .A2(new_n1061), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n973), .A2(new_n1204), .A3(new_n996), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1205), .A2(G384), .A3(G381), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT124), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1103), .A2(new_n1207), .A3(new_n1123), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n1103), .B2(new_n1123), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(G375), .A2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(G393), .A2(G396), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1206), .A2(new_n1211), .A3(new_n1212), .ZN(G407));
  NAND2_X1  g1013(.A1(new_n1211), .A2(new_n630), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(G407), .A2(G213), .A3(new_n1214), .ZN(G409));
  NAND3_X1  g1015(.A1(new_n1148), .A2(G378), .A3(new_n1181), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1125), .A2(new_n1141), .A3(new_n962), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1181), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n630), .A2(G213), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT60), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1034), .B(new_n1098), .C1(new_n1183), .C2(new_n1222), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1183), .A2(new_n1222), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1202), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(G384), .ZN(new_n1226));
  AND4_X1   g1026(.A1(KEYINPUT62), .A2(new_n1220), .A3(new_n1221), .A4(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT125), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1220), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1216), .A2(new_n1219), .A3(KEYINPUT125), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1229), .A2(new_n1221), .A3(new_n1226), .A4(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT62), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1227), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT61), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n630), .A2(G213), .A3(G2897), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1226), .B(new_n1235), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1234), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n973), .A2(new_n1204), .A3(new_n996), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1204), .B1(new_n996), .B2(new_n973), .ZN(new_n1240));
  OAI21_X1  g1040(.A(KEYINPUT127), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n970), .A2(new_n908), .A3(new_n971), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n908), .B1(new_n970), .B2(new_n971), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n964), .B1(new_n961), .B2(new_n962), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n996), .ZN(new_n1246));
  OAI21_X1  g1046(.A(G390), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT127), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n1248), .A3(new_n1205), .ZN(new_n1249));
  XOR2_X1   g1049(.A(G393), .B(G396), .Z(new_n1250));
  AND3_X1   g1050(.A1(new_n1241), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1250), .B1(new_n1241), .B2(new_n1249), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n1233), .A2(new_n1238), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT63), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1231), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT126), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1231), .A2(KEYINPUT126), .A3(new_n1254), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1229), .A2(new_n1221), .A3(new_n1230), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1235), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1226), .B(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT61), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1250), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(new_n1239), .A2(new_n1240), .A3(KEYINPUT127), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1248), .B1(new_n1247), .B2(new_n1205), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1264), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1241), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1237), .A2(KEYINPUT63), .A3(new_n1226), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1263), .A2(new_n1267), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1253), .B1(new_n1259), .B2(new_n1270), .ZN(G405));
  OAI21_X1  g1071(.A(G375), .B1(new_n1209), .B2(new_n1208), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1272), .A2(new_n1216), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1226), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1273), .B(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1275), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1273), .B(new_n1226), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(new_n1268), .A3(new_n1267), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1278), .ZN(G402));
endmodule


