//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT64), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n465), .A2(new_n470), .ZN(G160));
  INV_X1    g046(.A(new_n461), .ZN(new_n472));
  INV_X1    g047(.A(new_n462), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n460), .B1(new_n472), .B2(new_n473), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  INV_X1    g056(.A(G138), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n483), .B1(new_n461), .B2(new_n462), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n483), .B(new_n486), .C1(new_n462), .C2(new_n461), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT65), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n491), .A2(new_n493), .A3(G2104), .ZN(new_n494));
  AND3_X1   g069(.A1(new_n489), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n490), .B1(new_n489), .B2(new_n494), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n488), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G88), .ZN(new_n506));
  INV_X1    g081(.A(G62), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n507), .B1(new_n501), .B2(new_n502), .ZN(new_n508));
  AND2_X1   g083(.A1(G75), .A2(G543), .ZN(new_n509));
  OAI21_X1  g084(.A(G651), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n500), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT66), .ZN(new_n514));
  AND3_X1   g089(.A1(new_n513), .A2(new_n514), .A3(G50), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n514), .B1(new_n513), .B2(G50), .ZN(new_n516));
  OAI211_X1 g091(.A(new_n506), .B(new_n510), .C1(new_n515), .C2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  INV_X1    g093(.A(G51), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n504), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT67), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT67), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n519), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n503), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n503), .A2(new_n504), .ZN(new_n528));
  INV_X1    g103(.A(G89), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n525), .B(new_n527), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n524), .A2(new_n530), .ZN(G168));
  INV_X1    g106(.A(KEYINPUT68), .ZN(new_n532));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n533), .B1(new_n521), .B2(new_n523), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G651), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n536), .A2(new_n537), .B1(new_n538), .B2(new_n528), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n532), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  NOR3_X1   g116(.A1(new_n534), .A2(new_n539), .A3(KEYINPUT68), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  INV_X1    g119(.A(new_n503), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  INV_X1    g121(.A(G68), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n545), .A2(new_n546), .B1(new_n547), .B2(new_n500), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(KEYINPUT69), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT69), .ZN(new_n550));
  OAI221_X1 g125(.A(new_n550), .B1(new_n547), .B2(new_n500), .C1(new_n545), .C2(new_n546), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n549), .A2(G651), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(G43), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n554), .B1(new_n521), .B2(new_n523), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n503), .A2(new_n504), .A3(G81), .ZN(new_n556));
  NOR3_X1   g131(.A1(new_n555), .A2(KEYINPUT70), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT70), .B1(new_n555), .B2(new_n556), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n553), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  NAND3_X1  g140(.A1(new_n504), .A2(G53), .A3(G543), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n566), .B(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n503), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G91), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n569), .A2(new_n537), .B1(new_n570), .B2(new_n528), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G299));
  INV_X1    g148(.A(G168), .ZN(G286));
  NAND2_X1  g149(.A1(new_n513), .A2(G49), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n503), .B2(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n503), .A2(new_n504), .A3(G87), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  INV_X1    g153(.A(G48), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT72), .B1(new_n520), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT72), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n513), .A2(new_n581), .A3(G48), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n580), .A2(new_n582), .B1(G86), .B2(new_n505), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n501), .B2(new_n502), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT71), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n589), .B1(new_n585), .B2(new_n586), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n583), .A2(new_n591), .ZN(G305));
  AND2_X1   g167(.A1(new_n503), .A2(G60), .ZN(new_n593));
  AND2_X1   g168(.A1(G72), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT73), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(G85), .B2(new_n505), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n595), .A2(new_n596), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n521), .A2(new_n523), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G47), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(G290));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NOR2_X1   g178(.A1(G301), .A2(new_n603), .ZN(new_n604));
  AND3_X1   g179(.A1(new_n521), .A2(KEYINPUT75), .A3(new_n523), .ZN(new_n605));
  AOI21_X1  g180(.A(KEYINPUT75), .B1(new_n521), .B2(new_n523), .ZN(new_n606));
  OAI21_X1  g181(.A(G54), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n503), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(new_n537), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  XOR2_X1   g185(.A(KEYINPUT74), .B(KEYINPUT10), .Z(new_n611));
  OR3_X1    g186(.A1(new_n528), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n528), .B2(new_n610), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n607), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n616), .A2(KEYINPUT76), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(KEYINPUT76), .ZN(new_n618));
  AND2_X1   g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n604), .B1(new_n619), .B2(new_n603), .ZN(G284));
  AOI21_X1  g195(.A(new_n604), .B1(new_n619), .B2(new_n603), .ZN(G321));
  NOR2_X1   g196(.A1(G286), .A2(new_n603), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n572), .B(KEYINPUT77), .Z(new_n623));
  AOI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(new_n603), .ZN(G297));
  AOI21_X1  g199(.A(new_n622), .B1(new_n623), .B2(new_n603), .ZN(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n619), .B1(new_n626), .B2(G860), .ZN(G148));
  NAND2_X1  g202(.A1(new_n619), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n560), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n474), .A2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n476), .A2(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n460), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT78), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2096), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT3), .B(G2104), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(new_n468), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n638), .A2(G2096), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n639), .A2(new_n644), .A3(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2427), .B(G2430), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(KEYINPUT14), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT79), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(new_n648), .B2(new_n649), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(G14), .B1(new_n658), .B2(new_n661), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(G401));
  INV_X1    g239(.A(KEYINPUT18), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2100), .ZN(new_n672));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n668), .B2(KEYINPUT18), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2096), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n672), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT80), .B(KEYINPUT20), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n679), .A2(new_n680), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n678), .A2(new_n681), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n678), .B2(new_n685), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1991), .B(G1996), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1981), .B(G1986), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT81), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n690), .B(new_n694), .ZN(G229));
  NOR2_X1   g270(.A1(G16), .A2(G24), .ZN(new_n696));
  XOR2_X1   g271(.A(G290), .B(KEYINPUT85), .Z(new_n697));
  AOI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(G16), .ZN(new_n698));
  INV_X1    g273(.A(G1986), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  MUX2_X1   g275(.A(G6), .B(G305), .S(G16), .Z(new_n701));
  XOR2_X1   g276(.A(KEYINPUT32), .B(G1981), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G22), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G166), .B2(new_n704), .ZN(new_n706));
  INV_X1    g281(.A(G1971), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n704), .A2(G23), .ZN(new_n709));
  INV_X1    g284(.A(G288), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n704), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT33), .B(G1976), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n703), .A2(new_n708), .A3(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT34), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n476), .A2(G119), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT82), .Z(new_n717));
  OAI21_X1  g292(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n718));
  INV_X1    g293(.A(G107), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(G2105), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n474), .B2(G131), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT83), .ZN(new_n723));
  MUX2_X1   g298(.A(G25), .B(new_n723), .S(G29), .Z(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT35), .B(G1991), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT84), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n724), .B(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n700), .A2(new_n715), .A3(new_n727), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT36), .Z(new_n729));
  NOR2_X1   g304(.A1(G4), .A2(G16), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT86), .Z(new_n731));
  INV_X1    g306(.A(new_n619), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(new_n704), .ZN(new_n733));
  INV_X1    g308(.A(G1348), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(G16), .A2(G19), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n560), .B2(G16), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(G1341), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(G1341), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n704), .A2(G20), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT23), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n572), .B2(new_n704), .ZN(new_n742));
  INV_X1    g317(.A(G1956), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G29), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G32), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT91), .B(KEYINPUT26), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n468), .A2(G105), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI22_X1  g326(.A1(G129), .A2(new_n476), .B1(new_n474), .B2(G141), .ZN(new_n752));
  AND3_X1   g327(.A1(new_n751), .A2(KEYINPUT92), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(KEYINPUT92), .B1(new_n751), .B2(new_n752), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n746), .B1(new_n755), .B2(new_n745), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT27), .B(G1996), .Z(new_n757));
  INV_X1    g332(.A(G2078), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n745), .A2(G27), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT94), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n497), .B2(G29), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n756), .A2(new_n757), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n738), .A2(new_n739), .A3(new_n744), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n474), .A2(G139), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT88), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT25), .Z(new_n767));
  AOI22_X1  g342(.A1(new_n640), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(new_n460), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n770), .A2(new_n745), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n745), .B2(G33), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(G2072), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT89), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n745), .A2(G35), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G162), .B2(new_n745), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT29), .Z(new_n778));
  INV_X1    g353(.A(G2090), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(KEYINPUT95), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n775), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G5), .A2(G16), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(KEYINPUT93), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n783), .A2(KEYINPUT93), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n784), .B(new_n785), .C1(G301), .C2(new_n704), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n780), .A2(KEYINPUT95), .B1(new_n787), .B2(G1961), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n778), .A2(new_n779), .ZN(new_n789));
  OAI22_X1  g364(.A1(new_n756), .A2(new_n757), .B1(new_n758), .B2(new_n761), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n745), .A2(G26), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT28), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n474), .A2(G140), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n476), .A2(G128), .ZN(new_n794));
  OR2_X1    g369(.A1(G104), .A2(G2105), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n795), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n792), .B1(new_n797), .B2(G29), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT87), .B(G2067), .Z(new_n799));
  OAI22_X1  g374(.A1(new_n638), .A2(new_n745), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g375(.A1(KEYINPUT24), .A2(G34), .ZN(new_n801));
  NOR2_X1   g376(.A1(KEYINPUT24), .A2(G34), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n745), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT90), .Z(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G160), .B2(G29), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G2084), .ZN(new_n806));
  NOR4_X1   g381(.A1(new_n789), .A2(new_n790), .A3(new_n800), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n773), .A2(G2072), .ZN(new_n808));
  NOR2_X1   g383(.A1(G168), .A2(new_n704), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n704), .B2(G21), .ZN(new_n810));
  INV_X1    g385(.A(G1966), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT30), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n813), .A2(G28), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n745), .B1(new_n813), .B2(G28), .ZN(new_n815));
  AND2_X1   g390(.A1(KEYINPUT31), .A2(G11), .ZN(new_n816));
  NOR2_X1   g391(.A1(KEYINPUT31), .A2(G11), .ZN(new_n817));
  OAI22_X1  g392(.A1(new_n814), .A2(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(new_n798), .B2(new_n799), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n810), .A2(new_n811), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n808), .A2(new_n812), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(G1961), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n821), .B1(new_n822), .B2(new_n786), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n782), .A2(new_n788), .A3(new_n807), .A4(new_n823), .ZN(new_n824));
  OR4_X1    g399(.A1(new_n729), .A2(new_n735), .A3(new_n763), .A4(new_n824), .ZN(G150));
  XNOR2_X1  g400(.A(G150), .B(KEYINPUT96), .ZN(G311));
  INV_X1    g401(.A(G55), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n521), .B2(new_n523), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n829));
  INV_X1    g404(.A(G93), .ZN(new_n830));
  OAI22_X1  g405(.A1(new_n829), .A2(new_n537), .B1(new_n830), .B2(new_n528), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n559), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n552), .B(new_n832), .C1(new_n833), .C2(new_n557), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n600), .A2(G55), .ZN(new_n835));
  NAND2_X1  g410(.A1(G80), .A2(G543), .ZN(new_n836));
  INV_X1    g411(.A(G67), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n545), .B2(new_n837), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n838), .A2(G651), .B1(new_n505), .B2(G93), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT97), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n835), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(KEYINPUT97), .B1(new_n828), .B2(new_n831), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n834), .B1(new_n560), .B2(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT38), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n619), .A2(G559), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n849), .A2(new_n850), .A3(G860), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n843), .A2(G860), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT98), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT37), .Z(new_n854));
  OR2_X1    g429(.A1(new_n851), .A2(new_n854), .ZN(G145));
  OAI21_X1  g430(.A(new_n797), .B1(new_n753), .B2(new_n754), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NOR3_X1   g432(.A1(new_n753), .A2(new_n754), .A3(new_n797), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n717), .B(new_n721), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n858), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n860), .A2(new_n722), .A3(new_n856), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n474), .A2(G142), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n476), .A2(G130), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n460), .A2(G118), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n863), .B(new_n864), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT100), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n642), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n862), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n487), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n486), .B1(new_n640), .B2(new_n483), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n489), .B(new_n494), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n859), .A2(new_n869), .A3(new_n861), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n871), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n874), .B1(new_n871), .B2(new_n875), .ZN(new_n877));
  OAI22_X1  g452(.A1(new_n876), .A2(new_n877), .B1(new_n765), .B2(new_n769), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n871), .A2(new_n875), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n489), .A2(new_n494), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n880), .B1(new_n485), .B2(new_n487), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n871), .A2(new_n874), .A3(new_n875), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n770), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n878), .A2(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(G160), .B(KEYINPUT99), .Z(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(G162), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n638), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(G37), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n878), .A2(new_n884), .A3(new_n888), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g468(.A1(new_n843), .A2(new_n603), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n628), .B(KEYINPUT101), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n845), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n616), .A2(G299), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n615), .A2(new_n898), .A3(new_n572), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n898), .B1(new_n615), .B2(new_n572), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT41), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n901), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT41), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n903), .A2(new_n904), .A3(new_n897), .A4(new_n899), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n896), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n900), .A2(new_n901), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n907), .B1(new_n896), .B2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(G290), .B(new_n710), .ZN(new_n910));
  XNOR2_X1  g485(.A(G305), .B(G166), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n910), .B(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT42), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n909), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n894), .B1(new_n914), .B2(new_n603), .ZN(G295));
  OAI21_X1  g490(.A(new_n894), .B1(new_n914), .B2(new_n603), .ZN(G331));
  OAI21_X1  g491(.A(new_n552), .B1(new_n833), .B2(new_n557), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n843), .ZN(new_n918));
  OAI21_X1  g493(.A(G286), .B1(new_n541), .B2(new_n542), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n535), .A2(new_n540), .A3(new_n532), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT68), .B1(new_n534), .B2(new_n539), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(G168), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n918), .A2(new_n923), .A3(new_n834), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n918), .A2(new_n923), .A3(KEYINPUT104), .A4(new_n834), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n919), .A2(new_n922), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n845), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n929), .B1(new_n845), .B2(new_n928), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n926), .B(new_n927), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n906), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n845), .A2(new_n928), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n935), .A3(new_n924), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n845), .A2(new_n928), .A3(KEYINPUT105), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n908), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n933), .A2(new_n939), .A3(new_n912), .ZN(new_n940));
  INV_X1    g515(.A(G37), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n938), .B1(new_n906), .B2(new_n932), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n943), .A2(new_n912), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT43), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g522(.A(KEYINPUT106), .B(KEYINPUT43), .C1(new_n942), .C2(new_n944), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n936), .A2(new_n937), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n902), .A2(new_n905), .ZN(new_n950));
  OAI22_X1  g525(.A1(new_n932), .A2(new_n908), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n912), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT107), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(G37), .B1(new_n943), .B2(new_n912), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n951), .A2(KEYINPUT107), .A3(new_n952), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n955), .A2(new_n956), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n947), .A2(new_n948), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n957), .B1(new_n942), .B2(new_n944), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n961), .B1(new_n962), .B2(new_n957), .ZN(new_n963));
  MUX2_X1   g538(.A(new_n960), .B(new_n963), .S(KEYINPUT44), .Z(G397));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n497), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT50), .ZN(new_n967));
  NAND2_X1  g542(.A1(G160), .A2(G40), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n489), .A2(new_n494), .ZN(new_n969));
  AOI21_X1  g544(.A(G1384), .B1(new_n488), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(G1348), .B1(new_n967), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G2067), .ZN(new_n974));
  INV_X1    g549(.A(G40), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n465), .A2(new_n470), .A3(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n970), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT114), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n970), .A2(new_n979), .A3(new_n976), .A4(new_n974), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT115), .B1(new_n973), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n874), .A2(new_n971), .A3(new_n965), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n976), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n971), .B1(new_n497), .B2(new_n965), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n734), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT115), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n986), .A2(new_n987), .A3(new_n978), .A4(new_n980), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n982), .A2(new_n616), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT116), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n982), .A2(new_n988), .A3(new_n991), .A4(new_n616), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n993), .B(KEYINPUT57), .C1(new_n568), .C2(new_n571), .ZN(new_n994));
  INV_X1    g569(.A(new_n571), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n566), .B(KEYINPUT9), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n993), .A2(KEYINPUT57), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n993), .A2(KEYINPUT57), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n995), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n994), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n497), .A2(new_n971), .A3(new_n965), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT50), .B1(new_n881), .B2(G1384), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n976), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n743), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n966), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n968), .B1(new_n970), .B2(KEYINPUT45), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT56), .B(G2072), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1000), .B1(new_n1004), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n990), .A2(new_n992), .A3(new_n1011), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n1004), .A2(new_n1009), .A3(new_n1000), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n982), .A2(new_n988), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(KEYINPUT60), .A3(new_n615), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1004), .A2(new_n1009), .A3(new_n1000), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1011), .A2(KEYINPUT61), .A3(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n874), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n976), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT45), .B1(new_n497), .B2(new_n965), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1019), .A2(new_n1020), .A3(G1996), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT58), .B(G1341), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1022), .B1(new_n970), .B2(new_n976), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n560), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT59), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(KEYINPUT117), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  OAI221_X1 g602(.A(new_n560), .B1(KEYINPUT117), .B2(new_n1025), .C1(new_n1021), .C2(new_n1023), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT61), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n1013), .B2(new_n1010), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1015), .A2(new_n1017), .A3(new_n1029), .A4(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT60), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n982), .A2(new_n1033), .A3(new_n988), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1033), .B1(new_n982), .B2(new_n988), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1034), .A2(new_n1035), .A3(new_n615), .ZN(new_n1036));
  OAI22_X1  g611(.A1(new_n1012), .A2(new_n1013), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT49), .ZN(new_n1038));
  INV_X1    g613(.A(G1981), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n583), .A2(new_n1039), .A3(new_n591), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1039), .B1(new_n583), .B2(new_n591), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1038), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G305), .A2(G1981), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(KEYINPUT49), .A3(new_n1040), .ZN(new_n1045));
  INV_X1    g620(.A(G8), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1046), .B1(new_n970), .B2(new_n976), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n710), .A2(G1976), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1049), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1052));
  INV_X1    g627(.A(G1976), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(G288), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1051), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n707), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1001), .A2(new_n779), .A3(new_n1002), .A4(new_n976), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1046), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g633(.A(KEYINPUT110), .B(KEYINPUT55), .Z(new_n1059));
  AND3_X1   g634(.A1(G303), .A2(G8), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT110), .ZN(new_n1061));
  AOI22_X1  g636(.A1(G303), .A2(G8), .B1(new_n1061), .B2(KEYINPUT55), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1048), .B(new_n1055), .C1(new_n1058), .C2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n967), .A2(new_n972), .A3(new_n779), .ZN(new_n1066));
  AOI211_X1 g641(.A(new_n1046), .B(new_n1063), .C1(new_n1056), .C2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1005), .B1(new_n881), .B2(G1384), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(G2078), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1069), .A2(new_n1018), .A3(new_n976), .A4(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n822), .B1(new_n984), .B2(new_n985), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1019), .A2(new_n1020), .A3(G2078), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1072), .B(new_n1073), .C1(new_n1074), .C2(KEYINPUT53), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(G171), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1006), .A2(new_n1007), .A3(new_n758), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n1070), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT45), .B1(new_n874), .B2(new_n965), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT111), .B1(new_n1079), .B2(new_n968), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT111), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1069), .A2(new_n1082), .A3(new_n976), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1080), .A2(new_n1081), .A3(new_n1083), .A4(new_n1071), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1078), .A2(new_n1084), .A3(G301), .A4(new_n1073), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1076), .A2(KEYINPUT54), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1068), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1078), .A2(new_n1084), .A3(new_n1073), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G171), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1089), .A2(KEYINPUT121), .A3(G171), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1075), .A2(G171), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1087), .B1(new_n1088), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1037), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1080), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n811), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n984), .A2(new_n985), .ZN(new_n1102));
  INV_X1    g677(.A(G2084), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1046), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(G168), .A2(new_n1046), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1105), .A2(KEYINPUT51), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1106), .B(KEYINPUT119), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1101), .A2(KEYINPUT118), .A3(new_n1104), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1110), .B1(new_n1115), .B2(G8), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT51), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1108), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1115), .A2(new_n1106), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1099), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n984), .A2(new_n985), .A3(G2084), .ZN(new_n1121));
  AOI211_X1 g696(.A(new_n1112), .B(new_n1121), .C1(new_n811), .C2(new_n1100), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT118), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1123));
  OAI21_X1  g698(.A(G8), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1117), .B1(new_n1124), .B2(new_n1109), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1099), .B(new_n1119), .C1(new_n1125), .C2(new_n1107), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1098), .B1(new_n1120), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(G288), .A2(G1976), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1041), .B1(new_n1048), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1048), .A2(new_n1055), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1131), .A2(new_n1047), .B1(new_n1132), .B2(new_n1067), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1105), .A2(G168), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1046), .B1(new_n1066), .B2(new_n1056), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n1064), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1135), .A2(KEYINPUT63), .A3(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1132), .B1(new_n1136), .B2(new_n1064), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n1139), .A2(KEYINPUT112), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(KEYINPUT112), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1138), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT63), .B1(new_n1135), .B2(new_n1068), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1133), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1128), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT62), .B1(new_n1120), .B2(new_n1127), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1119), .B1(new_n1125), .B2(new_n1107), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT120), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1150), .A2(new_n1151), .A3(new_n1126), .ZN(new_n1152));
  AOI211_X1 g727(.A(new_n1067), .B(new_n1065), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1148), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1097), .B1(new_n1150), .B2(new_n1126), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT122), .B1(new_n1155), .B2(new_n1144), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1147), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n755), .B(G1996), .ZN(new_n1158));
  XOR2_X1   g733(.A(new_n722), .B(new_n725), .Z(new_n1159));
  XNOR2_X1  g734(.A(new_n797), .B(new_n974), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1069), .A2(new_n968), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n1162), .A2(KEYINPUT108), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(KEYINPUT108), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(G290), .A2(G1986), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT109), .ZN(new_n1169));
  NOR2_X1   g744(.A1(G290), .A2(G1986), .ZN(new_n1170));
  OR3_X1    g745(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1165), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1172), .B1(new_n1169), .B2(new_n1168), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1166), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1157), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(G1996), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1165), .A2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT46), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n755), .A2(new_n1160), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1178), .B1(new_n1172), .B2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1180), .B(KEYINPUT47), .ZN(new_n1181));
  OR2_X1    g756(.A1(new_n1181), .A2(KEYINPUT123), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(KEYINPUT123), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n723), .A2(new_n725), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1184), .A2(new_n1160), .A3(new_n1158), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n797), .A2(G2067), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1172), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(KEYINPUT48), .B1(new_n1165), .B2(new_n1170), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1166), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1165), .A2(KEYINPUT48), .A3(new_n1170), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1187), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  AND3_X1   g766(.A1(new_n1182), .A2(new_n1183), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1175), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT124), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1175), .A2(KEYINPUT124), .A3(new_n1192), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1195), .A2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g772(.A(KEYINPUT125), .ZN(new_n1199));
  NOR3_X1   g773(.A1(G229), .A2(new_n458), .A3(G227), .ZN(new_n1200));
  OAI21_X1  g774(.A(new_n1200), .B1(new_n662), .B2(new_n663), .ZN(new_n1201));
  AOI21_X1  g775(.A(new_n1201), .B1(new_n890), .B2(new_n891), .ZN(new_n1202));
  AND3_X1   g776(.A1(new_n960), .A2(new_n1199), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g777(.A(new_n1199), .B1(new_n960), .B2(new_n1202), .ZN(new_n1204));
  INV_X1    g778(.A(KEYINPUT126), .ZN(new_n1205));
  NOR3_X1   g779(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g780(.A1(new_n933), .A2(new_n939), .ZN(new_n1207));
  NAND2_X1  g781(.A1(new_n1207), .A2(new_n952), .ZN(new_n1208));
  AOI21_X1  g782(.A(new_n957), .B1(new_n956), .B2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g783(.A(new_n959), .B1(new_n1209), .B2(KEYINPUT106), .ZN(new_n1210));
  INV_X1    g784(.A(new_n948), .ZN(new_n1211));
  OAI21_X1  g785(.A(new_n1202), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g786(.A1(new_n1212), .A2(KEYINPUT125), .ZN(new_n1213));
  NAND3_X1  g787(.A1(new_n960), .A2(new_n1199), .A3(new_n1202), .ZN(new_n1214));
  AOI21_X1  g788(.A(KEYINPUT126), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g789(.A1(new_n1206), .A2(new_n1215), .ZN(G308));
  NAND2_X1  g790(.A1(new_n1213), .A2(new_n1214), .ZN(G225));
endmodule


