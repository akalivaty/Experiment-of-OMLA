

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878;

  BUF_X1 U373 ( .A(n804), .Z(n351) );
  NAND2_X1 U374 ( .A1(n355), .A2(n426), .ZN(n421) );
  AND2_X1 U375 ( .A1(n427), .A2(n369), .ZN(n355) );
  BUF_X1 U376 ( .A(n669), .Z(n657) );
  OR2_X1 U377 ( .A1(n798), .A2(n352), .ZN(n704) );
  OR2_X1 U378 ( .A1(n615), .A2(n616), .ZN(n679) );
  XNOR2_X1 U379 ( .A(n617), .B(KEYINPUT97), .ZN(n868) );
  BUF_X1 U380 ( .A(G143), .Z(n350) );
  XNOR2_X1 U381 ( .A(n549), .B(n548), .ZN(n617) );
  XNOR2_X1 U382 ( .A(n484), .B(G131), .ZN(n549) );
  XNOR2_X1 U383 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n484) );
  AND2_X2 U384 ( .A1(n501), .A2(n482), .ZN(n365) );
  NAND2_X2 U385 ( .A1(n808), .A2(n667), .ZN(n736) );
  AND2_X2 U386 ( .A1(n400), .A2(n399), .ZN(n398) );
  NAND2_X2 U387 ( .A1(n713), .A2(n497), .ZN(n496) );
  XNOR2_X2 U388 ( .A(n682), .B(n681), .ZN(n703) );
  OR2_X1 U389 ( .A1(n376), .A2(n758), .ZN(n498) );
  NOR2_X1 U390 ( .A1(G953), .A2(G237), .ZN(n544) );
  NAND2_X1 U391 ( .A1(n693), .A2(n819), .ZN(n822) );
  INV_X1 U392 ( .A(G953), .ZN(n870) );
  AND2_X1 U393 ( .A1(n414), .A2(n643), .ZN(n352) );
  AND2_X2 U394 ( .A1(n406), .A2(n405), .ZN(n404) );
  OR2_X2 U395 ( .A1(n669), .A2(n822), .ZN(n696) );
  XNOR2_X2 U396 ( .A(n436), .B(n639), .ZN(n645) );
  XNOR2_X1 U397 ( .A(n739), .B(n738), .ZN(n807) );
  NOR2_X1 U398 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U399 ( .A1(n473), .A2(n470), .ZN(n700) );
  NAND2_X1 U400 ( .A1(n740), .A2(n807), .ZN(n742) );
  NOR2_X1 U401 ( .A1(n726), .A2(n725), .ZN(n380) );
  AND2_X1 U402 ( .A1(n506), .A2(n488), .ZN(n411) );
  AND2_X1 U403 ( .A1(n425), .A2(n424), .ZN(n423) );
  XNOR2_X1 U404 ( .A(n692), .B(n370), .ZN(n376) );
  XNOR2_X1 U405 ( .A(n642), .B(KEYINPUT39), .ZN(n660) );
  XNOR2_X1 U406 ( .A(n456), .B(KEYINPUT22), .ZN(n707) );
  INV_X1 U407 ( .A(n474), .ZN(n473) );
  XNOR2_X1 U408 ( .A(n520), .B(n491), .ZN(n644) );
  OR2_X1 U409 ( .A1(n799), .A2(n783), .ZN(n705) );
  XNOR2_X1 U410 ( .A(n580), .B(n551), .ZN(n428) );
  INV_X1 U411 ( .A(n404), .ZN(n383) );
  INV_X1 U412 ( .A(n758), .ZN(n499) );
  XNOR2_X1 U413 ( .A(n478), .B(KEYINPUT89), .ZN(n635) );
  NOR2_X1 U414 ( .A1(n762), .A2(n357), .ZN(n478) );
  INV_X1 U415 ( .A(n468), .ZN(n467) );
  INV_X1 U416 ( .A(G469), .ZN(n619) );
  XNOR2_X1 U417 ( .A(n517), .B(n516), .ZN(n519) );
  NOR2_X1 U418 ( .A1(n393), .A2(n376), .ZN(n493) );
  NAND2_X1 U419 ( .A1(n499), .A2(n394), .ZN(n393) );
  NOR2_X1 U420 ( .A1(n490), .A2(n489), .ZN(n458) );
  AND2_X1 U421 ( .A1(n635), .A2(n637), .ZN(n489) );
  NOR2_X1 U422 ( .A1(n465), .A2(n464), .ZN(n463) );
  NOR2_X1 U423 ( .A1(n834), .A2(n469), .ZN(n464) );
  AND2_X1 U424 ( .A1(n428), .A2(n460), .ZN(n465) );
  NOR2_X1 U425 ( .A1(n468), .A2(n472), .ZN(n460) );
  INV_X1 U426 ( .A(G237), .ZN(n592) );
  NAND2_X1 U427 ( .A1(G902), .A2(G472), .ZN(n475) );
  OR2_X1 U428 ( .A1(n428), .A2(n477), .ZN(n476) );
  XOR2_X1 U429 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n522) );
  XNOR2_X1 U430 ( .A(G116), .B(G122), .ZN(n521) );
  XNOR2_X1 U431 ( .A(G134), .B(G107), .ZN(n524) );
  XNOR2_X1 U432 ( .A(n700), .B(n654), .ZN(n686) );
  NOR2_X1 U433 ( .A1(n693), .A2(n625), .ZN(n576) );
  XNOR2_X1 U434 ( .A(G137), .B(G134), .ZN(n548) );
  XNOR2_X1 U435 ( .A(G119), .B(KEYINPUT3), .ZN(n542) );
  XNOR2_X1 U436 ( .A(n558), .B(n559), .ZN(n749) );
  NAND2_X1 U437 ( .A1(G234), .A2(G237), .ZN(n567) );
  NAND2_X1 U438 ( .A1(n649), .A2(n407), .ZN(n405) );
  NAND2_X1 U439 ( .A1(n403), .A2(n402), .ZN(n401) );
  NOR2_X1 U440 ( .A1(n649), .A2(n407), .ZN(n402) );
  XNOR2_X1 U441 ( .A(n629), .B(KEYINPUT80), .ZN(n641) );
  NOR2_X1 U442 ( .A1(n626), .A2(n625), .ZN(n628) );
  NOR2_X2 U443 ( .A1(n685), .A2(n684), .ZN(n456) );
  XOR2_X1 U444 ( .A(n749), .B(KEYINPUT123), .Z(n750) );
  XNOR2_X1 U445 ( .A(n533), .B(n412), .ZN(n768) );
  XNOR2_X1 U446 ( .A(n527), .B(n413), .ZN(n412) );
  INV_X1 U447 ( .A(KEYINPUT104), .ZN(n413) );
  XNOR2_X1 U448 ( .A(n753), .B(n754), .ZN(n755) );
  XNOR2_X1 U449 ( .A(n631), .B(n744), .ZN(n745) );
  AND2_X1 U450 ( .A1(n390), .A2(n408), .ZN(n389) );
  INV_X1 U451 ( .A(KEYINPUT44), .ZN(n394) );
  NAND2_X1 U452 ( .A1(n397), .A2(n396), .ZN(n395) );
  NOR2_X1 U453 ( .A1(n384), .A2(n383), .ZN(n396) );
  INV_X1 U454 ( .A(KEYINPUT30), .ZN(n469) );
  NAND2_X1 U455 ( .A1(n834), .A2(n469), .ZN(n468) );
  AND2_X1 U456 ( .A1(n354), .A2(n446), .ZN(n440) );
  NOR2_X1 U457 ( .A1(n836), .A2(n356), .ZN(n482) );
  NAND2_X1 U458 ( .A1(G953), .A2(G902), .ZN(n673) );
  XOR2_X1 U459 ( .A(G125), .B(G140), .Z(n518) );
  XNOR2_X1 U460 ( .A(KEYINPUT4), .B(G146), .ZN(n539) );
  XOR2_X1 U461 ( .A(G119), .B(KEYINPUT23), .Z(n554) );
  XOR2_X1 U462 ( .A(KEYINPUT8), .B(n528), .Z(n552) );
  NAND2_X1 U463 ( .A1(n870), .A2(G234), .ZN(n528) );
  XNOR2_X1 U464 ( .A(G113), .B(G122), .ZN(n508) );
  XNOR2_X1 U465 ( .A(G125), .B(KEYINPUT84), .ZN(n585) );
  XOR2_X1 U466 ( .A(KEYINPUT17), .B(KEYINPUT83), .Z(n586) );
  INV_X1 U467 ( .A(KEYINPUT48), .ZN(n659) );
  OR2_X1 U468 ( .A1(n645), .A2(n502), .ZN(n483) );
  NAND2_X1 U469 ( .A1(n834), .A2(KEYINPUT111), .ZN(n502) );
  NAND2_X1 U470 ( .A1(n645), .A2(n646), .ZN(n501) );
  INV_X1 U471 ( .A(n647), .ZN(n479) );
  INV_X1 U472 ( .A(KEYINPUT42), .ZN(n407) );
  INV_X1 U473 ( .A(n700), .ZN(n824) );
  AND2_X1 U474 ( .A1(n466), .A2(n463), .ZN(n462) );
  XNOR2_X1 U475 ( .A(n656), .B(KEYINPUT1), .ZN(n669) );
  INV_X1 U476 ( .A(KEYINPUT5), .ZN(n545) );
  BUF_X1 U477 ( .A(n808), .Z(n869) );
  INV_X1 U478 ( .A(G104), .ZN(n577) );
  XNOR2_X1 U479 ( .A(G110), .B(G107), .ZN(n578) );
  XNOR2_X1 U480 ( .A(KEYINPUT16), .B(G122), .ZN(n582) );
  XNOR2_X1 U481 ( .A(n524), .B(n523), .ZN(n525) );
  INV_X1 U482 ( .A(KEYINPUT102), .ZN(n523) );
  XNOR2_X1 U483 ( .A(n868), .B(n358), .ZN(n500) );
  INV_X1 U484 ( .A(KEYINPUT40), .ZN(n409) );
  AND2_X1 U485 ( .A1(n686), .A2(n834), .ZN(n373) );
  NAND2_X1 U486 ( .A1(n420), .A2(n448), .ZN(n426) );
  INV_X1 U487 ( .A(KEYINPUT35), .ZN(n422) );
  AND2_X1 U488 ( .A1(n417), .A2(KEYINPUT35), .ZN(n416) );
  NAND2_X1 U489 ( .A1(n419), .A2(n353), .ZN(n418) );
  AND2_X1 U490 ( .A1(n689), .A2(n392), .ZN(n690) );
  INV_X1 U491 ( .A(n651), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n492), .B(G475), .ZN(n491) );
  INV_X1 U493 ( .A(KEYINPUT13), .ZN(n492) );
  XNOR2_X1 U494 ( .A(n535), .B(n534), .ZN(n643) );
  NAND2_X1 U495 ( .A1(n747), .A2(G953), .ZN(n770) );
  NOR2_X1 U496 ( .A1(n641), .A2(n634), .ZN(n762) );
  NAND2_X1 U497 ( .A1(n435), .A2(n361), .ZN(n634) );
  NAND2_X1 U498 ( .A1(n630), .A2(n644), .ZN(n787) );
  INV_X1 U499 ( .A(KEYINPUT124), .ZN(n450) );
  XNOR2_X1 U500 ( .A(n769), .B(n459), .ZN(n771) );
  INV_X1 U501 ( .A(n768), .ZN(n459) );
  INV_X1 U502 ( .A(KEYINPUT60), .ZN(n454) );
  INV_X1 U503 ( .A(KEYINPUT56), .ZN(n452) );
  INV_X1 U504 ( .A(G137), .ZN(n391) );
  INV_X1 U505 ( .A(G131), .ZN(n386) );
  XNOR2_X1 U506 ( .A(n506), .B(n374), .ZN(n802) );
  INV_X1 U507 ( .A(G125), .ZN(n374) );
  INV_X1 U508 ( .A(G119), .ZN(n372) );
  AND2_X1 U509 ( .A1(n447), .A2(n361), .ZN(n353) );
  AND2_X1 U510 ( .A1(n445), .A2(n716), .ZN(n354) );
  AND2_X1 U511 ( .A1(n503), .A2(n646), .ZN(n356) );
  AND2_X1 U512 ( .A1(n838), .A2(KEYINPUT47), .ZN(n357) );
  XOR2_X1 U513 ( .A(n618), .B(G140), .Z(n358) );
  XOR2_X1 U514 ( .A(KEYINPUT24), .B(G110), .Z(n359) );
  AND2_X1 U515 ( .A1(n470), .A2(KEYINPUT30), .ZN(n360) );
  AND2_X1 U516 ( .A1(n414), .A2(n630), .ZN(n361) );
  NAND2_X1 U517 ( .A1(n614), .A2(n728), .ZN(n362) );
  AND2_X1 U518 ( .A1(n808), .A2(KEYINPUT2), .ZN(n363) );
  AND2_X1 U519 ( .A1(n501), .A2(n429), .ZN(n364) );
  AND2_X1 U520 ( .A1(n448), .A2(KEYINPUT35), .ZN(n366) );
  INV_X1 U521 ( .A(n472), .ZN(n471) );
  NAND2_X1 U522 ( .A1(n593), .A2(n477), .ZN(n472) );
  INV_X1 U523 ( .A(G902), .ZN(n593) );
  OR2_X1 U524 ( .A1(n652), .A2(n409), .ZN(n367) );
  NOR2_X1 U525 ( .A1(n803), .A2(n759), .ZN(n368) );
  AND2_X1 U526 ( .A1(n353), .A2(n422), .ZN(n369) );
  XNOR2_X1 U527 ( .A(n691), .B(KEYINPUT68), .ZN(n370) );
  INV_X1 U528 ( .A(KEYINPUT111), .ZN(n646) );
  INV_X1 U529 ( .A(KEYINPUT34), .ZN(n449) );
  INV_X1 U530 ( .A(KEYINPUT46), .ZN(n410) );
  XNOR2_X1 U531 ( .A(n376), .B(n372), .ZN(G21) );
  NAND2_X1 U532 ( .A1(n653), .A2(n373), .ZN(n661) );
  NAND2_X1 U533 ( .A1(n658), .A2(n392), .ZN(n506) );
  NAND2_X1 U534 ( .A1(n382), .A2(n375), .ZN(n379) );
  NAND2_X2 U535 ( .A1(n439), .A2(n441), .ZN(n375) );
  INV_X1 U536 ( .A(n375), .ZN(n811) );
  NAND2_X1 U537 ( .A1(n363), .A2(n375), .ZN(n739) );
  NOR2_X2 U538 ( .A1(n378), .A2(n377), .ZN(n381) );
  AND2_X2 U539 ( .A1(n717), .A2(n811), .ZN(n377) );
  NAND2_X1 U540 ( .A1(n380), .A2(n379), .ZN(n378) );
  NAND2_X1 U541 ( .A1(n381), .A2(n737), .ZN(n740) );
  NAND2_X1 U542 ( .A1(n734), .A2(n733), .ZN(n382) );
  NAND2_X1 U543 ( .A1(n401), .A2(KEYINPUT46), .ZN(n384) );
  NAND2_X2 U544 ( .A1(n404), .A2(n401), .ZN(n385) );
  NAND2_X1 U545 ( .A1(n385), .A2(n410), .ZN(n399) );
  XNOR2_X1 U546 ( .A(n385), .B(n391), .ZN(G39) );
  INV_X1 U547 ( .A(n387), .ZN(n397) );
  NAND2_X1 U548 ( .A1(n387), .A2(n410), .ZN(n400) );
  XNOR2_X1 U549 ( .A(n387), .B(n386), .ZN(G33) );
  NAND2_X2 U550 ( .A1(n389), .A2(n388), .ZN(n387) );
  OR2_X1 U551 ( .A1(n660), .A2(n367), .ZN(n388) );
  NAND2_X1 U552 ( .A1(n660), .A2(n409), .ZN(n390) );
  XNOR2_X1 U553 ( .A(n657), .B(KEYINPUT95), .ZN(n392) );
  NAND2_X1 U554 ( .A1(n398), .A2(n395), .ZN(n650) );
  INV_X1 U555 ( .A(n805), .ZN(n403) );
  NAND2_X1 U556 ( .A1(n805), .A2(n407), .ZN(n406) );
  NAND2_X1 U557 ( .A1(n652), .A2(n409), .ZN(n408) );
  NAND2_X1 U558 ( .A1(n411), .A2(n485), .ZN(n490) );
  INV_X1 U559 ( .A(n643), .ZN(n630) );
  INV_X1 U560 ( .A(n644), .ZN(n414) );
  NAND2_X1 U561 ( .A1(n415), .A2(n793), .ZN(n622) );
  XNOR2_X1 U562 ( .A(n538), .B(n537), .ZN(n415) );
  NAND2_X2 U563 ( .A1(n432), .A2(n431), .ZN(n805) );
  NAND2_X1 U564 ( .A1(n804), .A2(KEYINPUT34), .ZN(n427) );
  NAND2_X1 U565 ( .A1(n418), .A2(n416), .ZN(n424) );
  NAND2_X1 U566 ( .A1(n353), .A2(n449), .ZN(n417) );
  INV_X1 U567 ( .A(n804), .ZN(n419) );
  NAND2_X1 U568 ( .A1(n420), .A2(n366), .ZN(n425) );
  INV_X1 U569 ( .A(n804), .ZN(n420) );
  NAND2_X2 U570 ( .A1(n423), .A2(n421), .ZN(n761) );
  NAND2_X1 U571 ( .A1(n428), .A2(n471), .ZN(n470) );
  XNOR2_X1 U572 ( .A(n428), .B(KEYINPUT62), .ZN(n763) );
  NAND2_X1 U573 ( .A1(n364), .A2(n483), .ZN(n431) );
  AND2_X1 U574 ( .A1(n482), .A2(n647), .ZN(n429) );
  NAND2_X1 U575 ( .A1(n430), .A2(n479), .ZN(n432) );
  NAND2_X1 U576 ( .A1(n365), .A2(n483), .ZN(n430) );
  XNOR2_X1 U577 ( .A(n433), .B(n500), .ZN(n773) );
  XNOR2_X2 U578 ( .A(n433), .B(n591), .ZN(n631) );
  XNOR2_X2 U579 ( .A(n580), .B(n579), .ZN(n433) );
  XNOR2_X1 U580 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U581 ( .A(n557), .B(n556), .ZN(n558) );
  NAND2_X1 U582 ( .A1(n438), .A2(n700), .ZN(n437) );
  XNOR2_X1 U583 ( .A(n437), .B(KEYINPUT28), .ZN(n648) );
  NAND2_X1 U584 ( .A1(n650), .A2(n458), .ZN(n505) );
  NAND2_X1 U585 ( .A1(n476), .A2(n475), .ZN(n474) );
  NAND2_X1 U586 ( .A1(n474), .A2(n467), .ZN(n466) );
  NOR2_X1 U587 ( .A1(n656), .A2(n822), .ZN(n627) );
  AND2_X1 U588 ( .A1(n701), .A2(n434), .ZN(n702) );
  AND2_X1 U589 ( .A1(n621), .A2(n434), .ZN(n793) );
  INV_X1 U590 ( .A(n656), .ZN(n434) );
  INV_X1 U591 ( .A(n436), .ZN(n435) );
  NOR2_X1 U592 ( .A1(n661), .A2(n436), .ZN(n655) );
  AND2_X1 U593 ( .A1(n436), .A2(n666), .ZN(n759) );
  XNOR2_X2 U594 ( .A(n633), .B(n632), .ZN(n436) );
  NAND2_X1 U595 ( .A1(n495), .A2(n440), .ZN(n439) );
  AND2_X2 U596 ( .A1(n444), .A2(n442), .ZN(n441) );
  NAND2_X1 U597 ( .A1(n443), .A2(n457), .ZN(n442) );
  NAND2_X1 U598 ( .A1(n446), .A2(n445), .ZN(n443) );
  NAND2_X1 U599 ( .A1(n496), .A2(n457), .ZN(n444) );
  NAND2_X1 U600 ( .A1(n761), .A2(KEYINPUT44), .ZN(n445) );
  NAND2_X1 U601 ( .A1(n494), .A2(n493), .ZN(n446) );
  NAND2_X1 U602 ( .A1(n685), .A2(KEYINPUT34), .ZN(n447) );
  NOR2_X1 U603 ( .A1(n685), .A2(KEYINPUT34), .ZN(n448) );
  XNOR2_X2 U604 ( .A(n672), .B(n671), .ZN(n804) );
  XNOR2_X1 U605 ( .A(n451), .B(n450), .ZN(G66) );
  NAND2_X1 U606 ( .A1(n752), .A2(n770), .ZN(n451) );
  XNOR2_X1 U607 ( .A(n453), .B(n452), .ZN(G51) );
  NAND2_X1 U608 ( .A1(n748), .A2(n770), .ZN(n453) );
  XNOR2_X1 U609 ( .A(n455), .B(n454), .ZN(G60) );
  NAND2_X1 U610 ( .A1(n757), .A2(n770), .ZN(n455) );
  XNOR2_X2 U611 ( .A(n698), .B(n697), .ZN(n830) );
  INV_X1 U612 ( .A(n716), .ZN(n457) );
  OR2_X2 U613 ( .A1(n773), .A2(G902), .ZN(n620) );
  AND2_X2 U614 ( .A1(n504), .A2(n368), .ZN(n808) );
  NAND2_X1 U615 ( .A1(n462), .A2(n461), .ZN(n626) );
  NAND2_X1 U616 ( .A1(n473), .A2(n360), .ZN(n461) );
  INV_X1 U617 ( .A(G472), .ZN(n477) );
  NAND2_X1 U618 ( .A1(n480), .A2(n483), .ZN(n837) );
  NOR2_X1 U619 ( .A1(n481), .A2(n356), .ZN(n480) );
  INV_X1 U620 ( .A(n501), .ZN(n481) );
  XNOR2_X1 U621 ( .A(n505), .B(n659), .ZN(n504) );
  INV_X1 U622 ( .A(n496), .ZN(n495) );
  OR2_X2 U623 ( .A1(n711), .A2(n710), .ZN(n760) );
  NAND2_X1 U624 ( .A1(n808), .A2(n729), .ZN(n734) );
  NOR2_X1 U625 ( .A1(n808), .A2(n719), .ZN(n726) );
  NAND2_X1 U626 ( .A1(n487), .A2(n486), .ZN(n485) );
  NOR2_X1 U627 ( .A1(n635), .A2(n637), .ZN(n486) );
  INV_X1 U628 ( .A(n636), .ZN(n487) );
  NAND2_X1 U629 ( .A1(n636), .A2(n637), .ZN(n488) );
  INV_X1 U630 ( .A(n761), .ZN(n494) );
  NAND2_X1 U631 ( .A1(n498), .A2(KEYINPUT44), .ZN(n497) );
  XNOR2_X2 U632 ( .A(n866), .B(n541), .ZN(n580) );
  XNOR2_X2 U633 ( .A(n540), .B(n539), .ZN(n866) );
  INV_X1 U634 ( .A(n640), .ZN(n833) );
  INV_X1 U635 ( .A(n834), .ZN(n503) );
  BUF_X1 U636 ( .A(n767), .Z(n772) );
  XNOR2_X2 U637 ( .A(n742), .B(n741), .ZN(n767) );
  NOR2_X1 U638 ( .A1(n842), .A2(n351), .ZN(n507) );
  INV_X1 U639 ( .A(KEYINPUT77), .ZN(n537) );
  INV_X1 U640 ( .A(KEYINPUT75), .ZN(n637) );
  XNOR2_X1 U641 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U642 ( .A(n549), .B(n515), .ZN(n516) );
  XNOR2_X1 U643 ( .A(n584), .B(n547), .ZN(n550) );
  XNOR2_X1 U644 ( .A(n526), .B(n525), .ZN(n527) );
  BUF_X1 U645 ( .A(n773), .Z(n776) );
  INV_X1 U646 ( .A(KEYINPUT47), .ZN(n536) );
  XOR2_X1 U647 ( .A(KEYINPUT100), .B(KEYINPUT11), .Z(n509) );
  XNOR2_X1 U648 ( .A(n509), .B(n508), .ZN(n513) );
  NAND2_X1 U649 ( .A1(G214), .A2(n544), .ZN(n511) );
  XOR2_X1 U650 ( .A(KEYINPUT99), .B(KEYINPUT101), .Z(n510) );
  XNOR2_X1 U651 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U652 ( .A(n513), .B(n512), .ZN(n517) );
  XOR2_X1 U653 ( .A(KEYINPUT12), .B(G104), .Z(n514) );
  XNOR2_X1 U654 ( .A(n514), .B(n350), .ZN(n515) );
  XNOR2_X1 U655 ( .A(KEYINPUT10), .B(n518), .ZN(n865) );
  XNOR2_X1 U656 ( .A(n865), .B(G146), .ZN(n559) );
  XNOR2_X1 U657 ( .A(n519), .B(n559), .ZN(n753) );
  NOR2_X1 U658 ( .A1(n753), .A2(G902), .ZN(n520) );
  XNOR2_X1 U659 ( .A(n522), .B(n521), .ZN(n526) );
  AND2_X1 U660 ( .A1(n552), .A2(G217), .ZN(n532) );
  XNOR2_X2 U661 ( .A(G128), .B(G143), .ZN(n530) );
  XNOR2_X2 U662 ( .A(KEYINPUT65), .B(KEYINPUT87), .ZN(n529) );
  XNOR2_X2 U663 ( .A(n530), .B(n529), .ZN(n540) );
  XNOR2_X1 U664 ( .A(n540), .B(KEYINPUT103), .ZN(n531) );
  XNOR2_X1 U665 ( .A(n532), .B(n531), .ZN(n533) );
  NAND2_X1 U666 ( .A1(n768), .A2(n593), .ZN(n535) );
  INV_X1 U667 ( .A(G478), .ZN(n534) );
  INV_X1 U668 ( .A(n787), .ZN(n798) );
  AND2_X1 U669 ( .A1(n536), .A2(n704), .ZN(n538) );
  XNOR2_X1 U670 ( .A(KEYINPUT70), .B(G101), .ZN(n541) );
  XOR2_X1 U671 ( .A(G113), .B(G116), .Z(n543) );
  XNOR2_X1 U672 ( .A(n543), .B(n542), .ZN(n584) );
  NAND2_X1 U673 ( .A1(n544), .A2(G210), .ZN(n546) );
  XNOR2_X1 U674 ( .A(n617), .B(n550), .ZN(n551) );
  NAND2_X1 U675 ( .A1(G221), .A2(n552), .ZN(n557) );
  XNOR2_X1 U676 ( .A(G128), .B(G137), .ZN(n553) );
  XNOR2_X1 U677 ( .A(n359), .B(n553), .ZN(n555) );
  NAND2_X1 U678 ( .A1(n749), .A2(n593), .ZN(n566) );
  XOR2_X1 U679 ( .A(KEYINPUT81), .B(KEYINPUT25), .Z(n562) );
  XNOR2_X2 U680 ( .A(G902), .B(KEYINPUT15), .ZN(n728) );
  NAND2_X1 U681 ( .A1(n728), .A2(G234), .ZN(n560) );
  XNOR2_X1 U682 ( .A(n560), .B(KEYINPUT20), .ZN(n574) );
  NAND2_X1 U683 ( .A1(n574), .A2(G217), .ZN(n561) );
  XNOR2_X1 U684 ( .A(n562), .B(n561), .ZN(n564) );
  INV_X1 U685 ( .A(KEYINPUT82), .ZN(n563) );
  XNOR2_X1 U686 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X2 U687 ( .A(n566), .B(n565), .ZN(n693) );
  XNOR2_X1 U688 ( .A(n567), .B(KEYINPUT14), .ZN(n817) );
  NOR2_X1 U689 ( .A1(G900), .A2(n673), .ZN(n568) );
  NAND2_X1 U690 ( .A1(n817), .A2(n568), .ZN(n569) );
  XOR2_X1 U691 ( .A(KEYINPUT108), .B(n569), .Z(n572) );
  INV_X1 U692 ( .A(n817), .ZN(n570) );
  NAND2_X1 U693 ( .A1(G952), .A2(n870), .ZN(n674) );
  NOR2_X1 U694 ( .A1(n570), .A2(n674), .ZN(n571) );
  NOR2_X1 U695 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U696 ( .A(KEYINPUT88), .B(n573), .ZN(n625) );
  AND2_X1 U697 ( .A1(n574), .A2(G221), .ZN(n575) );
  XNOR2_X1 U698 ( .A(n575), .B(KEYINPUT21), .ZN(n819) );
  NAND2_X1 U699 ( .A1(n576), .A2(n819), .ZN(n651) );
  XNOR2_X1 U700 ( .A(n578), .B(n577), .ZN(n854) );
  XNOR2_X1 U701 ( .A(n854), .B(KEYINPUT73), .ZN(n579) );
  INV_X1 U702 ( .A(KEYINPUT74), .ZN(n581) );
  XNOR2_X1 U703 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U704 ( .A(n584), .B(n583), .ZN(n852) );
  XNOR2_X1 U705 ( .A(n586), .B(n585), .ZN(n589) );
  NAND2_X1 U706 ( .A1(n870), .A2(G224), .ZN(n587) );
  XNOR2_X1 U707 ( .A(n587), .B(KEYINPUT18), .ZN(n588) );
  XNOR2_X1 U708 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U709 ( .A(n852), .B(n590), .ZN(n591) );
  NAND2_X1 U710 ( .A1(n593), .A2(n592), .ZN(n601) );
  INV_X1 U711 ( .A(n601), .ZN(n609) );
  INV_X1 U712 ( .A(KEYINPUT19), .ZN(n594) );
  NAND2_X1 U713 ( .A1(n609), .A2(n594), .ZN(n596) );
  INV_X1 U714 ( .A(G210), .ZN(n607) );
  NAND2_X1 U715 ( .A1(n607), .A2(n594), .ZN(n595) );
  AND2_X1 U716 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U717 ( .A1(n601), .A2(G210), .ZN(n632) );
  INV_X1 U718 ( .A(G214), .ZN(n597) );
  NAND2_X1 U719 ( .A1(n597), .A2(KEYINPUT19), .ZN(n606) );
  OR2_X1 U720 ( .A1(n632), .A2(n606), .ZN(n598) );
  NAND2_X1 U721 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U722 ( .A1(n631), .A2(n600), .ZN(n605) );
  INV_X1 U723 ( .A(n728), .ZN(n735) );
  NAND2_X1 U724 ( .A1(n600), .A2(n735), .ZN(n603) );
  NAND2_X1 U725 ( .A1(n601), .A2(G214), .ZN(n834) );
  OR2_X1 U726 ( .A1(n834), .A2(KEYINPUT19), .ZN(n602) );
  AND2_X1 U727 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U728 ( .A1(n605), .A2(n604), .ZN(n616) );
  INV_X1 U729 ( .A(n606), .ZN(n608) );
  NAND2_X1 U730 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U731 ( .A1(n609), .A2(KEYINPUT19), .ZN(n610) );
  AND2_X1 U732 ( .A1(n611), .A2(n610), .ZN(n613) );
  OR2_X1 U733 ( .A1(n632), .A2(KEYINPUT19), .ZN(n612) );
  NAND2_X1 U734 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U735 ( .A1(n631), .A2(n362), .ZN(n615) );
  NOR2_X1 U736 ( .A1(n648), .A2(n679), .ZN(n621) );
  NAND2_X1 U737 ( .A1(n870), .A2(G227), .ZN(n618) );
  XNOR2_X2 U738 ( .A(n620), .B(n619), .ZN(n656) );
  XNOR2_X1 U739 ( .A(n622), .B(KEYINPUT76), .ZN(n624) );
  INV_X1 U740 ( .A(n793), .ZN(n788) );
  NAND2_X1 U741 ( .A1(n788), .A2(KEYINPUT47), .ZN(n623) );
  NAND2_X1 U742 ( .A1(n624), .A2(n623), .ZN(n636) );
  NAND2_X1 U743 ( .A1(n628), .A2(n627), .ZN(n629) );
  OR2_X2 U744 ( .A1(n631), .A2(n735), .ZN(n633) );
  INV_X1 U745 ( .A(n704), .ZN(n838) );
  INV_X1 U746 ( .A(KEYINPUT78), .ZN(n638) );
  XNOR2_X1 U747 ( .A(n638), .B(KEYINPUT38), .ZN(n639) );
  BUF_X1 U748 ( .A(n645), .Z(n640) );
  INV_X1 U749 ( .A(n352), .ZN(n652) );
  NAND2_X1 U750 ( .A1(n644), .A2(n643), .ZN(n836) );
  XNOR2_X1 U751 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n647) );
  OR2_X1 U752 ( .A1(n656), .A2(n648), .ZN(n649) );
  NOR2_X1 U753 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U754 ( .A(KEYINPUT105), .B(KEYINPUT6), .ZN(n654) );
  XNOR2_X1 U755 ( .A(n655), .B(KEYINPUT36), .ZN(n658) );
  NOR2_X1 U756 ( .A1(n787), .A2(n660), .ZN(n803) );
  XOR2_X1 U757 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n664) );
  INV_X1 U758 ( .A(n661), .ZN(n662) );
  NAND2_X1 U759 ( .A1(n662), .A2(n657), .ZN(n663) );
  XNOR2_X1 U760 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U761 ( .A(n665), .B(KEYINPUT110), .ZN(n666) );
  INV_X1 U762 ( .A(KEYINPUT91), .ZN(n730) );
  NOR2_X1 U763 ( .A1(n730), .A2(KEYINPUT67), .ZN(n667) );
  NAND2_X1 U764 ( .A1(n730), .A2(KEYINPUT67), .ZN(n722) );
  OR2_X1 U765 ( .A1(n722), .A2(KEYINPUT2), .ZN(n668) );
  NAND2_X1 U766 ( .A1(n736), .A2(n668), .ZN(n717) );
  XNOR2_X1 U767 ( .A(n696), .B(KEYINPUT107), .ZN(n670) );
  NAND2_X1 U768 ( .A1(n670), .A2(n686), .ZN(n672) );
  INV_X1 U769 ( .A(KEYINPUT33), .ZN(n671) );
  NOR2_X1 U770 ( .A1(G898), .A2(n673), .ZN(n676) );
  INV_X1 U771 ( .A(n674), .ZN(n675) );
  OR2_X1 U772 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U773 ( .A1(n817), .A2(n677), .ZN(n678) );
  NOR2_X2 U774 ( .A1(n679), .A2(n678), .ZN(n682) );
  INV_X1 U775 ( .A(KEYINPUT69), .ZN(n680) );
  XNOR2_X1 U776 ( .A(n680), .B(KEYINPUT0), .ZN(n681) );
  INV_X1 U777 ( .A(n703), .ZN(n685) );
  INV_X1 U778 ( .A(n836), .ZN(n683) );
  NAND2_X1 U779 ( .A1(n683), .A2(n819), .ZN(n684) );
  INV_X1 U780 ( .A(n686), .ZN(n706) );
  XNOR2_X1 U781 ( .A(n706), .B(KEYINPUT86), .ZN(n688) );
  XNOR2_X1 U782 ( .A(n693), .B(KEYINPUT106), .ZN(n818) );
  INV_X1 U783 ( .A(n818), .ZN(n687) );
  AND2_X1 U784 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U785 ( .A1(n707), .A2(n690), .ZN(n692) );
  XNOR2_X1 U786 ( .A(KEYINPUT85), .B(KEYINPUT32), .ZN(n691) );
  NOR2_X1 U787 ( .A1(n700), .A2(n693), .ZN(n694) );
  AND2_X1 U788 ( .A1(n657), .A2(n694), .ZN(n695) );
  AND2_X1 U789 ( .A1(n707), .A2(n695), .ZN(n758) );
  OR2_X1 U790 ( .A1(n696), .A2(n824), .ZN(n698) );
  INV_X1 U791 ( .A(KEYINPUT98), .ZN(n697) );
  NAND2_X1 U792 ( .A1(n830), .A2(n703), .ZN(n699) );
  XNOR2_X1 U793 ( .A(n699), .B(KEYINPUT31), .ZN(n799) );
  NOR2_X1 U794 ( .A1(n700), .A2(n822), .ZN(n701) );
  AND2_X1 U795 ( .A1(n703), .A2(n702), .ZN(n783) );
  NAND2_X1 U796 ( .A1(n705), .A2(n704), .ZN(n712) );
  NAND2_X1 U797 ( .A1(n707), .A2(n706), .ZN(n709) );
  INV_X1 U798 ( .A(KEYINPUT93), .ZN(n708) );
  XNOR2_X1 U799 ( .A(n709), .B(n708), .ZN(n711) );
  NAND2_X1 U800 ( .A1(n657), .A2(n818), .ZN(n710) );
  AND2_X1 U801 ( .A1(n712), .A2(n760), .ZN(n713) );
  XNOR2_X1 U802 ( .A(KEYINPUT92), .B(KEYINPUT45), .ZN(n715) );
  INV_X1 U803 ( .A(KEYINPUT64), .ZN(n714) );
  XNOR2_X1 U804 ( .A(n715), .B(n714), .ZN(n716) );
  INV_X1 U805 ( .A(KEYINPUT2), .ZN(n812) );
  OR2_X1 U806 ( .A1(n728), .A2(n812), .ZN(n718) );
  NAND2_X1 U807 ( .A1(n718), .A2(KEYINPUT67), .ZN(n719) );
  INV_X1 U808 ( .A(KEYINPUT67), .ZN(n720) );
  NAND2_X1 U809 ( .A1(n720), .A2(KEYINPUT2), .ZN(n721) );
  NAND2_X1 U810 ( .A1(n735), .A2(n721), .ZN(n724) );
  NAND2_X1 U811 ( .A1(n728), .A2(n722), .ZN(n723) );
  AND2_X1 U812 ( .A1(n724), .A2(n723), .ZN(n725) );
  OR2_X1 U813 ( .A1(KEYINPUT91), .A2(KEYINPUT67), .ZN(n727) );
  NOR2_X1 U814 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U815 ( .A1(n812), .A2(KEYINPUT67), .ZN(n731) );
  NOR2_X1 U816 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U817 ( .A1(n735), .A2(n732), .ZN(n733) );
  OR2_X1 U818 ( .A1(n736), .A2(n735), .ZN(n737) );
  INV_X1 U819 ( .A(KEYINPUT79), .ZN(n738) );
  INV_X1 U820 ( .A(KEYINPUT66), .ZN(n741) );
  NAND2_X1 U821 ( .A1(n767), .A2(G210), .ZN(n746) );
  XNOR2_X1 U822 ( .A(KEYINPUT94), .B(KEYINPUT54), .ZN(n743) );
  XNOR2_X1 U823 ( .A(n743), .B(KEYINPUT55), .ZN(n744) );
  XNOR2_X1 U824 ( .A(n746), .B(n745), .ZN(n748) );
  INV_X1 U825 ( .A(G952), .ZN(n747) );
  NAND2_X1 U826 ( .A1(n767), .A2(G217), .ZN(n751) );
  XNOR2_X1 U827 ( .A(n751), .B(n750), .ZN(n752) );
  NAND2_X1 U828 ( .A1(n767), .A2(G475), .ZN(n756) );
  XNOR2_X1 U829 ( .A(KEYINPUT96), .B(KEYINPUT59), .ZN(n754) );
  XNOR2_X1 U830 ( .A(n756), .B(n755), .ZN(n757) );
  XOR2_X1 U831 ( .A(G110), .B(n758), .Z(G12) );
  XOR2_X1 U832 ( .A(n759), .B(G140), .Z(G42) );
  XNOR2_X1 U833 ( .A(n760), .B(G101), .ZN(G3) );
  XOR2_X1 U834 ( .A(n761), .B(G122), .Z(G24) );
  XOR2_X1 U835 ( .A(n350), .B(n762), .Z(G45) );
  NAND2_X1 U836 ( .A1(n767), .A2(G472), .ZN(n764) );
  XNOR2_X1 U837 ( .A(n764), .B(n763), .ZN(n765) );
  NAND2_X1 U838 ( .A1(n765), .A2(n770), .ZN(n766) );
  XNOR2_X1 U839 ( .A(n766), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U840 ( .A1(n772), .A2(G478), .ZN(n769) );
  INV_X1 U841 ( .A(n770), .ZN(n779) );
  NOR2_X1 U842 ( .A1(n771), .A2(n779), .ZN(G63) );
  NAND2_X1 U843 ( .A1(n772), .A2(G469), .ZN(n778) );
  XOR2_X1 U844 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n774) );
  XNOR2_X1 U845 ( .A(n774), .B(KEYINPUT58), .ZN(n775) );
  XNOR2_X1 U846 ( .A(n776), .B(n775), .ZN(n777) );
  XNOR2_X1 U847 ( .A(n778), .B(n777), .ZN(n780) );
  NOR2_X1 U848 ( .A1(n780), .A2(n779), .ZN(G54) );
  XOR2_X1 U849 ( .A(G104), .B(KEYINPUT113), .Z(n782) );
  NAND2_X1 U850 ( .A1(n783), .A2(n352), .ZN(n781) );
  XNOR2_X1 U851 ( .A(n782), .B(n781), .ZN(G6) );
  XOR2_X1 U852 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n785) );
  NAND2_X1 U853 ( .A1(n783), .A2(n798), .ZN(n784) );
  XNOR2_X1 U854 ( .A(n785), .B(n784), .ZN(n786) );
  XNOR2_X1 U855 ( .A(G107), .B(n786), .ZN(G9) );
  NOR2_X1 U856 ( .A1(n788), .A2(n787), .ZN(n792) );
  XOR2_X1 U857 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n790) );
  XNOR2_X1 U858 ( .A(G128), .B(KEYINPUT29), .ZN(n789) );
  XNOR2_X1 U859 ( .A(n790), .B(n789), .ZN(n791) );
  XNOR2_X1 U860 ( .A(n792), .B(n791), .ZN(G30) );
  NAND2_X1 U861 ( .A1(n793), .A2(n352), .ZN(n794) );
  XNOR2_X1 U862 ( .A(n794), .B(KEYINPUT116), .ZN(n795) );
  XNOR2_X1 U863 ( .A(G146), .B(n795), .ZN(G48) );
  XOR2_X1 U864 ( .A(G113), .B(KEYINPUT117), .Z(n797) );
  NAND2_X1 U865 ( .A1(n799), .A2(n352), .ZN(n796) );
  XNOR2_X1 U866 ( .A(n797), .B(n796), .ZN(G15) );
  NAND2_X1 U867 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U868 ( .A(n800), .B(KEYINPUT118), .ZN(n801) );
  XNOR2_X1 U869 ( .A(G116), .B(n801), .ZN(G18) );
  XNOR2_X1 U870 ( .A(n802), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U871 ( .A(G134), .B(n803), .Z(G36) );
  NOR2_X1 U872 ( .A1(n351), .A2(n805), .ZN(n806) );
  NOR2_X1 U873 ( .A1(n806), .A2(G953), .ZN(n850) );
  INV_X1 U874 ( .A(n807), .ZN(n816) );
  INV_X1 U875 ( .A(n869), .ZN(n809) );
  NAND2_X1 U876 ( .A1(n809), .A2(n812), .ZN(n810) );
  XNOR2_X1 U877 ( .A(n810), .B(KEYINPUT90), .ZN(n814) );
  BUF_X1 U878 ( .A(n811), .Z(n857) );
  NAND2_X1 U879 ( .A1(n857), .A2(n812), .ZN(n813) );
  NAND2_X1 U880 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U881 ( .A1(n816), .A2(n815), .ZN(n848) );
  NAND2_X1 U882 ( .A1(G952), .A2(n817), .ZN(n846) );
  NOR2_X1 U883 ( .A1(n819), .A2(n818), .ZN(n821) );
  XNOR2_X1 U884 ( .A(KEYINPUT49), .B(KEYINPUT119), .ZN(n820) );
  XNOR2_X1 U885 ( .A(n821), .B(n820), .ZN(n827) );
  NAND2_X1 U886 ( .A1(n657), .A2(n822), .ZN(n823) );
  XNOR2_X1 U887 ( .A(n823), .B(KEYINPUT50), .ZN(n825) );
  NAND2_X1 U888 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U889 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U890 ( .A(n828), .B(KEYINPUT120), .ZN(n829) );
  NOR2_X1 U891 ( .A1(n830), .A2(n829), .ZN(n831) );
  XOR2_X1 U892 ( .A(KEYINPUT51), .B(n831), .Z(n832) );
  NOR2_X1 U893 ( .A1(n805), .A2(n832), .ZN(n843) );
  NOR2_X1 U894 ( .A1(n834), .A2(n833), .ZN(n835) );
  NOR2_X1 U895 ( .A1(n836), .A2(n835), .ZN(n841) );
  NOR2_X1 U896 ( .A1(n838), .A2(n837), .ZN(n839) );
  XOR2_X1 U897 ( .A(KEYINPUT121), .B(n839), .Z(n840) );
  NOR2_X1 U898 ( .A1(n841), .A2(n840), .ZN(n842) );
  NOR2_X1 U899 ( .A1(n843), .A2(n507), .ZN(n844) );
  XNOR2_X1 U900 ( .A(n844), .B(KEYINPUT52), .ZN(n845) );
  NOR2_X1 U901 ( .A1(n846), .A2(n845), .ZN(n847) );
  NOR2_X1 U902 ( .A1(n848), .A2(n847), .ZN(n849) );
  NAND2_X1 U903 ( .A1(n850), .A2(n849), .ZN(n851) );
  XOR2_X1 U904 ( .A(KEYINPUT53), .B(n851), .Z(G75) );
  XOR2_X1 U905 ( .A(G101), .B(n852), .Z(n853) );
  XNOR2_X1 U906 ( .A(n854), .B(n853), .ZN(n856) );
  NOR2_X1 U907 ( .A1(G898), .A2(n870), .ZN(n855) );
  NOR2_X1 U908 ( .A1(n856), .A2(n855), .ZN(n864) );
  NOR2_X1 U909 ( .A1(n857), .A2(G953), .ZN(n858) );
  XNOR2_X1 U910 ( .A(n858), .B(KEYINPUT125), .ZN(n862) );
  NAND2_X1 U911 ( .A1(G953), .A2(G224), .ZN(n859) );
  XNOR2_X1 U912 ( .A(KEYINPUT61), .B(n859), .ZN(n860) );
  NAND2_X1 U913 ( .A1(n860), .A2(G898), .ZN(n861) );
  NAND2_X1 U914 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U915 ( .A(n864), .B(n863), .ZN(G69) );
  XNOR2_X1 U916 ( .A(n866), .B(n865), .ZN(n867) );
  XNOR2_X1 U917 ( .A(n868), .B(n867), .ZN(n873) );
  XOR2_X1 U918 ( .A(n873), .B(n869), .Z(n871) );
  NAND2_X1 U919 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U920 ( .A(n872), .B(KEYINPUT126), .ZN(n878) );
  XNOR2_X1 U921 ( .A(G227), .B(n873), .ZN(n874) );
  NAND2_X1 U922 ( .A1(n874), .A2(G900), .ZN(n875) );
  XOR2_X1 U923 ( .A(KEYINPUT127), .B(n875), .Z(n876) );
  NAND2_X1 U924 ( .A1(G953), .A2(n876), .ZN(n877) );
  NAND2_X1 U925 ( .A1(n878), .A2(n877), .ZN(G72) );
endmodule

