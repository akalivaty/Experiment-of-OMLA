//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n544, new_n545,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n593, new_n594, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT66), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  NAND2_X1  g033(.A1(new_n453), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(new_n456), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT67), .ZN(G319));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n463), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n463), .A2(G137), .ZN(new_n467));
  NAND2_X1  g042(.A1(G101), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(G160));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n473), .A2(new_n465), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  OAI211_X1 g056(.A(G138), .B(new_n465), .C1(new_n471), .C2(new_n472), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n463), .A2(KEYINPUT4), .A3(G138), .A4(new_n465), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g061(.A(G126), .B(G2105), .C1(new_n471), .C2(new_n472), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n486), .A2(new_n491), .ZN(G164));
  NAND2_X1  g067(.A1(KEYINPUT68), .A2(G651), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT6), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT69), .A2(G651), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n495), .A2(new_n496), .A3(KEYINPUT6), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n498), .A2(G50), .A3(G543), .A4(new_n499), .ZN(new_n500));
  XNOR2_X1  g075(.A(new_n500), .B(KEYINPUT70), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n498), .A2(new_n499), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(G75), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G62), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n506), .A2(G88), .B1(new_n509), .B2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n501), .A2(new_n510), .ZN(G303));
  INV_X1    g086(.A(G303), .ZN(G166));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n502), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G51), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n506), .A2(G89), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n517), .A2(KEYINPUT7), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(KEYINPUT7), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(new_n513), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(G63), .A2(G651), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n518), .A2(new_n519), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n515), .A2(new_n516), .A3(new_n525), .ZN(G168));
  NAND2_X1  g101(.A1(new_n514), .A2(G52), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n506), .A2(G90), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G651), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n527), .A2(new_n528), .A3(new_n531), .ZN(G301));
  INV_X1    g107(.A(G301), .ZN(G171));
  AOI22_X1  g108(.A1(G43), .A2(new_n514), .B1(new_n506), .B2(G81), .ZN(new_n534));
  NAND2_X1  g109(.A1(G68), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G56), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n505), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n530), .B1(new_n537), .B2(KEYINPUT71), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n538), .B1(KEYINPUT71), .B2(new_n537), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND4_X1  g120(.A1(G319), .A2(G483), .A3(G661), .A4(new_n545), .ZN(G188));
  AOI22_X1  g121(.A1(new_n496), .A2(new_n495), .B1(new_n493), .B2(KEYINPUT6), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n495), .A2(new_n496), .A3(KEYINPUT6), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g124(.A1(new_n549), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n498), .A2(G53), .A3(G543), .A4(new_n499), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT9), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n549), .A2(G91), .A3(new_n523), .ZN(new_n554));
  INV_X1    g129(.A(G65), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n505), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g131(.A1(G78), .A2(G543), .ZN(new_n557));
  OAI21_X1  g132(.A(G651), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n550), .A2(new_n553), .A3(new_n554), .A4(new_n558), .ZN(G299));
  NAND3_X1  g134(.A1(new_n515), .A2(new_n516), .A3(new_n525), .ZN(G286));
  NAND2_X1  g135(.A1(new_n514), .A2(G49), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n506), .A2(G87), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(G288));
  INV_X1    g139(.A(G61), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n565), .B1(new_n521), .B2(new_n522), .ZN(new_n566));
  AND2_X1   g141(.A1(G73), .A2(G543), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n498), .A2(G86), .A3(new_n499), .A4(new_n523), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n498), .A2(G48), .A3(G543), .A4(new_n499), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G305));
  NAND2_X1  g146(.A1(new_n514), .A2(G47), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n549), .A2(new_n523), .ZN(new_n574));
  XNOR2_X1  g149(.A(KEYINPUT72), .B(G85), .ZN(new_n575));
  OAI221_X1 g150(.A(new_n572), .B1(new_n530), .B2(new_n573), .C1(new_n574), .C2(new_n575), .ZN(G290));
  NAND2_X1  g151(.A1(G301), .A2(G868), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n498), .A2(G92), .A3(new_n499), .A4(new_n523), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT10), .ZN(new_n579));
  INV_X1    g154(.A(G66), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n580), .B1(new_n521), .B2(new_n522), .ZN(new_n581));
  NAND2_X1  g156(.A1(G79), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT73), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT73), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n585), .B(new_n582), .C1(new_n505), .C2(new_n580), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(G651), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n549), .A2(G54), .A3(G543), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n579), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n577), .B1(new_n590), .B2(G868), .ZN(G321));
  XOR2_X1   g166(.A(G321), .B(KEYINPUT74), .Z(G284));
  INV_X1    g167(.A(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(G299), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(G168), .B2(new_n593), .ZN(G297));
  OAI21_X1  g170(.A(new_n594), .B1(G168), .B2(new_n593), .ZN(G280));
  INV_X1    g171(.A(G559), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n590), .B1(new_n597), .B2(G860), .ZN(G148));
  NAND2_X1  g173(.A1(new_n590), .A2(new_n597), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT75), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(new_n593), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n541), .A2(new_n593), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(KEYINPUT11), .Z(G282));
  INV_X1    g179(.A(new_n603), .ZN(G323));
  NAND2_X1  g180(.A1(new_n474), .A2(G2104), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT13), .ZN(new_n608));
  XOR2_X1   g183(.A(KEYINPUT76), .B(G2100), .Z(new_n609));
  OR2_X1    g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n474), .A2(G135), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n476), .A2(G123), .ZN(new_n613));
  NOR2_X1   g188(.A1(G99), .A2(G2105), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(new_n465), .B2(G111), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n612), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G2096), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n610), .A2(new_n611), .A3(new_n618), .ZN(G156));
  XNOR2_X1  g194(.A(G2427), .B(G2430), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT77), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(KEYINPUT14), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G1341), .B(G1348), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2443), .B(G2446), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2451), .B(G2454), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT78), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n630), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(G14), .A3(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(G401));
  XOR2_X1   g212(.A(G2072), .B(G2078), .Z(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT17), .Z(new_n639));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  INV_X1    g218(.A(new_n640), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(new_n638), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n642), .B(new_n643), .C1(new_n641), .C2(new_n645), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n643), .A2(new_n638), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT18), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(new_n617), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2100), .ZN(G227));
  XNOR2_X1  g226(.A(G1961), .B(G1966), .ZN(new_n652));
  AND2_X1   g227(.A1(new_n652), .A2(KEYINPUT79), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(KEYINPUT79), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1956), .B(G2474), .ZN(new_n655));
  OR3_X1    g230(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT20), .Z(new_n660));
  OAI21_X1  g235(.A(new_n655), .B1(new_n653), .B2(new_n654), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n661), .A2(new_n658), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT80), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n656), .A2(new_n661), .A3(new_n658), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n660), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G1986), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  INV_X1    g246(.A(G1981), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n668), .A2(new_n669), .A3(new_n673), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(G229));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G23), .ZN(new_n679));
  INV_X1    g254(.A(G288), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(new_n678), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT33), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G1976), .ZN(new_n683));
  MUX2_X1   g258(.A(G6), .B(G305), .S(G16), .Z(new_n684));
  XOR2_X1   g259(.A(KEYINPUT32), .B(G1981), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT84), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(new_n687));
  NOR2_X1   g262(.A1(G16), .A2(G22), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(G166), .B2(G16), .ZN(new_n689));
  INV_X1    g264(.A(G1971), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n683), .A2(new_n687), .A3(new_n691), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n692), .A2(KEYINPUT34), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(KEYINPUT34), .ZN(new_n694));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n695), .A2(G25), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n476), .A2(G119), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT81), .ZN(new_n698));
  OR2_X1    g273(.A1(G95), .A2(G2105), .ZN(new_n699));
  INV_X1    g274(.A(G2104), .ZN(new_n700));
  INV_X1    g275(.A(G107), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(G2105), .ZN(new_n702));
  AOI22_X1  g277(.A1(new_n474), .A2(G131), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n696), .B1(new_n704), .B2(G29), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT82), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT35), .B(G1991), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n706), .B(new_n707), .Z(new_n708));
  AND3_X1   g283(.A1(new_n678), .A2(KEYINPUT83), .A3(G24), .ZN(new_n709));
  AOI21_X1  g284(.A(KEYINPUT83), .B1(new_n678), .B2(G24), .ZN(new_n710));
  AOI211_X1 g285(.A(new_n709), .B(new_n710), .C1(G290), .C2(G16), .ZN(new_n711));
  INV_X1    g286(.A(G1986), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT36), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(KEYINPUT85), .B2(new_n715), .ZN(new_n716));
  NOR3_X1   g291(.A1(new_n708), .A2(new_n713), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n693), .A2(new_n694), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n718), .A2(KEYINPUT85), .A3(new_n715), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n717), .A2(new_n694), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n715), .A2(KEYINPUT85), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n720), .A2(new_n721), .A3(new_n693), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n678), .A2(G19), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(new_n541), .B2(new_n678), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(G1341), .Z(new_n725));
  NAND2_X1  g300(.A1(new_n695), .A2(G26), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT28), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n474), .A2(G140), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n476), .A2(G128), .ZN(new_n729));
  OR2_X1    g304(.A1(G104), .A2(G2105), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n730), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n728), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G29), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n733), .A2(KEYINPUT86), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(KEYINPUT86), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n727), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G2067), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n590), .A2(new_n678), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G4), .B2(new_n678), .ZN(new_n740));
  INV_X1    g315(.A(G1348), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n725), .A2(new_n738), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT87), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n695), .A2(G35), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G162), .B2(new_n695), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT93), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT29), .ZN(new_n749));
  INV_X1    g324(.A(G2090), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(KEYINPUT94), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n695), .A2(G32), .ZN(new_n753));
  NAND3_X1  g328(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT26), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n476), .A2(G129), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n465), .A2(G105), .A3(G2104), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT91), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  AOI211_X1 g334(.A(new_n755), .B(new_n759), .C1(G141), .C2(new_n474), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n753), .B1(new_n760), .B2(new_n695), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT27), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1996), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n695), .B1(KEYINPUT24), .B2(G34), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(KEYINPUT24), .B2(G34), .ZN(new_n765));
  INV_X1    g340(.A(G160), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n765), .B1(new_n766), .B2(G29), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT90), .ZN(new_n768));
  INV_X1    g343(.A(G2084), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n695), .A2(G27), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G164), .B2(new_n695), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2078), .ZN(new_n773));
  INV_X1    g348(.A(G1961), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n678), .A2(G5), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G301), .B2(G16), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n773), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n752), .A2(new_n763), .A3(new_n770), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n678), .A2(G21), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G168), .B2(new_n678), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(G1966), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n616), .A2(new_n695), .ZN(new_n782));
  INV_X1    g357(.A(G28), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(KEYINPUT30), .ZN(new_n784));
  AOI21_X1  g359(.A(G29), .B1(new_n783), .B2(KEYINPUT30), .ZN(new_n785));
  OR2_X1    g360(.A1(KEYINPUT31), .A2(G11), .ZN(new_n786));
  NAND2_X1  g361(.A1(KEYINPUT31), .A2(G11), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n784), .A2(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n781), .A2(new_n782), .A3(new_n788), .ZN(new_n789));
  OAI22_X1  g364(.A1(new_n780), .A2(G1966), .B1(new_n776), .B2(new_n774), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT92), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n751), .B2(KEYINPUT94), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT88), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT25), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(G115), .A2(G2104), .ZN(new_n798));
  INV_X1    g373(.A(G127), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n473), .B2(new_n799), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n800), .A2(G2105), .B1(new_n474), .B2(G139), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n795), .A2(new_n796), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n797), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(KEYINPUT89), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT89), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n797), .A2(new_n801), .A3(new_n805), .A4(new_n802), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  MUX2_X1   g382(.A(G33), .B(new_n807), .S(G29), .Z(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(G2072), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n678), .A2(G20), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT23), .ZN(new_n811));
  AND4_X1   g386(.A1(new_n550), .A2(new_n553), .A3(new_n554), .A4(new_n558), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(new_n678), .ZN(new_n813));
  INV_X1    g388(.A(G1956), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n809), .B(new_n815), .C1(new_n749), .C2(new_n750), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n778), .A2(new_n793), .A3(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n719), .A2(new_n722), .A3(new_n745), .A4(new_n817), .ZN(G150));
  INV_X1    g393(.A(G150), .ZN(G311));
  NAND2_X1  g394(.A1(new_n514), .A2(G55), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n506), .A2(G93), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n820), .B(new_n821), .C1(new_n530), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G860), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT96), .B(KEYINPUT37), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n540), .A2(new_n823), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n540), .A2(new_n823), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n590), .A2(G559), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n831), .B(new_n832), .Z(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n835));
  INV_X1    g410(.A(G860), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n834), .B2(KEYINPUT39), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n826), .B1(new_n835), .B2(new_n837), .ZN(G145));
  NAND2_X1  g413(.A1(new_n474), .A2(G142), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n476), .A2(G130), .ZN(new_n840));
  NOR2_X1   g415(.A1(G106), .A2(G2105), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(new_n465), .B2(G118), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n839), .B(new_n840), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n760), .B(new_n843), .Z(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n732), .B1(new_n804), .B2(new_n806), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT97), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n491), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n487), .A2(new_n490), .A3(KEYINPUT97), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n849), .A2(new_n484), .A3(new_n485), .A4(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n804), .A2(new_n806), .A3(new_n732), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n847), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n704), .B(new_n607), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  AND3_X1   g431(.A1(new_n804), .A2(new_n806), .A3(new_n732), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n851), .B1(new_n857), .B2(new_n846), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n854), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n856), .B1(new_n854), .B2(new_n858), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n845), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n854), .A2(new_n858), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n855), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n854), .A2(new_n856), .A3(new_n858), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(new_n844), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(G160), .B(new_n616), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(G162), .ZN(new_n868));
  AOI21_X1  g443(.A(G37), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n861), .A2(new_n865), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT98), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT98), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n869), .A2(new_n874), .A3(new_n871), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n873), .A2(KEYINPUT40), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT40), .B1(new_n873), .B2(new_n875), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(G395));
  XNOR2_X1  g453(.A(new_n600), .B(new_n829), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(new_n590), .B2(G299), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n590), .A2(G299), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT10), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n578), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n578), .A2(new_n883), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n588), .B(new_n587), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n886), .A2(new_n812), .A3(KEYINPUT99), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n881), .A2(new_n882), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n879), .A2(new_n888), .ZN(new_n889));
  XOR2_X1   g464(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n890));
  OR2_X1    g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n886), .A2(new_n812), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n886), .A2(new_n812), .A3(KEYINPUT99), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT99), .B1(new_n886), .B2(new_n812), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n881), .A2(KEYINPUT100), .A3(new_n887), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n892), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n891), .B1(new_n898), .B2(KEYINPUT41), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n889), .B1(new_n900), .B2(new_n879), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT42), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n904));
  OAI221_X1 g479(.A(new_n889), .B1(KEYINPUT102), .B2(new_n904), .C1(new_n900), .C2(new_n879), .ZN(new_n905));
  XNOR2_X1  g480(.A(G290), .B(new_n680), .ZN(new_n906));
  XNOR2_X1  g481(.A(G303), .B(G305), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n908), .B1(KEYINPUT102), .B2(new_n904), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n903), .A2(new_n905), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n909), .B1(new_n903), .B2(new_n905), .ZN(new_n911));
  OAI21_X1  g486(.A(G868), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n823), .A2(new_n593), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(G295));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n913), .ZN(G331));
  INV_X1    g490(.A(new_n888), .ZN(new_n916));
  XNOR2_X1  g491(.A(G301), .B(G286), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n829), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n827), .A3(new_n828), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  AOI211_X1 g497(.A(new_n921), .B(new_n908), .C1(new_n899), .C2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G37), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n921), .B1(new_n899), .B2(new_n922), .ZN(new_n925));
  INV_X1    g500(.A(new_n908), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n923), .B1(new_n927), .B2(KEYINPUT103), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n929), .B(new_n924), .C1(new_n925), .C2(new_n926), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT43), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n925), .A2(new_n926), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n924), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n888), .A2(new_n890), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT104), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n898), .A2(KEYINPUT41), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n922), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n921), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n926), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n933), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT44), .B1(new_n931), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n940), .B1(new_n928), .B2(new_n930), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n933), .A2(new_n939), .A3(KEYINPUT43), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n942), .A2(new_n946), .ZN(G397));
  INV_X1    g522(.A(G1384), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT45), .B1(new_n851), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(KEYINPUT105), .B(G40), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n466), .A2(new_n469), .A3(new_n950), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n732), .B(G2067), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT108), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G1996), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n760), .B(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n952), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT109), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n704), .A2(new_n707), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n704), .A2(new_n707), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n952), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(G290), .A2(G1986), .ZN(new_n964));
  XOR2_X1   g539(.A(new_n964), .B(KEYINPUT106), .Z(new_n965));
  NAND2_X1  g540(.A1(G290), .A2(G1986), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT107), .ZN(new_n967));
  OR2_X1    g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n963), .B1(new_n952), .B2(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n568), .A2(new_n569), .A3(new_n570), .A4(new_n672), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n971));
  OR2_X1    g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n971), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XOR2_X1   g549(.A(KEYINPUT112), .B(G86), .Z(new_n975));
  OAI211_X1 g550(.A(new_n568), .B(new_n570), .C1(new_n574), .C2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(G1981), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n974), .A2(KEYINPUT49), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n972), .A2(new_n973), .B1(G1981), .B2(new_n976), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(KEYINPUT114), .A3(KEYINPUT49), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n951), .A2(new_n851), .A3(new_n948), .ZN(new_n984));
  XOR2_X1   g559(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(G8), .B(new_n984), .C1(new_n981), .C2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(G288), .A2(G1976), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n989), .A2(new_n990), .B1(new_n973), .B2(new_n972), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n984), .A2(G8), .ZN(new_n992));
  INV_X1    g567(.A(G137), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n468), .B1(new_n473), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n465), .ZN(new_n995));
  INV_X1    g570(.A(new_n950), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n995), .B(new_n996), .C1(new_n465), .C2(new_n464), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n948), .B1(new_n486), .B2(new_n491), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n997), .B1(KEYINPUT50), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n851), .A2(new_n1000), .A3(new_n948), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n999), .A2(new_n1001), .A3(new_n750), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n997), .B1(new_n1003), .B2(new_n998), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n851), .A2(KEYINPUT45), .A3(new_n948), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1971), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT110), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n1007), .A2(G8), .ZN(new_n1008));
  NAND2_X1  g583(.A1(G303), .A2(G8), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1006), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n999), .A2(new_n750), .A3(new_n1001), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1008), .A2(new_n1011), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1976), .ZN(new_n1017));
  NOR2_X1   g592(.A1(G288), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n992), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT52), .B1(G288), .B2(new_n1017), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT52), .B1(new_n992), .B2(new_n1018), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n989), .A2(new_n1023), .ZN(new_n1024));
  OAI22_X1  g599(.A1(new_n991), .A2(new_n992), .B1(new_n1016), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n987), .B1(new_n980), .B2(new_n982), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n989), .A2(new_n1023), .A3(KEYINPUT116), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n851), .A2(new_n948), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT50), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(new_n1033), .A3(new_n951), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1000), .B1(new_n851), .B2(new_n948), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT115), .B1(new_n1035), .B2(new_n997), .ZN(new_n1036));
  INV_X1    g611(.A(new_n998), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n1000), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1034), .A2(new_n1036), .A3(new_n750), .A4(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n1012), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(G8), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1011), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1016), .A2(new_n1029), .A3(new_n1030), .A4(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1966), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n951), .B1(new_n998), .B2(new_n1003), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1045), .B1(new_n1046), .B2(new_n949), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n999), .A2(new_n769), .A3(new_n1001), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(new_n1048), .A3(G168), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G8), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT51), .B1(new_n1050), .B2(KEYINPUT122), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT62), .ZN(new_n1052));
  AOI21_X1  g627(.A(G168), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1053));
  NOR2_X1   g628(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n1054));
  OAI211_X1 g629(.A(G8), .B(new_n1049), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1051), .A2(new_n1052), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G2078), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT53), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1046), .A2(new_n949), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n999), .A2(new_n1001), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1059), .B1(new_n774), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT124), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1004), .A2(new_n1057), .A3(new_n1005), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1063), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1061), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1056), .A2(G171), .A3(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1044), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT127), .B1(new_n1070), .B2(KEYINPUT62), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT127), .ZN(new_n1072));
  AOI211_X1 g647(.A(new_n1072), .B(new_n1052), .C1(new_n1051), .C2(new_n1055), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1025), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g650(.A(G301), .B(KEYINPUT54), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1061), .B(new_n1076), .C1(new_n1066), .C2(new_n1065), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1060), .A2(new_n774), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n469), .B(KEYINPUT125), .ZN(new_n1079));
  INV_X1    g654(.A(G40), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n466), .A2(new_n1080), .A3(new_n1058), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1005), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1078), .B1(new_n949), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1065), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1063), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1077), .B1(new_n1086), .B2(new_n1076), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n1070), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT126), .B1(new_n1044), .B2(new_n1088), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1076), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1066), .A2(new_n1065), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1091), .B1(new_n1092), .B2(new_n1083), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1093), .A2(new_n1077), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT126), .ZN(new_n1095));
  AND4_X1   g670(.A1(G8), .A2(new_n1015), .A3(new_n1011), .A4(new_n1007), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1011), .B1(new_n1040), .B2(G8), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1090), .A2(new_n1094), .A3(new_n1095), .A4(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1034), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n814), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n1102));
  NOR2_X1   g677(.A1(G299), .A2(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1103), .B(KEYINPUT120), .ZN(new_n1104));
  NAND2_X1  g679(.A1(G299), .A2(new_n1102), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT119), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT56), .B(G2072), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1101), .A2(new_n1107), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(G1348), .B1(new_n999), .B2(new_n1001), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n984), .A2(G2067), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(new_n886), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1107), .B1(new_n1101), .B2(new_n1111), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1113), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1114), .A2(new_n1115), .A3(new_n590), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT60), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT61), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1004), .A2(new_n956), .A3(new_n1005), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT58), .B(G1341), .Z(new_n1124));
  NAND2_X1  g699(.A1(new_n984), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n540), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  AND2_X1   g701(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1127));
  NOR2_X1   g702(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1128));
  OR3_X1    g703(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n886), .A2(KEYINPUT60), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1126), .A2(new_n1127), .B1(new_n1116), .B2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1121), .A2(new_n1122), .A3(new_n1129), .A4(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1121), .A2(KEYINPUT61), .A3(new_n1129), .A4(new_n1131), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1119), .A2(new_n1132), .B1(new_n1133), .B2(new_n1113), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1089), .A2(new_n1099), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1075), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(G168), .A2(G8), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1016), .A2(KEYINPUT63), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1024), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1008), .A2(new_n1015), .ZN(new_n1141));
  OAI211_X1 g716(.A(KEYINPUT118), .B(new_n1140), .C1(new_n1141), .C2(new_n1011), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT118), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1011), .B1(new_n1008), .B2(new_n1015), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1143), .B1(new_n1144), .B2(new_n1024), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1139), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1098), .A2(new_n1029), .A3(new_n1030), .A4(new_n1138), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT117), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT63), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1090), .A2(KEYINPUT117), .A3(new_n1098), .A4(new_n1138), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1146), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n969), .B1(new_n1136), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n954), .A2(new_n760), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT46), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n952), .A2(new_n956), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1153), .A2(new_n952), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1156), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT47), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n965), .A2(new_n952), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT48), .Z(new_n1160));
  OAI21_X1  g735(.A(new_n1158), .B1(new_n963), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n959), .A2(new_n961), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1162), .B1(G2067), .B2(new_n732), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1161), .B1(new_n952), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1152), .A2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g740(.A1(new_n944), .A2(new_n945), .ZN(new_n1167));
  NOR2_X1   g741(.A1(G227), .A2(new_n461), .ZN(new_n1168));
  NAND2_X1  g742(.A1(new_n1168), .A2(new_n636), .ZN(new_n1169));
  AOI21_X1  g743(.A(new_n1169), .B1(new_n675), .B2(new_n676), .ZN(new_n1170));
  INV_X1    g744(.A(new_n875), .ZN(new_n1171));
  AOI21_X1  g745(.A(new_n874), .B1(new_n869), .B2(new_n871), .ZN(new_n1172));
  OAI21_X1  g746(.A(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g747(.A1(new_n1167), .A2(new_n1173), .ZN(G308));
  OAI221_X1 g748(.A(new_n1170), .B1(new_n1171), .B2(new_n1172), .C1(new_n944), .C2(new_n945), .ZN(G225));
endmodule


