

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580;

  XNOR2_X1 U322 ( .A(KEYINPUT97), .B(n397), .ZN(n545) );
  XOR2_X1 U323 ( .A(KEYINPUT84), .B(G134GAT), .Z(n291) );
  XNOR2_X1 U324 ( .A(KEYINPUT85), .B(G127GAT), .ZN(n290) );
  XNOR2_X1 U325 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U326 ( .A(KEYINPUT0), .B(n292), .Z(n379) );
  XNOR2_X1 U327 ( .A(G120GAT), .B(G148GAT), .ZN(n293) );
  XNOR2_X1 U328 ( .A(n293), .B(G57GAT), .ZN(n335) );
  XOR2_X1 U329 ( .A(n335), .B(G85GAT), .Z(n295) );
  XOR2_X1 U330 ( .A(G113GAT), .B(G1GAT), .Z(n324) );
  XNOR2_X1 U331 ( .A(G29GAT), .B(n324), .ZN(n294) );
  XNOR2_X1 U332 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U333 ( .A(n379), .B(n296), .ZN(n310) );
  XOR2_X1 U334 ( .A(KEYINPUT96), .B(KEYINPUT6), .Z(n298) );
  XNOR2_X1 U335 ( .A(KEYINPUT94), .B(KEYINPUT5), .ZN(n297) );
  XNOR2_X1 U336 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U337 ( .A(KEYINPUT4), .B(n299), .Z(n301) );
  NAND2_X1 U338 ( .A1(G225GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U339 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U340 ( .A(n302), .B(KEYINPUT1), .Z(n308) );
  XNOR2_X1 U341 ( .A(G155GAT), .B(KEYINPUT92), .ZN(n303) );
  XNOR2_X1 U342 ( .A(n303), .B(KEYINPUT3), .ZN(n304) );
  XOR2_X1 U343 ( .A(n304), .B(KEYINPUT2), .Z(n306) );
  XNOR2_X1 U344 ( .A(G141GAT), .B(G162GAT), .ZN(n305) );
  XNOR2_X1 U345 ( .A(n306), .B(n305), .ZN(n347) );
  XNOR2_X1 U346 ( .A(n347), .B(KEYINPUT95), .ZN(n307) );
  XNOR2_X1 U347 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U348 ( .A(n310), .B(n309), .ZN(n397) );
  XOR2_X1 U349 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n312) );
  NAND2_X1 U350 ( .A1(G229GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U351 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U352 ( .A(n313), .B(KEYINPUT67), .Z(n321) );
  XOR2_X1 U353 ( .A(KEYINPUT8), .B(G50GAT), .Z(n315) );
  XNOR2_X1 U354 ( .A(G43GAT), .B(G29GAT), .ZN(n314) );
  XNOR2_X1 U355 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U356 ( .A(KEYINPUT7), .B(n316), .Z(n419) );
  XOR2_X1 U357 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n318) );
  XNOR2_X1 U358 ( .A(G197GAT), .B(G141GAT), .ZN(n317) );
  XNOR2_X1 U359 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U360 ( .A(n419), .B(n319), .ZN(n320) );
  XNOR2_X1 U361 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U362 ( .A(G15GAT), .B(G22GAT), .Z(n425) );
  XOR2_X1 U363 ( .A(n322), .B(n425), .Z(n326) );
  XNOR2_X1 U364 ( .A(G169GAT), .B(G36GAT), .ZN(n323) );
  XNOR2_X1 U365 ( .A(n323), .B(G8GAT), .ZN(n387) );
  XNOR2_X1 U366 ( .A(n324), .B(n387), .ZN(n325) );
  XNOR2_X1 U367 ( .A(n326), .B(n325), .ZN(n567) );
  XOR2_X1 U368 ( .A(n567), .B(KEYINPUT70), .Z(n551) );
  XNOR2_X1 U369 ( .A(G99GAT), .B(G85GAT), .ZN(n327) );
  XNOR2_X1 U370 ( .A(n327), .B(KEYINPUT75), .ZN(n402) );
  XOR2_X1 U371 ( .A(KEYINPUT72), .B(n402), .Z(n329) );
  NAND2_X1 U372 ( .A1(G230GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U373 ( .A(n329), .B(n328), .ZN(n339) );
  XOR2_X1 U374 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n331) );
  XNOR2_X1 U375 ( .A(KEYINPUT32), .B(KEYINPUT73), .ZN(n330) );
  XNOR2_X1 U376 ( .A(n331), .B(n330), .ZN(n333) );
  XNOR2_X1 U377 ( .A(G71GAT), .B(KEYINPUT71), .ZN(n332) );
  XNOR2_X1 U378 ( .A(n332), .B(KEYINPUT13), .ZN(n429) );
  XOR2_X1 U379 ( .A(n333), .B(n429), .Z(n337) );
  XNOR2_X1 U380 ( .A(G106GAT), .B(G78GAT), .ZN(n334) );
  XNOR2_X1 U381 ( .A(n334), .B(KEYINPUT74), .ZN(n354) );
  XNOR2_X1 U382 ( .A(n354), .B(n335), .ZN(n336) );
  XNOR2_X1 U383 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U384 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U385 ( .A(G92GAT), .B(G64GAT), .Z(n341) );
  XNOR2_X1 U386 ( .A(G176GAT), .B(KEYINPUT76), .ZN(n340) );
  XNOR2_X1 U387 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U388 ( .A(G204GAT), .B(n342), .ZN(n384) );
  XNOR2_X1 U389 ( .A(n343), .B(n384), .ZN(n571) );
  NAND2_X1 U390 ( .A1(n551), .A2(n571), .ZN(n457) );
  INV_X1 U391 ( .A(n457), .ZN(n443) );
  XOR2_X1 U392 ( .A(KEYINPUT98), .B(KEYINPUT26), .Z(n381) );
  XOR2_X1 U393 ( .A(KEYINPUT91), .B(G218GAT), .Z(n345) );
  XNOR2_X1 U394 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n344) );
  XNOR2_X1 U395 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U396 ( .A(G197GAT), .B(n346), .Z(n386) );
  XNOR2_X1 U397 ( .A(n386), .B(n347), .ZN(n361) );
  XOR2_X1 U398 ( .A(G148GAT), .B(KEYINPUT22), .Z(n349) );
  XNOR2_X1 U399 ( .A(G22GAT), .B(KEYINPUT24), .ZN(n348) );
  XNOR2_X1 U400 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U401 ( .A(G204GAT), .B(KEYINPUT89), .Z(n351) );
  XNOR2_X1 U402 ( .A(KEYINPUT23), .B(KEYINPUT90), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U404 ( .A(n353), .B(n352), .Z(n359) );
  XOR2_X1 U405 ( .A(KEYINPUT93), .B(n354), .Z(n356) );
  NAND2_X1 U406 ( .A1(G228GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U407 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U408 ( .A(G50GAT), .B(n357), .ZN(n358) );
  XNOR2_X1 U409 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U410 ( .A(n361), .B(n360), .ZN(n547) );
  XOR2_X1 U411 ( .A(G71GAT), .B(KEYINPUT20), .Z(n363) );
  XNOR2_X1 U412 ( .A(G113GAT), .B(G15GAT), .ZN(n362) );
  XNOR2_X1 U413 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U414 ( .A(G120GAT), .B(G176GAT), .Z(n365) );
  XNOR2_X1 U415 ( .A(G169GAT), .B(G43GAT), .ZN(n364) );
  XNOR2_X1 U416 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U417 ( .A(n367), .B(n366), .ZN(n377) );
  XOR2_X1 U418 ( .A(KEYINPUT86), .B(KEYINPUT17), .Z(n369) );
  XNOR2_X1 U419 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n368) );
  XNOR2_X1 U420 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U421 ( .A(KEYINPUT19), .B(n370), .Z(n390) );
  XOR2_X1 U422 ( .A(G190GAT), .B(G99GAT), .Z(n372) );
  XNOR2_X1 U423 ( .A(KEYINPUT88), .B(KEYINPUT87), .ZN(n371) );
  XNOR2_X1 U424 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U425 ( .A(n390), .B(n373), .Z(n375) );
  NAND2_X1 U426 ( .A1(G227GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U427 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U428 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U429 ( .A(n379), .B(n378), .ZN(n550) );
  NAND2_X1 U430 ( .A1(n547), .A2(n550), .ZN(n380) );
  XNOR2_X1 U431 ( .A(n381), .B(n380), .ZN(n565) );
  XOR2_X1 U432 ( .A(G190GAT), .B(KEYINPUT80), .Z(n403) );
  XOR2_X1 U433 ( .A(KEYINPUT81), .B(n403), .Z(n383) );
  NAND2_X1 U434 ( .A1(G226GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U435 ( .A(n383), .B(n382), .ZN(n385) );
  XNOR2_X1 U436 ( .A(n385), .B(n384), .ZN(n389) );
  XNOR2_X1 U437 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U438 ( .A(n389), .B(n388), .ZN(n391) );
  XNOR2_X1 U439 ( .A(n391), .B(n390), .ZN(n540) );
  XOR2_X1 U440 ( .A(n540), .B(KEYINPUT27), .Z(n398) );
  AND2_X1 U441 ( .A1(n565), .A2(n398), .ZN(n526) );
  NOR2_X1 U442 ( .A1(n550), .A2(n540), .ZN(n392) );
  NOR2_X1 U443 ( .A1(n547), .A2(n392), .ZN(n393) );
  XNOR2_X1 U444 ( .A(n393), .B(KEYINPUT25), .ZN(n394) );
  XNOR2_X1 U445 ( .A(KEYINPUT99), .B(n394), .ZN(n395) );
  NOR2_X1 U446 ( .A1(n526), .A2(n395), .ZN(n396) );
  NOR2_X1 U447 ( .A1(n397), .A2(n396), .ZN(n401) );
  INV_X1 U448 ( .A(n550), .ZN(n511) );
  XNOR2_X1 U449 ( .A(n547), .B(KEYINPUT28), .ZN(n450) );
  NOR2_X1 U450 ( .A1(n545), .A2(n450), .ZN(n399) );
  NAND2_X1 U451 ( .A1(n399), .A2(n398), .ZN(n513) );
  NOR2_X1 U452 ( .A1(n511), .A2(n513), .ZN(n400) );
  NOR2_X1 U453 ( .A1(n401), .A2(n400), .ZN(n453) );
  XOR2_X1 U454 ( .A(KEYINPUT16), .B(KEYINPUT83), .Z(n441) );
  XOR2_X1 U455 ( .A(n403), .B(n402), .Z(n405) );
  XNOR2_X1 U456 ( .A(G218GAT), .B(G162GAT), .ZN(n404) );
  XNOR2_X1 U457 ( .A(n405), .B(n404), .ZN(n418) );
  XOR2_X1 U458 ( .A(KEYINPUT11), .B(KEYINPUT78), .Z(n407) );
  XNOR2_X1 U459 ( .A(G134GAT), .B(KEYINPUT79), .ZN(n406) );
  XNOR2_X1 U460 ( .A(n407), .B(n406), .ZN(n411) );
  XOR2_X1 U461 ( .A(KEYINPUT77), .B(KEYINPUT10), .Z(n409) );
  XNOR2_X1 U462 ( .A(KEYINPUT9), .B(KEYINPUT66), .ZN(n408) );
  XNOR2_X1 U463 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U464 ( .A(n411), .B(n410), .Z(n416) );
  XOR2_X1 U465 ( .A(G92GAT), .B(G106GAT), .Z(n413) );
  NAND2_X1 U466 ( .A1(G232GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U467 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U468 ( .A(G36GAT), .B(n414), .ZN(n415) );
  XNOR2_X1 U469 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U470 ( .A(n418), .B(n417), .ZN(n421) );
  INV_X1 U471 ( .A(n419), .ZN(n420) );
  XOR2_X1 U472 ( .A(n421), .B(n420), .Z(n538) );
  XOR2_X1 U473 ( .A(G78GAT), .B(G211GAT), .Z(n423) );
  XNOR2_X1 U474 ( .A(G127GAT), .B(G183GAT), .ZN(n422) );
  XNOR2_X1 U475 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U476 ( .A(n425), .B(n424), .Z(n427) );
  NAND2_X1 U477 ( .A1(G231GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U478 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U479 ( .A(n428), .B(KEYINPUT81), .Z(n431) );
  XNOR2_X1 U480 ( .A(n429), .B(KEYINPUT12), .ZN(n430) );
  XNOR2_X1 U481 ( .A(n431), .B(n430), .ZN(n439) );
  XOR2_X1 U482 ( .A(G57GAT), .B(G155GAT), .Z(n433) );
  XNOR2_X1 U483 ( .A(G1GAT), .B(G8GAT), .ZN(n432) );
  XNOR2_X1 U484 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U485 ( .A(KEYINPUT82), .B(KEYINPUT14), .Z(n435) );
  XNOR2_X1 U486 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n434) );
  XNOR2_X1 U487 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U488 ( .A(n437), .B(n436), .Z(n438) );
  XNOR2_X1 U489 ( .A(n439), .B(n438), .ZN(n557) );
  NAND2_X1 U490 ( .A1(n538), .A2(n557), .ZN(n440) );
  XNOR2_X1 U491 ( .A(n441), .B(n440), .ZN(n442) );
  NOR2_X1 U492 ( .A1(n453), .A2(n442), .ZN(n471) );
  NAND2_X1 U493 ( .A1(n443), .A2(n471), .ZN(n451) );
  NOR2_X1 U494 ( .A1(n545), .A2(n451), .ZN(n444) );
  XOR2_X1 U495 ( .A(KEYINPUT34), .B(n444), .Z(n445) );
  XNOR2_X1 U496 ( .A(G1GAT), .B(n445), .ZN(G1324GAT) );
  NOR2_X1 U497 ( .A1(n540), .A2(n451), .ZN(n446) );
  XOR2_X1 U498 ( .A(G8GAT), .B(n446), .Z(G1325GAT) );
  NOR2_X1 U499 ( .A1(n550), .A2(n451), .ZN(n448) );
  XNOR2_X1 U500 ( .A(KEYINPUT100), .B(KEYINPUT35), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U502 ( .A(G15GAT), .B(n449), .ZN(G1326GAT) );
  INV_X1 U503 ( .A(n450), .ZN(n495) );
  NOR2_X1 U504 ( .A1(n495), .A2(n451), .ZN(n452) );
  XOR2_X1 U505 ( .A(G22GAT), .B(n452), .Z(G1327GAT) );
  INV_X1 U506 ( .A(n557), .ZN(n575) );
  XNOR2_X1 U507 ( .A(KEYINPUT36), .B(n538), .ZN(n578) );
  NOR2_X1 U508 ( .A1(n578), .A2(n453), .ZN(n454) );
  NAND2_X1 U509 ( .A1(n575), .A2(n454), .ZN(n455) );
  XNOR2_X1 U510 ( .A(KEYINPUT37), .B(n455), .ZN(n456) );
  XNOR2_X1 U511 ( .A(KEYINPUT101), .B(n456), .ZN(n486) );
  NOR2_X1 U512 ( .A1(n486), .A2(n457), .ZN(n458) );
  XOR2_X1 U513 ( .A(KEYINPUT38), .B(n458), .Z(n467) );
  NOR2_X1 U514 ( .A1(n467), .A2(n545), .ZN(n460) );
  XNOR2_X1 U515 ( .A(KEYINPUT102), .B(KEYINPUT39), .ZN(n459) );
  XNOR2_X1 U516 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U517 ( .A(G29GAT), .B(n461), .ZN(G1328GAT) );
  NOR2_X1 U518 ( .A1(n467), .A2(n540), .ZN(n462) );
  XOR2_X1 U519 ( .A(G36GAT), .B(n462), .Z(G1329GAT) );
  XOR2_X1 U520 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n464) );
  XNOR2_X1 U521 ( .A(G43GAT), .B(KEYINPUT104), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n464), .B(n463), .ZN(n466) );
  NOR2_X1 U523 ( .A1(n467), .A2(n550), .ZN(n465) );
  XOR2_X1 U524 ( .A(n466), .B(n465), .Z(G1330GAT) );
  XNOR2_X1 U525 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n469) );
  NOR2_X1 U526 ( .A1(n495), .A2(n467), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n469), .B(n468), .ZN(G1331GAT) );
  XNOR2_X1 U528 ( .A(KEYINPUT65), .B(KEYINPUT41), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n470), .B(n571), .ZN(n528) );
  XNOR2_X1 U530 ( .A(KEYINPUT107), .B(n528), .ZN(n553) );
  NAND2_X1 U531 ( .A1(n567), .A2(n553), .ZN(n485) );
  INV_X1 U532 ( .A(n485), .ZN(n472) );
  NAND2_X1 U533 ( .A1(n472), .A2(n471), .ZN(n481) );
  NOR2_X1 U534 ( .A1(n481), .A2(n545), .ZN(n476) );
  XOR2_X1 U535 ( .A(KEYINPUT106), .B(KEYINPUT108), .Z(n474) );
  XNOR2_X1 U536 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n473) );
  XNOR2_X1 U537 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U538 ( .A(n476), .B(n475), .ZN(G1332GAT) );
  NOR2_X1 U539 ( .A1(n540), .A2(n481), .ZN(n478) );
  XNOR2_X1 U540 ( .A(G64GAT), .B(KEYINPUT109), .ZN(n477) );
  XNOR2_X1 U541 ( .A(n478), .B(n477), .ZN(G1333GAT) );
  NOR2_X1 U542 ( .A1(n550), .A2(n481), .ZN(n479) );
  XOR2_X1 U543 ( .A(KEYINPUT110), .B(n479), .Z(n480) );
  XNOR2_X1 U544 ( .A(G71GAT), .B(n480), .ZN(G1334GAT) );
  NOR2_X1 U545 ( .A1(n495), .A2(n481), .ZN(n483) );
  XNOR2_X1 U546 ( .A(KEYINPUT111), .B(KEYINPUT43), .ZN(n482) );
  XNOR2_X1 U547 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U548 ( .A(G78GAT), .B(n484), .Z(G1335GAT) );
  NOR2_X1 U549 ( .A1(n486), .A2(n485), .ZN(n487) );
  XOR2_X1 U550 ( .A(KEYINPUT112), .B(n487), .Z(n494) );
  NOR2_X1 U551 ( .A1(n494), .A2(n545), .ZN(n488) );
  XOR2_X1 U552 ( .A(G85GAT), .B(n488), .Z(G1336GAT) );
  NOR2_X1 U553 ( .A1(n494), .A2(n540), .ZN(n490) );
  XNOR2_X1 U554 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n489) );
  XNOR2_X1 U555 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U556 ( .A(G92GAT), .B(n491), .ZN(G1337GAT) );
  NOR2_X1 U557 ( .A1(n494), .A2(n550), .ZN(n493) );
  XNOR2_X1 U558 ( .A(G99GAT), .B(KEYINPUT115), .ZN(n492) );
  XNOR2_X1 U559 ( .A(n493), .B(n492), .ZN(G1338GAT) );
  XNOR2_X1 U560 ( .A(KEYINPUT44), .B(KEYINPUT116), .ZN(n497) );
  NOR2_X1 U561 ( .A1(n495), .A2(n494), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U563 ( .A(G106GAT), .B(n498), .Z(G1339GAT) );
  NOR2_X1 U564 ( .A1(n567), .A2(n528), .ZN(n500) );
  XNOR2_X1 U565 ( .A(KEYINPUT117), .B(KEYINPUT46), .ZN(n499) );
  XNOR2_X1 U566 ( .A(n500), .B(n499), .ZN(n502) );
  INV_X1 U567 ( .A(n538), .ZN(n561) );
  NOR2_X1 U568 ( .A1(n561), .A2(n557), .ZN(n501) );
  NAND2_X1 U569 ( .A1(n502), .A2(n501), .ZN(n503) );
  XNOR2_X1 U570 ( .A(n503), .B(KEYINPUT47), .ZN(n508) );
  NOR2_X1 U571 ( .A1(n575), .A2(n578), .ZN(n504) );
  XNOR2_X1 U572 ( .A(n504), .B(KEYINPUT45), .ZN(n505) );
  NAND2_X1 U573 ( .A1(n505), .A2(n571), .ZN(n506) );
  NOR2_X1 U574 ( .A1(n506), .A2(n551), .ZN(n507) );
  NOR2_X1 U575 ( .A1(n508), .A2(n507), .ZN(n509) );
  XOR2_X1 U576 ( .A(n509), .B(KEYINPUT64), .Z(n510) );
  XNOR2_X1 U577 ( .A(KEYINPUT48), .B(n510), .ZN(n541) );
  NAND2_X1 U578 ( .A1(n511), .A2(n541), .ZN(n512) );
  NOR2_X1 U579 ( .A1(n513), .A2(n512), .ZN(n520) );
  NAND2_X1 U580 ( .A1(n520), .A2(n551), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n514), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U582 ( .A(G120GAT), .B(KEYINPUT49), .Z(n516) );
  NAND2_X1 U583 ( .A1(n520), .A2(n553), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n516), .B(n515), .ZN(G1341GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n518) );
  NAND2_X1 U586 ( .A1(n520), .A2(n557), .ZN(n517) );
  XNOR2_X1 U587 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U588 ( .A(G127GAT), .B(n519), .Z(G1342GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n522) );
  NAND2_X1 U590 ( .A1(n520), .A2(n561), .ZN(n521) );
  XNOR2_X1 U591 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U592 ( .A(G134GAT), .B(n523), .Z(G1343GAT) );
  INV_X1 U593 ( .A(n541), .ZN(n524) );
  NOR2_X1 U594 ( .A1(n524), .A2(n545), .ZN(n525) );
  NAND2_X1 U595 ( .A1(n526), .A2(n525), .ZN(n537) );
  NOR2_X1 U596 ( .A1(n567), .A2(n537), .ZN(n527) );
  XOR2_X1 U597 ( .A(G141GAT), .B(n527), .Z(G1344GAT) );
  NOR2_X1 U598 ( .A1(n528), .A2(n537), .ZN(n533) );
  XOR2_X1 U599 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n530) );
  XNOR2_X1 U600 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n529) );
  XNOR2_X1 U601 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U602 ( .A(KEYINPUT52), .B(n531), .ZN(n532) );
  XNOR2_X1 U603 ( .A(n533), .B(n532), .ZN(G1345GAT) );
  NOR2_X1 U604 ( .A1(n575), .A2(n537), .ZN(n535) );
  XNOR2_X1 U605 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n534) );
  XNOR2_X1 U606 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U607 ( .A(G155GAT), .B(n536), .ZN(G1346GAT) );
  NOR2_X1 U608 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U609 ( .A(G162GAT), .B(n539), .Z(G1347GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT124), .B(n540), .Z(n542) );
  NAND2_X1 U611 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n543), .B(KEYINPUT125), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n544), .B(KEYINPUT54), .ZN(n546) );
  NAND2_X1 U614 ( .A1(n546), .A2(n545), .ZN(n564) );
  NOR2_X1 U615 ( .A1(n547), .A2(n564), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n548), .B(KEYINPUT55), .ZN(n549) );
  NOR2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n560), .A2(n551), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n552), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n555) );
  NAND2_X1 U621 ( .A1(n553), .A2(n560), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(n556), .ZN(G1349GAT) );
  NAND2_X1 U624 ( .A1(n557), .A2(n560), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(KEYINPUT126), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G183GAT), .B(n559), .ZN(G1350GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT58), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(n563), .ZN(G1351GAT) );
  INV_X1 U630 ( .A(n564), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n577) );
  NOR2_X1 U632 ( .A1(n567), .A2(n577), .ZN(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(n570), .ZN(G1352GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n577), .ZN(n573) );
  XNOR2_X1 U637 ( .A(KEYINPUT61), .B(KEYINPUT127), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(G204GAT), .B(n574), .Z(G1353GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n577), .ZN(n576) );
  XOR2_X1 U641 ( .A(G211GAT), .B(n576), .Z(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT62), .B(n579), .Z(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

