//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n812, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029;
  XNOR2_X1  g000(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G78gat), .B(G106gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G22gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(KEYINPUT84), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n209), .B1(new_n206), .B2(new_n205), .ZN(new_n210));
  NAND2_X1  g009(.A1(G228gat), .A2(G233gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT79), .B(G155gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G162gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT2), .ZN(new_n214));
  INV_X1    g013(.A(G141gat), .ZN(new_n215));
  INV_X1    g014(.A(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218));
  AND2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n217), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(KEYINPUT78), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT78), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G155gat), .B2(G162gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226));
  AND3_X1   g025(.A1(new_n223), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n217), .A2(new_n228), .A3(new_n218), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n214), .A2(new_n222), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G197gat), .B(G204gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT22), .ZN(new_n232));
  INV_X1    g031(.A(G211gat), .ZN(new_n233));
  INV_X1    g032(.A(G218gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G211gat), .B(G218gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n231), .A3(new_n235), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT29), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n230), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n239), .A2(KEYINPUT76), .A3(new_n240), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT76), .B1(new_n239), .B2(new_n240), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n229), .A2(new_n226), .A3(new_n223), .A4(new_n225), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n228), .B1(new_n212), .B2(G162gat), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n249), .B(new_n244), .C1(new_n250), .C2(new_n221), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n242), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT83), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n245), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n248), .A2(KEYINPUT83), .A3(new_n252), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n211), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n253), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n236), .A2(KEYINPUT82), .A3(new_n238), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n242), .B(new_n259), .C1(new_n241), .C2(KEYINPUT82), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n230), .B1(new_n260), .B2(new_n244), .ZN(new_n261));
  INV_X1    g060(.A(new_n211), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n258), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n210), .B1(new_n257), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n252), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT76), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n241), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n239), .A2(KEYINPUT76), .A3(new_n240), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n254), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n245), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n256), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(new_n262), .ZN(new_n273));
  OR3_X1    g072(.A1(new_n258), .A2(new_n261), .A3(new_n262), .ZN(new_n274));
  INV_X1    g073(.A(new_n210), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n264), .A2(new_n276), .A3(KEYINPUT85), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT85), .B1(new_n264), .B2(new_n276), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G226gat), .A2(G233gat), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g082(.A(KEYINPUT69), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT26), .ZN(new_n288));
  NOR2_X1   g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G183gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT27), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT27), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G183gat), .ZN(new_n297));
  INV_X1    g096(.A(G190gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n295), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n293), .B1(new_n299), .B2(KEYINPUT28), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT68), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(new_n296), .ZN(new_n302));
  NAND2_X1  g101(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(G183gat), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n295), .A2(KEYINPUT67), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT67), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n306), .A2(new_n294), .A3(KEYINPUT27), .ZN(new_n307));
  NOR2_X1   g106(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n304), .A2(new_n305), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n291), .A2(new_n300), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n298), .A3(KEYINPUT65), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT65), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(G183gat), .B2(G190gat), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT64), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n312), .A2(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AND3_X1   g116(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT24), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n292), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n318), .B1(new_n320), .B2(KEYINPUT64), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT66), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n317), .A2(new_n321), .A3(KEYINPUT66), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n289), .A2(KEYINPUT23), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT23), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n327), .B1(G169gat), .B2(G176gat), .ZN(new_n328));
  AND4_X1   g127(.A1(KEYINPUT25), .A2(new_n326), .A3(new_n286), .A4(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n326), .A2(new_n286), .A3(new_n328), .ZN(new_n331));
  NAND3_X1  g130(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n320), .B(new_n332), .C1(G183gat), .C2(G190gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT25), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n311), .B1(new_n330), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n280), .B1(new_n337), .B2(KEYINPUT29), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n325), .A2(new_n329), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT66), .B1(new_n317), .B2(new_n321), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n336), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n310), .A2(KEYINPUT70), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT70), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n291), .A2(new_n300), .A3(new_n309), .A4(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n341), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n346));
  INV_X1    g145(.A(new_n280), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n346), .B1(new_n345), .B2(new_n347), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n269), .B(new_n338), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G8gat), .B(G36gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(G64gat), .ZN(new_n352));
  INV_X1    g151(.A(G92gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n347), .A2(KEYINPUT29), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n345), .A2(new_n355), .B1(new_n337), .B2(new_n347), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n248), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n350), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT30), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n350), .A2(KEYINPUT30), .A3(new_n354), .A4(new_n357), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n350), .A2(new_n357), .ZN(new_n362));
  INV_X1    g161(.A(new_n354), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AND3_X1   g163(.A1(new_n360), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n221), .B1(new_n213), .B2(KEYINPUT2), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n223), .A2(new_n225), .A3(new_n226), .ZN(new_n367));
  INV_X1    g166(.A(new_n218), .ZN(new_n368));
  NOR2_X1   g167(.A1(G141gat), .A2(G148gat), .ZN(new_n369));
  NOR3_X1   g168(.A1(new_n368), .A2(new_n369), .A3(KEYINPUT2), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT3), .B1(new_n366), .B2(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(G127gat), .B(G134gat), .Z(new_n373));
  INV_X1    g172(.A(G120gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G113gat), .ZN(new_n375));
  INV_X1    g174(.A(G113gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(G120gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT71), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n375), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT1), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n378), .B1(new_n375), .B2(new_n377), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n373), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n373), .A2(KEYINPUT1), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT72), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n375), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n374), .A2(KEYINPUT72), .A3(G113gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n386), .A2(new_n377), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n383), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n372), .A2(new_n390), .A3(new_n251), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n230), .A2(KEYINPUT4), .A3(new_n383), .A4(new_n389), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n249), .B1(new_n250), .B2(new_n221), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G225gat), .A2(G233gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n391), .B(new_n392), .C1(new_n394), .C2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n390), .B(new_n230), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n399), .B(KEYINPUT5), .C1(new_n395), .C2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n397), .B1(new_n390), .B2(new_n393), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n396), .A2(KEYINPUT5), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n402), .A2(new_n391), .A3(new_n392), .A4(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT80), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n404), .A2(new_n405), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n401), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G1gat), .B(G29gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(KEYINPUT0), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(G57gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(G85gat), .ZN(new_n412));
  INV_X1    g211(.A(G57gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n410), .B(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(G85gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n408), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT6), .ZN(new_n419));
  INV_X1    g218(.A(new_n417), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n401), .B(new_n420), .C1(new_n406), .C2(new_n407), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n418), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n408), .A2(KEYINPUT6), .A3(new_n417), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n279), .B1(new_n365), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n264), .A2(new_n276), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT86), .B1(new_n412), .B2(new_n416), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n416), .A3(KEYINPUT86), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n402), .A2(new_n391), .A3(new_n392), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT87), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n432), .A3(new_n396), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n432), .B1(new_n431), .B2(new_n396), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT39), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n437), .B1(new_n400), .B2(new_n395), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n430), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n437), .B1(new_n434), .B2(new_n435), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT40), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n431), .A2(new_n396), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT87), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n443), .A2(new_n438), .A3(new_n433), .ZN(new_n444));
  INV_X1    g243(.A(new_n429), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n445), .A2(new_n427), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n440), .A2(new_n444), .A3(KEYINPUT40), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n408), .A2(new_n430), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n441), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n360), .A2(new_n361), .A3(new_n364), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n426), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(KEYINPUT88), .B(KEYINPUT38), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n362), .A2(new_n354), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n453), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n248), .B(new_n338), .C1(new_n348), .C2(new_n349), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT37), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n457), .B1(new_n356), .B2(new_n269), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n455), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n350), .A2(new_n457), .A3(new_n357), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n454), .B1(new_n461), .B2(new_n354), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n423), .A2(KEYINPUT89), .ZN(new_n463));
  OR2_X1    g262(.A1(new_n404), .A2(new_n405), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n404), .A2(new_n405), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT5), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n390), .B(new_n393), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n466), .B1(new_n467), .B2(new_n396), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n464), .A2(new_n465), .B1(new_n468), .B2(new_n399), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n421), .B(new_n419), .C1(new_n469), .C2(new_n446), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT89), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n408), .A2(new_n471), .A3(KEYINPUT6), .A4(new_n417), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n463), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n460), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n457), .B1(new_n350), .B2(new_n357), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n455), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n462), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n425), .B1(new_n452), .B2(new_n477), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n383), .A2(new_n389), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT25), .B1(new_n331), .B2(new_n333), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n325), .A2(new_n329), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n480), .B1(new_n481), .B2(new_n324), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n342), .A2(new_n344), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n479), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(G227gat), .A2(G233gat), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n341), .A2(new_n390), .A3(new_n342), .A4(new_n344), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  XOR2_X1   g287(.A(G71gat), .B(G99gat), .Z(new_n489));
  XNOR2_X1  g288(.A(G15gat), .B(G43gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT33), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n488), .A2(KEYINPUT32), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT73), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT73), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n488), .A2(new_n495), .A3(KEYINPUT32), .A4(new_n492), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n488), .A2(KEYINPUT32), .ZN(new_n498));
  INV_X1    g297(.A(new_n488), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n498), .B(new_n491), .C1(new_n499), .C2(KEYINPUT33), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n487), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n485), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT34), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(KEYINPUT74), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n486), .B1(new_n484), .B2(new_n487), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT74), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT34), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n501), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT75), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n497), .A2(new_n509), .A3(new_n500), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT36), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n497), .A2(new_n509), .A3(new_n500), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT75), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n511), .A2(KEYINPUT36), .A3(new_n513), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n478), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n463), .A2(new_n470), .A3(new_n472), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n451), .A2(KEYINPUT35), .A3(new_n426), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n509), .B1(new_n497), .B2(new_n500), .ZN(new_n524));
  NOR3_X1   g323(.A1(new_n516), .A2(new_n524), .A3(KEYINPUT75), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n513), .A2(new_n512), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n522), .B(new_n523), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n426), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n513), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n365), .A2(new_n424), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT35), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n521), .A2(KEYINPUT90), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT90), .B1(new_n521), .B2(new_n532), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G43gat), .B(G50gat), .ZN(new_n536));
  INV_X1    g335(.A(G29gat), .ZN(new_n537));
  INV_X1    g336(.A(G36gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT14), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT14), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(G29gat), .B2(G36gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT92), .ZN(new_n543));
  OAI22_X1  g342(.A1(new_n542), .A2(new_n543), .B1(new_n537), .B2(new_n538), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT92), .B1(new_n539), .B2(new_n541), .ZN(new_n545));
  OAI211_X1 g344(.A(KEYINPUT15), .B(new_n536), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n536), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n547));
  INV_X1    g346(.A(new_n542), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n547), .B(new_n548), .C1(KEYINPUT15), .C2(new_n536), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n546), .A2(new_n549), .A3(KEYINPUT17), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT17), .B1(new_n546), .B2(new_n549), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT95), .ZN(new_n553));
  XNOR2_X1  g352(.A(G15gat), .B(G22gat), .ZN(new_n554));
  INV_X1    g353(.A(G1gat), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(KEYINPUT93), .A3(KEYINPUT16), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT93), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT16), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n558), .B1(new_n559), .B2(G1gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n554), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT94), .ZN(new_n562));
  INV_X1    g361(.A(G8gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n556), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n562), .A2(new_n563), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n566), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n556), .A2(new_n568), .A3(new_n561), .A4(new_n564), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n552), .A2(new_n553), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n546), .A2(new_n549), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n546), .A2(new_n549), .A3(KEYINPUT17), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(new_n575), .A3(new_n570), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT95), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT18), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n570), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n567), .A2(KEYINPUT96), .A3(new_n569), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n583), .B1(new_n587), .B2(new_n572), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n578), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT97), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT97), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n578), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n579), .B(KEYINPUT13), .Z(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n587), .A2(new_n572), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n585), .A2(new_n546), .A3(new_n549), .A4(new_n586), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n578), .A2(new_n579), .A3(new_n596), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(new_n599), .B2(new_n581), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n593), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G169gat), .B(G197gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(G113gat), .B(G141gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n599), .A2(new_n581), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n607), .B1(new_n608), .B2(KEYINPUT98), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n601), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT98), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n611), .B1(new_n599), .B2(new_n581), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n593), .B(new_n600), .C1(new_n612), .C2(new_n607), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n610), .A2(KEYINPUT99), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT99), .B1(new_n610), .B2(new_n613), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n587), .ZN(new_n618));
  OR2_X1    g417(.A1(G57gat), .A2(G64gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(G57gat), .A2(G64gat), .ZN(new_n620));
  AND2_X1   g419(.A1(G71gat), .A2(G78gat), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(KEYINPUT9), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G71gat), .B(G78gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n624), .B(new_n625), .Z(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT21), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n618), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(G183gat), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n618), .A2(new_n294), .A3(new_n627), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n632));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n632), .B(new_n633), .Z(new_n634));
  OR2_X1    g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n626), .A2(KEYINPUT21), .ZN(new_n638));
  XNOR2_X1  g437(.A(G127gat), .B(G155gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G211gat), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n635), .A2(new_n641), .A3(new_n636), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(G85gat), .A2(G92gat), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(KEYINPUT7), .ZN(new_n648));
  NAND2_X1  g447(.A1(G85gat), .A2(G92gat), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(G99gat), .ZN(new_n651));
  INV_X1    g450(.A(G106gat), .ZN(new_n652));
  OAI21_X1  g451(.A(KEYINPUT8), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n650), .B(new_n653), .C1(new_n649), .C2(new_n648), .ZN(new_n654));
  XOR2_X1   g453(.A(G99gat), .B(G106gat), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n552), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n654), .A2(new_n655), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AND2_X1   g459(.A1(G232gat), .A2(G233gat), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n660), .A2(new_n572), .B1(KEYINPUT41), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n657), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G134gat), .B(G162gat), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n663), .B(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n661), .A2(KEYINPUT41), .ZN(new_n667));
  XNOR2_X1  g466(.A(G190gat), .B(G218gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n666), .B(new_n669), .Z(new_n670));
  AND2_X1   g469(.A1(new_n645), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n626), .A2(new_n660), .A3(KEYINPUT10), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n626), .A2(new_n660), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n624), .B(new_n625), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n656), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n672), .B1(new_n676), .B2(KEYINPUT10), .ZN(new_n677));
  NAND2_X1  g476(.A1(G230gat), .A2(G233gat), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n678), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(G120gat), .B(G148gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G176gat), .ZN(new_n683));
  INV_X1    g482(.A(G204gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n679), .A2(new_n681), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n679), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n677), .A2(KEYINPUT102), .A3(new_n678), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n681), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n686), .B1(new_n692), .B2(new_n685), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n671), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n535), .A2(new_n617), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT103), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n424), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n422), .A2(KEYINPUT104), .A3(new_n423), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g504(.A(KEYINPUT105), .B(KEYINPUT16), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(new_n563), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n698), .A2(new_n451), .A3(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n698), .A2(new_n451), .ZN(new_n710));
  AOI22_X1  g509(.A1(new_n708), .A2(new_n709), .B1(new_n710), .B2(G8gat), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(new_n709), .B2(new_n708), .ZN(G1325gat));
  INV_X1    g511(.A(new_n698), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n525), .A2(new_n526), .ZN(new_n714));
  OR3_X1    g513(.A1(new_n713), .A2(G15gat), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(G15gat), .B1(new_n713), .B2(new_n520), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(G1326gat));
  INV_X1    g516(.A(new_n279), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n698), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(KEYINPUT43), .B(G22gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1327gat));
  NAND2_X1  g520(.A1(new_n521), .A2(new_n532), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT90), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n521), .A2(KEYINPUT90), .A3(new_n532), .ZN(new_n725));
  INV_X1    g524(.A(new_n645), .ZN(new_n726));
  INV_X1    g525(.A(new_n670), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n693), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n724), .A2(new_n725), .A3(new_n617), .A4(new_n729), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n730), .A2(G29gat), .A3(new_n702), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT45), .Z(new_n732));
  XOR2_X1   g531(.A(new_n645), .B(KEYINPUT106), .Z(new_n733));
  NAND2_X1  g532(.A1(new_n610), .A2(new_n613), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(new_n734), .A3(new_n694), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT44), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n426), .A2(KEYINPUT35), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n365), .A2(new_n522), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n740), .B1(new_n517), .B2(new_n514), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT35), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n516), .A2(new_n524), .A3(new_n426), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n451), .B1(new_n423), .B2(new_n422), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n738), .B1(new_n741), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n527), .A2(KEYINPUT107), .A3(new_n531), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n746), .A2(new_n521), .A3(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n746), .A2(new_n521), .A3(new_n747), .A4(KEYINPUT108), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n670), .A2(KEYINPUT44), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n735), .B1(new_n737), .B2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(G29gat), .B1(new_n755), .B2(new_n702), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n732), .A2(new_n756), .ZN(G1328gat));
  NOR2_X1   g556(.A1(new_n365), .A2(G36gat), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n730), .A2(KEYINPUT46), .A3(new_n759), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT110), .Z(new_n761));
  OAI21_X1  g560(.A(KEYINPUT46), .B1(new_n730), .B2(new_n759), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT109), .ZN(new_n763));
  OAI21_X1  g562(.A(G36gat), .B1(new_n755), .B2(new_n365), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n761), .A2(new_n763), .A3(new_n764), .ZN(G1329gat));
  NOR3_X1   g564(.A1(new_n730), .A2(G43gat), .A3(new_n714), .ZN(new_n766));
  INV_X1    g565(.A(new_n520), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n754), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n766), .B1(new_n768), .B2(G43gat), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g569(.A(KEYINPUT48), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n533), .A2(new_n534), .A3(new_n670), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n753), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n735), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(new_n426), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G50gat), .ZN(new_n777));
  INV_X1    g576(.A(G50gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n718), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n730), .B2(KEYINPUT111), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n535), .A2(new_n781), .A3(new_n617), .A4(new_n729), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n771), .B1(new_n777), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n778), .B1(new_n754), .B2(new_n718), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n771), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT112), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  AOI211_X1 g587(.A(new_n279), .B(new_n735), .C1(new_n737), .C2(new_n753), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n771), .B(new_n783), .C1(new_n789), .C2(new_n778), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n776), .A2(G50gat), .B1(new_n782), .B2(new_n780), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n790), .B(new_n791), .C1(new_n771), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n788), .A2(new_n793), .ZN(G1331gat));
  AND2_X1   g593(.A1(new_n750), .A2(new_n751), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n694), .A2(new_n734), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n671), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n798), .A2(new_n702), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(new_n413), .ZN(G1332gat));
  XNOR2_X1  g599(.A(new_n451), .B(KEYINPUT113), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n804));
  AND2_X1   g603(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n803), .B2(new_n804), .ZN(G1333gat));
  OAI21_X1  g606(.A(G71gat), .B1(new_n798), .B2(new_n520), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n714), .A2(G71gat), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n808), .B1(new_n798), .B2(new_n809), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n810), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g610(.A1(new_n798), .A2(new_n279), .ZN(new_n812));
  XOR2_X1   g611(.A(new_n812), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g612(.A1(new_n728), .A2(new_n734), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n748), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT51), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n694), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(new_n415), .A3(new_n703), .ZN(new_n818));
  INV_X1    g617(.A(new_n774), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n796), .A2(new_n726), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n819), .A2(new_n702), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n818), .B1(new_n821), .B2(new_n415), .ZN(G1336gat));
  NOR2_X1   g621(.A1(new_n802), .A2(G92gat), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(new_n817), .B2(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n819), .A2(new_n802), .A3(new_n820), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n825), .B2(new_n353), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n819), .A2(new_n820), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n451), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n828), .A2(G92gat), .B1(new_n817), .B2(new_n823), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n826), .B1(new_n829), .B2(new_n830), .ZN(G1337gat));
  INV_X1    g630(.A(new_n714), .ZN(new_n832));
  AOI21_X1  g631(.A(G99gat), .B1(new_n817), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n520), .A2(new_n651), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n833), .B1(new_n827), .B2(new_n834), .ZN(G1338gat));
  NOR2_X1   g634(.A1(new_n528), .A2(G106gat), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT53), .B1(new_n817), .B2(new_n836), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n819), .A2(new_n528), .A3(new_n820), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n837), .B1(new_n838), .B2(new_n652), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n827), .A2(new_n718), .ZN(new_n840));
  AOI22_X1  g639(.A1(new_n840), .A2(G106gat), .B1(new_n817), .B2(new_n836), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(G1339gat));
  NOR2_X1   g642(.A1(new_n695), .A2(new_n734), .ZN(new_n844));
  XOR2_X1   g643(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n845));
  NAND3_X1  g644(.A1(new_n688), .A2(new_n689), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n847), .B1(new_n677), .B2(new_n678), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n672), .B(new_n680), .C1(new_n676), .C2(KEYINPUT10), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n685), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT55), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n846), .A2(KEYINPUT55), .A3(new_n850), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n853), .A2(new_n686), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n734), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n593), .A2(new_n607), .A3(new_n600), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT115), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n578), .A2(new_n596), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n596), .A2(new_n597), .ZN(new_n860));
  AOI22_X1  g659(.A1(new_n859), .A2(new_n580), .B1(new_n860), .B2(new_n595), .ZN(new_n861));
  INV_X1    g660(.A(new_n606), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n858), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n861), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(KEYINPUT115), .A3(new_n606), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n693), .A2(new_n857), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n856), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n670), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n865), .A2(new_n863), .A3(new_n857), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT116), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n727), .B(new_n855), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n844), .B1(new_n874), .B2(new_n733), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(new_n714), .A3(new_n718), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n801), .A2(new_n702), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n878), .A2(new_n376), .A3(new_n616), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n875), .A2(new_n702), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n743), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(new_n801), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n734), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n879), .B1(new_n883), .B2(new_n376), .ZN(G1340gat));
  NOR3_X1   g683(.A1(new_n878), .A2(new_n374), .A3(new_n694), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n882), .A2(new_n693), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(new_n374), .ZN(G1341gat));
  INV_X1    g686(.A(G127gat), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n882), .A2(new_n888), .A3(new_n645), .ZN(new_n889));
  OAI21_X1  g688(.A(G127gat), .B1(new_n878), .B2(new_n733), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT117), .ZN(G1342gat));
  NAND2_X1  g691(.A1(new_n727), .A2(new_n365), .ZN(new_n893));
  OR3_X1    g692(.A1(new_n881), .A2(G134gat), .A3(new_n893), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n894), .A2(KEYINPUT56), .ZN(new_n895));
  OAI21_X1  g694(.A(G134gat), .B1(new_n878), .B2(new_n670), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(KEYINPUT56), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G1343gat));
  NAND2_X1  g697(.A1(new_n520), .A2(new_n877), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n855), .A2(new_n727), .ZN(new_n900));
  INV_X1    g699(.A(new_n872), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n869), .A2(new_n870), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n727), .B1(new_n856), .B2(new_n866), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n733), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n844), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n426), .ZN(new_n908));
  XNOR2_X1  g707(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n855), .B1(new_n614), .B2(new_n615), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n727), .B1(new_n911), .B2(new_n866), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n726), .B1(new_n912), .B2(new_n903), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n906), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(KEYINPUT57), .A3(new_n718), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n899), .B1(new_n910), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n734), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n767), .A2(new_n528), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n880), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n919), .A2(new_n801), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n616), .A2(G141gat), .ZN(new_n921));
  AOI22_X1  g720(.A1(new_n917), .A2(G141gat), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT58), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n920), .A2(new_n921), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n923), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n215), .B1(new_n916), .B2(new_n617), .ZN(new_n926));
  OAI22_X1  g725(.A1(new_n922), .A2(new_n923), .B1(new_n925), .B2(new_n926), .ZN(G1344gat));
  NAND3_X1  g726(.A1(new_n920), .A2(new_n216), .A3(new_n693), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT59), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n696), .A2(new_n616), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n913), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n718), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT57), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n909), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n907), .A2(new_n426), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n694), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(new_n520), .A3(new_n877), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n929), .B1(new_n938), .B2(G148gat), .ZN(new_n939));
  AOI211_X1 g738(.A(KEYINPUT59), .B(new_n216), .C1(new_n916), .C2(new_n693), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n928), .B1(new_n939), .B2(new_n940), .ZN(G1345gat));
  INV_X1    g740(.A(new_n916), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n212), .B1(new_n942), .B2(new_n733), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n726), .A2(new_n212), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n920), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1346gat));
  OAI21_X1  g745(.A(G162gat), .B1(new_n942), .B2(new_n670), .ZN(new_n947));
  OR3_X1    g746(.A1(new_n919), .A2(G162gat), .A3(new_n893), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1347gat));
  NAND2_X1  g748(.A1(new_n801), .A2(new_n743), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT120), .ZN(new_n951));
  OAI21_X1  g750(.A(KEYINPUT119), .B1(new_n875), .B2(new_n703), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT119), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n907), .A2(new_n953), .A3(new_n702), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n951), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(G169gat), .B1(new_n955), .B2(new_n734), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n703), .A2(new_n365), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n876), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(G169gat), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n958), .A2(new_n959), .A3(new_n616), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n956), .A2(new_n960), .ZN(G1348gat));
  OAI21_X1  g760(.A(G176gat), .B1(new_n958), .B2(new_n694), .ZN(new_n962));
  INV_X1    g761(.A(new_n955), .ZN(new_n963));
  OR2_X1    g762(.A1(new_n694), .A2(G176gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(G1349gat));
  OAI21_X1  g764(.A(G183gat), .B1(new_n958), .B2(new_n733), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT121), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n645), .A2(new_n295), .A3(new_n297), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n955), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n967), .B1(new_n955), .B2(new_n968), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(KEYINPUT60), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT60), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n973), .B(new_n966), .C1(new_n969), .C2(new_n970), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n974), .ZN(G1350gat));
  OAI21_X1  g774(.A(G190gat), .B1(new_n958), .B2(new_n670), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT122), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT122), .ZN(new_n978));
  OAI211_X1 g777(.A(new_n978), .B(G190gat), .C1(new_n958), .C2(new_n670), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n977), .A2(KEYINPUT61), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n955), .A2(new_n298), .A3(new_n727), .ZN(new_n981));
  OAI211_X1 g780(.A(new_n980), .B(new_n981), .C1(KEYINPUT61), .C2(new_n977), .ZN(G1351gat));
  INV_X1    g781(.A(G197gat), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n279), .B1(new_n913), .B2(new_n930), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n936), .B1(KEYINPUT57), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n957), .A2(new_n520), .ZN(new_n986));
  XOR2_X1   g785(.A(new_n986), .B(KEYINPUT123), .Z(new_n987));
  NAND3_X1  g786(.A1(new_n985), .A2(new_n617), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n983), .B1(new_n988), .B2(KEYINPUT124), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n989), .B1(KEYINPUT124), .B2(new_n988), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n952), .A2(new_n954), .ZN(new_n991));
  NOR3_X1   g790(.A1(new_n767), .A2(new_n528), .A3(new_n802), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n993), .A2(new_n983), .A3(new_n734), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n990), .A2(new_n994), .ZN(G1352gat));
  NAND2_X1  g794(.A1(new_n937), .A2(new_n987), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(G204gat), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT125), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n694), .A2(G204gat), .ZN(new_n999));
  NOR3_X1   g798(.A1(new_n875), .A2(KEYINPUT119), .A3(new_n703), .ZN(new_n1000));
  AOI21_X1  g799(.A(new_n953), .B1(new_n907), .B2(new_n702), .ZN(new_n1001));
  OAI211_X1 g800(.A(new_n992), .B(new_n999), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1002), .A2(KEYINPUT62), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT62), .ZN(new_n1004));
  NAND4_X1  g803(.A1(new_n991), .A2(new_n1004), .A3(new_n992), .A4(new_n999), .ZN(new_n1005));
  NAND4_X1  g804(.A1(new_n997), .A2(new_n998), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1007));
  AOI21_X1  g806(.A(new_n684), .B1(new_n937), .B2(new_n987), .ZN(new_n1008));
  OAI21_X1  g807(.A(KEYINPUT125), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1006), .A2(new_n1009), .ZN(G1353gat));
  NAND3_X1  g809(.A1(new_n993), .A2(new_n233), .A3(new_n645), .ZN(new_n1011));
  AOI21_X1  g810(.A(KEYINPUT57), .B1(new_n931), .B2(new_n718), .ZN(new_n1012));
  AOI211_X1 g811(.A(new_n528), .B(new_n909), .C1(new_n905), .C2(new_n906), .ZN(new_n1013));
  OAI211_X1 g812(.A(new_n645), .B(new_n987), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  INV_X1    g813(.A(KEYINPUT126), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g815(.A1(new_n985), .A2(KEYINPUT126), .A3(new_n645), .A4(new_n987), .ZN(new_n1017));
  AND4_X1   g816(.A1(KEYINPUT63), .A2(new_n1016), .A3(G211gat), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g817(.A(new_n233), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1019));
  AOI21_X1  g818(.A(KEYINPUT63), .B1(new_n1019), .B2(new_n1017), .ZN(new_n1020));
  OAI21_X1  g819(.A(new_n1011), .B1(new_n1018), .B2(new_n1020), .ZN(G1354gat));
  NAND3_X1  g820(.A1(new_n991), .A2(new_n727), .A3(new_n992), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1022), .A2(new_n234), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n985), .A2(new_n987), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n727), .A2(G218gat), .ZN(new_n1025));
  OAI21_X1  g824(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1026), .A2(KEYINPUT127), .ZN(new_n1027));
  INV_X1    g826(.A(KEYINPUT127), .ZN(new_n1028));
  OAI211_X1 g827(.A(new_n1023), .B(new_n1028), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1027), .A2(new_n1029), .ZN(G1355gat));
endmodule


