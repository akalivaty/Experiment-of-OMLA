//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1332, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1401,
    new_n1402, new_n1403, new_n1404, new_n1405, new_n1406;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  OAI21_X1  g0008(.A(G50), .B1(G58), .B2(G68), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND3_X1  g0012(.A1(new_n210), .A2(G20), .A3(new_n212), .ZN(new_n213));
  XOR2_X1   g0013(.A(KEYINPUT64), .B(G77), .Z(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G116), .A2(G270), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n205), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n208), .B(new_n213), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0024(.A(G250), .B(G257), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT67), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(G270), .Z(new_n228));
  XNOR2_X1  g0028(.A(G226), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT66), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n228), .B(new_n234), .Z(G358));
  XNOR2_X1  g0035(.A(G87), .B(G97), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT68), .ZN(new_n237));
  INV_X1    g0037(.A(G107), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g0039(.A(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  INV_X1    g0045(.A(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G20), .ZN(new_n247));
  INV_X1    g0047(.A(G20), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G33), .ZN(new_n249));
  INV_X1    g0049(.A(G50), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  OAI221_X1 g0052(.A(new_n247), .B1(new_n249), .B2(new_n202), .C1(new_n250), .C2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n211), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n253), .A2(KEYINPUT11), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G13), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G1), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT12), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n256), .B1(KEYINPUT12), .B2(new_n259), .C1(new_n247), .C2(new_n262), .ZN(new_n263));
  AND3_X1   g0063(.A1(new_n258), .A2(new_n211), .A3(new_n254), .ZN(new_n264));
  OAI21_X1  g0064(.A(KEYINPUT72), .B1(new_n248), .B2(G1), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT72), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(new_n257), .A3(G20), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n246), .B1(new_n269), .B2(KEYINPUT12), .ZN(new_n270));
  AOI21_X1  g0070(.A(KEYINPUT11), .B1(new_n253), .B2(new_n255), .ZN(new_n271));
  OR3_X1    g0071(.A1(new_n263), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT14), .ZN(new_n273));
  INV_X1    g0073(.A(G169), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(KEYINPUT80), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT13), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  INV_X1    g0077(.A(G45), .ZN(new_n278));
  AOI21_X1  g0078(.A(G1), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(G1), .A3(G13), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(new_n281), .A3(G274), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT79), .ZN(new_n283));
  INV_X1    g0083(.A(G274), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n284), .B1(new_n212), .B2(new_n280), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT79), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(new_n286), .A3(new_n279), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n281), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n283), .A2(new_n287), .B1(G238), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G226), .A2(G1698), .ZN(new_n292));
  INV_X1    g0092(.A(G232), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(G1698), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT3), .B(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G97), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n281), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(KEYINPUT78), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n294), .A2(new_n295), .B1(G33), .B2(G97), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT78), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n300), .A2(new_n301), .A3(new_n281), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n276), .B(new_n291), .C1(new_n299), .C2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n298), .A2(KEYINPUT78), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n301), .B1(new_n300), .B2(new_n281), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n276), .B1(new_n307), .B2(new_n291), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n273), .B(new_n275), .C1(new_n304), .C2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n291), .B1(new_n299), .B2(new_n302), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT13), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n311), .A2(G179), .A3(new_n303), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n303), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n273), .B1(new_n314), .B2(new_n275), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n272), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n272), .B1(new_n314), .B2(G200), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n311), .A2(G190), .A3(new_n303), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n282), .B1(new_n293), .B2(new_n289), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n323));
  OR2_X1    g0123(.A1(G223), .A2(G1698), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT3), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G33), .ZN(new_n326));
  INV_X1    g0126(.A(G226), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G1698), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n323), .A2(new_n324), .A3(new_n326), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G33), .A2(G87), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n322), .A2(new_n333), .A3(G179), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n281), .B1(new_n329), .B2(new_n330), .ZN(new_n335));
  OAI21_X1  g0135(.A(G169), .B1(new_n321), .B2(new_n335), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n334), .A2(KEYINPUT83), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT83), .B1(new_n334), .B2(new_n336), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT8), .B(G58), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n259), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n254), .A2(new_n211), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(KEYINPUT71), .A3(new_n258), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT71), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n344), .B1(new_n259), .B2(new_n255), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n345), .A3(new_n268), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n341), .B1(new_n346), .B2(new_n340), .ZN(new_n347));
  INV_X1    g0147(.A(G58), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n348), .A2(new_n246), .ZN(new_n349));
  NOR2_X1   g0149(.A1(G58), .A2(G68), .ZN(new_n350));
  OAI21_X1  g0150(.A(G20), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(G20), .A2(G33), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n352), .A2(KEYINPUT81), .A3(G159), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT81), .B1(new_n352), .B2(G159), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n351), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT7), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n295), .B2(G20), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n323), .A2(new_n326), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n359), .A2(KEYINPUT7), .A3(new_n248), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n356), .B1(new_n361), .B2(G68), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n342), .B1(new_n362), .B2(KEYINPUT16), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT16), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT82), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n325), .B2(G33), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n251), .A2(KEYINPUT82), .A3(KEYINPUT3), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n326), .A3(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n357), .A2(G20), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n246), .B1(new_n370), .B2(new_n358), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n364), .B1(new_n371), .B2(new_n356), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n347), .B1(new_n363), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT18), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n339), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n334), .A2(new_n336), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT83), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n334), .A2(new_n336), .A3(KEYINPUT83), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n295), .A2(new_n357), .A3(G20), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT7), .B1(new_n359), .B2(new_n248), .ZN(new_n382));
  OAI21_X1  g0182(.A(G68), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n356), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(KEYINPUT16), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n372), .A2(new_n385), .A3(new_n255), .ZN(new_n386));
  INV_X1    g0186(.A(new_n347), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT18), .B1(new_n380), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT17), .ZN(new_n390));
  INV_X1    g0190(.A(G200), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(new_n322), .B2(new_n333), .ZN(new_n392));
  INV_X1    g0192(.A(G190), .ZN(new_n393));
  NOR3_X1   g0193(.A1(new_n321), .A2(new_n335), .A3(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n390), .B1(new_n373), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n386), .A2(new_n395), .A3(new_n387), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n397), .A2(KEYINPUT17), .ZN(new_n398));
  OAI22_X1  g0198(.A1(new_n375), .A2(new_n389), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n320), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G1698), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n295), .A2(G222), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT69), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n404), .B(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n359), .A2(new_n403), .ZN(new_n407));
  XNOR2_X1  g0207(.A(KEYINPUT64), .B(G77), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n407), .A2(G223), .B1(new_n408), .B2(new_n359), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n281), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n282), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(G226), .B2(new_n290), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n274), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g0214(.A(new_n404), .B(KEYINPUT69), .ZN(new_n415));
  INV_X1    g0215(.A(new_n409), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n332), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G179), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n418), .A3(new_n412), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n343), .A2(new_n345), .A3(G50), .A4(new_n268), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n259), .A2(new_n250), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n352), .A2(G150), .ZN(new_n424));
  OAI221_X1 g0224(.A(new_n424), .B1(new_n201), .B2(new_n248), .C1(new_n340), .C2(new_n249), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n255), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT70), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n426), .A2(KEYINPUT70), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n423), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n414), .A2(new_n419), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  OR2_X1    g0232(.A1(new_n426), .A2(KEYINPUT70), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n422), .B1(new_n433), .B2(new_n427), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT75), .B1(new_n434), .B2(KEYINPUT9), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT75), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT9), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n430), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(G200), .B1(new_n410), .B2(new_n413), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n423), .B(KEYINPUT9), .C1(new_n428), .C2(new_n429), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n417), .A2(G190), .A3(new_n412), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT76), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT10), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n439), .A2(new_n447), .A3(new_n443), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n432), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n295), .A2(G232), .A3(new_n403), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n238), .B2(new_n295), .ZN(new_n453));
  INV_X1    g0253(.A(G238), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n359), .A2(new_n454), .A3(new_n403), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n332), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n411), .B1(G244), .B2(new_n290), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G190), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT73), .ZN(new_n461));
  XOR2_X1   g0261(.A(KEYINPUT15), .B(G87), .Z(new_n462));
  INV_X1    g0262(.A(new_n249), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n462), .A2(new_n463), .B1(new_n408), .B2(G20), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n340), .A2(new_n252), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n342), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n264), .A2(G77), .A3(new_n268), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n214), .A2(new_n259), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n461), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT15), .B(G87), .ZN(new_n472));
  OAI22_X1  g0272(.A1(new_n214), .A2(new_n248), .B1(new_n472), .B2(new_n249), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n255), .B1(new_n473), .B2(new_n465), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n474), .A2(KEYINPUT73), .A3(new_n469), .A4(new_n468), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n458), .A2(G200), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n460), .A2(new_n471), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n471), .A2(new_n475), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n458), .A2(new_n274), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT74), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n471), .A2(new_n475), .B1(new_n458), .B2(new_n274), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n484), .A2(KEYINPUT74), .B1(new_n418), .B2(new_n459), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n478), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT77), .B1(new_n451), .B2(new_n486), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n439), .A2(new_n443), .A3(new_n447), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n447), .B1(new_n439), .B2(new_n443), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n431), .B(new_n486), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT77), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n402), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n258), .A2(G97), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n257), .A2(G33), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n258), .A2(new_n495), .A3(new_n211), .A4(new_n254), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n494), .B1(new_n497), .B2(G97), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n323), .A2(new_n326), .A3(G244), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(G1698), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n295), .A2(G244), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G283), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n501), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n295), .A2(G250), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n403), .B1(new_n506), .B2(KEYINPUT4), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n332), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n257), .B(G45), .C1(new_n277), .C2(KEYINPUT5), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n277), .A2(KEYINPUT5), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(new_n332), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n512), .A2(G257), .B1(new_n285), .B2(new_n511), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT86), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n393), .B1(new_n514), .B2(new_n391), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n508), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(G200), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n517), .B1(new_n508), .B2(new_n513), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT85), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n252), .A2(new_n202), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT6), .ZN(new_n522));
  INV_X1    g0322(.A(G97), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n523), .A2(new_n238), .ZN(new_n524));
  NOR2_X1   g0324(.A1(G97), .A2(G107), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n238), .A2(KEYINPUT6), .A3(G97), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n521), .B1(new_n528), .B2(G20), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n238), .B1(new_n370), .B2(new_n358), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT84), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n325), .A2(G33), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n248), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n357), .A2(new_n535), .B1(new_n368), .B2(new_n369), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n536), .A2(KEYINPUT84), .A3(new_n238), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n520), .B(new_n255), .C1(new_n532), .C2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(KEYINPUT84), .B1(new_n536), .B2(new_n238), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n370), .A2(new_n358), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(new_n531), .A3(G107), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n542), .A3(new_n529), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n520), .B1(new_n543), .B2(new_n255), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n498), .B(new_n519), .C1(new_n539), .C2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n498), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n255), .B1(new_n532), .B2(new_n537), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT85), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n546), .B1(new_n548), .B2(new_n538), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n274), .B1(new_n508), .B2(new_n513), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n508), .A2(new_n513), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n550), .B1(new_n552), .B2(G179), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n545), .B1(new_n549), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g0354(.A(KEYINPUT91), .B(KEYINPUT92), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT25), .ZN(new_n556));
  AOI211_X1 g0356(.A(G107), .B(new_n258), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n555), .A2(new_n556), .ZN(new_n558));
  XNOR2_X1  g0358(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n497), .A2(G107), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n323), .A2(new_n326), .A3(new_n248), .A4(G87), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT22), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT22), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n295), .A2(new_n565), .A3(new_n248), .A4(G87), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n248), .A2(KEYINPUT23), .A3(G107), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT23), .ZN(new_n569));
  OAI22_X1  g0369(.A1(new_n568), .A2(KEYINPUT89), .B1(new_n569), .B2(new_n238), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n238), .A3(G20), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT89), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n573));
  OAI22_X1  g0373(.A1(new_n571), .A2(new_n572), .B1(new_n573), .B2(G20), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n567), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT24), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT24), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n567), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT90), .B1(new_n580), .B2(new_n255), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n567), .A2(new_n575), .A3(new_n578), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n578), .B1(new_n567), .B2(new_n575), .ZN(new_n583));
  OAI211_X1 g0383(.A(KEYINPUT90), .B(new_n255), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n562), .B1(new_n581), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n295), .A2(G250), .A3(new_n403), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G33), .A2(G294), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n323), .A2(new_n326), .A3(G257), .A4(G1698), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n332), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n511), .A2(new_n285), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n512), .A2(G264), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n274), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(G179), .B2(new_n594), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n586), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n259), .A2(new_n240), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n496), .B2(new_n240), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n504), .B(new_n248), .C1(G33), .C2(new_n523), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n240), .A2(G20), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(new_n255), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT20), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n601), .A2(KEYINPUT20), .A3(new_n255), .A4(new_n602), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n600), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(G270), .B(new_n281), .C1(new_n509), .C2(new_n510), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n403), .A2(G257), .ZN(new_n609));
  NAND2_X1  g0409(.A1(G264), .A2(G1698), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n295), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n332), .B1(new_n295), .B2(G303), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n592), .B(new_n608), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n607), .A2(new_n614), .A3(new_n418), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(G200), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n617), .B(new_n607), .C1(new_n393), .C2(new_n614), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n614), .A2(G169), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n619), .A2(new_n607), .A3(KEYINPUT21), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT21), .ZN(new_n621));
  INV_X1    g0421(.A(new_n607), .ZN(new_n622));
  INV_X1    g0422(.A(G303), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n281), .B1(new_n359), .B2(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n624), .A2(new_n611), .B1(new_n285), .B2(new_n511), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n274), .B1(new_n625), .B2(new_n608), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n621), .B1(new_n622), .B2(new_n626), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n616), .B(new_n618), .C1(new_n620), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n454), .A2(new_n403), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n215), .A2(G1698), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n323), .A2(new_n629), .A3(new_n326), .A4(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n251), .A2(new_n240), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n281), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(G250), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n278), .B2(G1), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n257), .A2(new_n284), .A3(G45), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n281), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(G169), .B1(new_n634), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(G238), .A2(G1698), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n641), .B1(new_n215), .B2(G1698), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n632), .B1(new_n642), .B2(new_n295), .ZN(new_n643));
  OAI211_X1 g0443(.A(G179), .B(new_n638), .C1(new_n643), .C2(new_n281), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n462), .A2(new_n258), .ZN(new_n646));
  INV_X1    g0446(.A(G87), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n647), .A2(new_n523), .A3(new_n238), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n297), .A2(new_n248), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT19), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n323), .A2(new_n326), .A3(new_n248), .A4(G68), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT19), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n249), .B2(new_n523), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n646), .B1(new_n654), .B2(new_n255), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n497), .A2(new_n462), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n655), .A2(KEYINPUT87), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT87), .B1(new_n655), .B2(new_n656), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n645), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(G200), .B1(new_n634), .B2(new_n639), .ZN(new_n660));
  OAI211_X1 g0460(.A(G190), .B(new_n638), .C1(new_n643), .C2(new_n281), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT88), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n264), .A2(new_n662), .A3(G87), .A4(new_n495), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT88), .B1(new_n496), .B2(new_n647), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n660), .A2(new_n661), .A3(new_n655), .A4(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n659), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n628), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n255), .B1(new_n582), .B2(new_n583), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT90), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n584), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n594), .A2(new_n391), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n590), .A2(new_n332), .B1(new_n512), .B2(G264), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n674), .A2(new_n393), .A3(new_n592), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n672), .A2(new_n562), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n598), .A2(new_n668), .A3(new_n677), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n493), .A2(new_n554), .A3(new_n678), .ZN(G372));
  NAND3_X1  g0479(.A1(new_n388), .A2(new_n376), .A3(new_n374), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n374), .B1(new_n388), .B2(new_n376), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n479), .A2(new_n480), .A3(KEYINPUT74), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n459), .A2(new_n418), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n484), .A2(KEYINPUT74), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n319), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n689), .A2(new_n316), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n397), .A2(KEYINPUT17), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n373), .A2(new_n390), .A3(new_n395), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  OAI211_X1 g0494(.A(KEYINPUT96), .B(new_n683), .C1(new_n690), .C2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n449), .A2(new_n450), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT96), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n694), .B1(new_n689), .B2(new_n316), .ZN(new_n698));
  INV_X1    g0498(.A(new_n682), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n680), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n697), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n695), .A2(new_n696), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n431), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT93), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n645), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n640), .A2(new_n644), .A3(KEYINPUT93), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n706), .B(new_n707), .C1(new_n658), .C2(new_n657), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n660), .A2(new_n655), .A3(new_n665), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT94), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n660), .A2(new_n655), .A3(new_n665), .A4(KEYINPUT94), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(new_n661), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n561), .B1(new_n671), .B2(new_n584), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(new_n676), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT21), .B1(new_n619), .B2(new_n607), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n622), .A2(new_n626), .A3(new_n621), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n615), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n715), .B2(new_n596), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n498), .B1(new_n539), .B2(new_n544), .ZN(new_n721));
  INV_X1    g0521(.A(new_n553), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n716), .A2(new_n720), .A3(new_n723), .A4(new_n545), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n708), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT95), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n549), .A2(new_n714), .A3(new_n553), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n726), .B1(new_n727), .B2(KEYINPUT26), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT26), .ZN(new_n729));
  NOR4_X1   g0529(.A1(new_n549), .A2(new_n729), .A3(new_n667), .A4(new_n553), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n548), .A2(new_n538), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n553), .B1(new_n731), .B2(new_n498), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n708), .A2(new_n713), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT26), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n730), .B1(new_n734), .B2(KEYINPUT95), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n725), .B1(new_n728), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n704), .B1(new_n493), .B2(new_n736), .ZN(G369));
  NAND2_X1  g0537(.A1(new_n261), .A2(new_n248), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n738), .A2(KEYINPUT27), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(KEYINPUT27), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n739), .A2(G213), .A3(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G343), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n607), .ZN(new_n745));
  MUX2_X1   g0545(.A(new_n628), .B(new_n719), .S(new_n745), .Z(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT97), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n747), .A2(G330), .ZN(new_n748));
  AOI221_X4 g0548(.A(new_n561), .B1(new_n675), .B2(new_n673), .C1(new_n671), .C2(new_n584), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n596), .B1(new_n672), .B2(new_n562), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(new_n715), .B2(new_n744), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(new_n598), .B2(new_n744), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n719), .A2(new_n743), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n750), .A2(new_n744), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n754), .A2(new_n760), .ZN(G399));
  INV_X1    g0561(.A(new_n206), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G41), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n648), .A2(G116), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n763), .A2(new_n765), .A3(new_n257), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(new_n210), .B2(new_n763), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT98), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT28), .Z(new_n769));
  INV_X1    g0569(.A(new_n730), .ZN(new_n770));
  OAI211_X1 g0570(.A(KEYINPUT95), .B(new_n729), .C1(new_n723), .C2(new_n714), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n728), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n708), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n677), .A2(new_n733), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n554), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n773), .B1(new_n775), .B2(new_n720), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT29), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n777), .A2(new_n778), .A3(new_n744), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n723), .A2(new_n545), .A3(new_n677), .A4(new_n733), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n720), .A2(KEYINPUT101), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT101), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n782), .B(new_n719), .C1(new_n715), .C2(new_n596), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n780), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n667), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n732), .A2(new_n729), .A3(new_n785), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n786), .B(new_n708), .C1(new_n729), .C2(new_n727), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n744), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(KEYINPUT29), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n779), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G330), .ZN(new_n792));
  INV_X1    g0592(.A(new_n554), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n793), .A2(new_n751), .A3(new_n668), .A4(new_n744), .ZN(new_n794));
  OAI21_X1  g0594(.A(KEYINPUT99), .B1(new_n634), .B2(new_n639), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT99), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n796), .B(new_n638), .C1(new_n643), .C2(new_n281), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(G179), .B1(new_n625), .B2(new_n608), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT100), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n800), .A2(new_n801), .A3(new_n551), .A4(new_n594), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n798), .A2(new_n594), .A3(new_n799), .ZN(new_n803));
  OAI21_X1  g0603(.A(KEYINPUT100), .B1(new_n803), .B2(new_n552), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT30), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n614), .A2(new_n644), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n674), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n805), .B1(new_n807), .B2(new_n551), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n552), .A2(KEYINPUT30), .A3(new_n674), .A4(new_n806), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n802), .A2(new_n804), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n743), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT31), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n808), .B(new_n809), .C1(new_n552), .C2(new_n803), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n744), .A2(new_n812), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n811), .A2(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n792), .B1(new_n794), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n791), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n769), .B1(new_n819), .B2(G1), .ZN(G364));
  NOR2_X1   g0620(.A1(new_n260), .A2(G20), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(G45), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT102), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n823), .A2(new_n257), .A3(new_n763), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n748), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(G330), .B2(new_n747), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n393), .A2(G179), .A3(G200), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n248), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n523), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n248), .A2(new_n418), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n393), .A2(new_n391), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n359), .B(new_n829), .C1(G50), .C2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n830), .ZN(new_n835));
  NOR3_X1   g0635(.A1(new_n835), .A2(new_n391), .A3(G190), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n248), .A2(G179), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n831), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n836), .A2(G68), .B1(G87), .B2(new_n839), .ZN(new_n840));
  NOR3_X1   g0640(.A1(new_n835), .A2(new_n393), .A3(G200), .ZN(new_n841));
  NOR2_X1   g0641(.A1(G190), .A2(G200), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n830), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n841), .A2(G58), .B1(new_n408), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n834), .A2(new_n840), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n837), .A2(new_n393), .A3(G200), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT103), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(G107), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n837), .A2(new_n842), .ZN(new_n850));
  INV_X1    g0650(.A(G159), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT32), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n828), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n855), .A2(G294), .B1(new_n833), .B2(G326), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT104), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n848), .A2(G283), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n295), .B1(new_n839), .B2(G303), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n841), .A2(G322), .B1(G311), .B2(new_n844), .ZN(new_n860));
  XNOR2_X1  g0660(.A(KEYINPUT33), .B(G317), .ZN(new_n861));
  INV_X1    g0661(.A(new_n850), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n836), .A2(new_n861), .B1(G329), .B2(new_n862), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n858), .A2(new_n859), .A3(new_n860), .A4(new_n863), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n846), .A2(new_n854), .B1(new_n857), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n211), .B1(G20), .B2(new_n274), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n824), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n244), .A2(G45), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n762), .A2(new_n295), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n869), .B(new_n870), .C1(G45), .C2(new_n209), .ZN(new_n871));
  INV_X1    g0671(.A(G355), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n295), .A2(new_n206), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n871), .B1(G116), .B2(new_n206), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(G13), .A2(G33), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n876), .A2(G20), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n877), .A2(new_n866), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n868), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n877), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n867), .B(new_n879), .C1(new_n747), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n826), .A2(new_n881), .ZN(G396));
  INV_X1    g0682(.A(KEYINPUT108), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n777), .A2(new_n744), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n479), .A2(new_n743), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n477), .B(new_n885), .C1(new_n686), .C2(new_n687), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n485), .A2(new_n479), .A3(new_n483), .A4(new_n743), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n883), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n888), .ZN(new_n890));
  AOI211_X1 g0690(.A(KEYINPUT108), .B(new_n890), .C1(new_n777), .C2(new_n744), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n486), .A2(new_n744), .ZN(new_n892));
  OAI22_X1  g0692(.A1(new_n889), .A2(new_n891), .B1(new_n736), .B2(new_n892), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n893), .A2(new_n817), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n824), .B1(new_n893), .B2(new_n817), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n866), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n876), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n824), .B1(G77), .B2(new_n898), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n836), .A2(KEYINPUT105), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n836), .A2(KEYINPUT105), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(G283), .ZN(new_n904));
  OAI22_X1  g0704(.A1(new_n238), .A2(new_n838), .B1(new_n843), .B2(new_n240), .ZN(new_n905));
  INV_X1    g0705(.A(G311), .ZN(new_n906));
  OAI22_X1  g0706(.A1(new_n832), .A2(new_n623), .B1(new_n850), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  AOI211_X1 g0708(.A(new_n295), .B(new_n829), .C1(G294), .C2(new_n841), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n848), .A2(G87), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n904), .A2(new_n908), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n843), .A2(new_n851), .ZN(new_n912));
  INV_X1    g0712(.A(G143), .ZN(new_n913));
  INV_X1    g0713(.A(new_n841), .ZN(new_n914));
  INV_X1    g0714(.A(new_n836), .ZN(new_n915));
  INV_X1    g0715(.A(G150), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n913), .A2(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI211_X1 g0717(.A(new_n912), .B(new_n917), .C1(G137), .C2(new_n833), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT34), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n848), .A2(G68), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n855), .A2(G58), .B1(new_n839), .B2(G50), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(G132), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n295), .B1(new_n850), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT106), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n918), .B2(KEYINPUT34), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n911), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n899), .B1(new_n927), .B2(new_n866), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n890), .B2(new_n876), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT107), .Z(new_n930));
  OR2_X1    g0730(.A1(new_n896), .A2(new_n930), .ZN(G384));
  NOR3_X1   g0731(.A1(new_n211), .A2(new_n248), .A3(new_n240), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n528), .B(KEYINPUT109), .Z(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT35), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n935), .B2(new_n934), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT36), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n408), .B(new_n210), .C1(new_n348), .C2(new_n246), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n250), .A2(G68), .ZN(new_n940));
  AOI211_X1 g0740(.A(new_n257), .B(G13), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n246), .B1(new_n358), .B2(new_n360), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n364), .B1(new_n943), .B2(new_n356), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n385), .A2(new_n944), .A3(new_n255), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n387), .ZN(new_n946));
  INV_X1    g0746(.A(new_n741), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n399), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n946), .A2(new_n376), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n951), .A2(new_n948), .A3(new_n397), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT37), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n388), .B1(new_n380), .B2(new_n947), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT37), .B1(new_n373), .B2(new_n395), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n950), .A2(new_n957), .A3(KEYINPUT38), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT38), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n374), .B1(new_n339), .B2(new_n373), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n380), .A2(new_n388), .A3(KEYINPUT18), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n948), .B1(new_n962), .B2(new_n693), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n952), .A2(KEYINPUT37), .B1(new_n954), .B2(new_n955), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n959), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n958), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(KEYINPUT39), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT39), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n388), .A2(new_n376), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n388), .A2(new_n947), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n969), .A2(new_n970), .A3(new_n397), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n971), .A2(KEYINPUT37), .B1(new_n954), .B2(new_n955), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n693), .A2(KEYINPUT110), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT110), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n691), .A2(new_n692), .A3(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n973), .A2(new_n683), .A3(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n970), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n972), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n968), .B(new_n958), .C1(new_n978), .C2(KEYINPUT38), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n967), .A2(new_n979), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n272), .B(new_n744), .C1(new_n313), .C2(new_n315), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n272), .A2(new_n743), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n316), .A2(new_n319), .A3(new_n984), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n272), .B(new_n743), .C1(new_n313), .C2(new_n315), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n892), .B1(new_n772), .B2(new_n776), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n688), .A2(new_n744), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n966), .B(new_n987), .C1(new_n988), .C2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n700), .A2(new_n741), .ZN(new_n992));
  AND3_X1   g0792(.A1(new_n983), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n493), .B1(new_n789), .B2(new_n779), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n994), .A2(new_n703), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n993), .B(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n811), .A2(new_n812), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n810), .A2(KEYINPUT31), .A3(new_n743), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n794), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n888), .B1(new_n985), .B2(new_n986), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n966), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT40), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n958), .B1(new_n978), .B2(KEYINPUT38), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1004), .A2(KEYINPUT40), .A3(new_n999), .A4(new_n1000), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n678), .A2(new_n554), .A3(new_n743), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n997), .A2(new_n998), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1006), .B1(new_n493), .B2(new_n1009), .ZN(new_n1010));
  AND3_X1   g0810(.A1(new_n999), .A2(new_n1000), .A3(KEYINPUT40), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n1011), .A2(new_n1004), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n451), .A2(KEYINPUT77), .A3(new_n486), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n490), .A2(new_n491), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n401), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1012), .A2(new_n1015), .A3(new_n999), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1010), .A2(new_n1016), .A3(G330), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n996), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n257), .B2(new_n821), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n996), .A2(new_n1017), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n942), .B1(new_n1019), .B2(new_n1020), .ZN(G367));
  NAND2_X1  g0821(.A1(new_n732), .A2(new_n743), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT111), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT112), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n793), .B1(new_n549), .B2(new_n744), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1024), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n750), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n743), .B1(new_n1029), .B2(new_n723), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1032), .A2(new_n751), .A3(new_n756), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT42), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT43), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n655), .A2(new_n665), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n743), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n733), .A2(new_n1038), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n708), .A2(new_n1038), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1031), .A2(new_n1035), .A3(new_n1036), .A4(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1036), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1041), .A2(KEYINPUT43), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(new_n1030), .C2(new_n1034), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1047), .B1(new_n754), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1048), .A2(new_n754), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1043), .A2(new_n1050), .A3(new_n1046), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n763), .B(KEYINPUT41), .Z(new_n1052));
  INV_X1    g0852(.A(new_n754), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT44), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1032), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1054), .B1(new_n1055), .B2(new_n759), .ZN(new_n1056));
  NOR3_X1   g0856(.A1(new_n1032), .A2(KEYINPUT44), .A3(new_n760), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT45), .ZN(new_n1059));
  NOR3_X1   g0859(.A1(new_n1055), .A2(new_n1059), .A3(new_n759), .ZN(new_n1060));
  AOI21_X1  g0860(.A(KEYINPUT45), .B1(new_n1032), .B2(new_n760), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1053), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n757), .B1(new_n753), .B2(new_n756), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(new_n748), .Z(new_n1065));
  NOR2_X1   g0865(.A1(new_n818), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1067), .B(new_n754), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1063), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1052), .B1(new_n1069), .B2(new_n819), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n823), .A2(new_n257), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1049), .B(new_n1051), .C1(new_n1070), .C2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n870), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n228), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n878), .B1(new_n206), .B2(new_n472), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n824), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(G137), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n914), .A2(new_n916), .B1(new_n850), .B2(new_n1078), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n359), .B(new_n1079), .C1(G50), .C2(new_n844), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n855), .A2(G68), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n903), .A2(G159), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n214), .A2(new_n847), .B1(new_n838), .B2(new_n348), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G143), .B2(new_n833), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .A4(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n903), .A2(G294), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n839), .A2(G116), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT46), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n847), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n295), .B(new_n1089), .C1(G97), .C2(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1087), .A2(new_n1088), .B1(new_n855), .B2(G107), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n832), .A2(new_n906), .ZN(new_n1093));
  INV_X1    g0893(.A(G283), .ZN(new_n1094));
  INV_X1    g0894(.A(G317), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n843), .A2(new_n1094), .B1(new_n850), .B2(new_n1095), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1093), .B(new_n1096), .C1(G303), .C2(new_n841), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1086), .A2(new_n1091), .A3(new_n1092), .A4(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1085), .A2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT47), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1077), .B1(new_n1100), .B2(new_n866), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n1041), .B2(new_n880), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1073), .A2(new_n1102), .ZN(G387));
  INV_X1    g0903(.A(new_n1066), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n818), .A2(new_n1065), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1104), .A2(new_n763), .A3(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1065), .A2(new_n1071), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n753), .A2(new_n880), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n873), .A2(new_n764), .B1(G107), .B2(new_n206), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n234), .A2(G45), .ZN(new_n1110));
  AOI211_X1 g0910(.A(G45), .B(new_n765), .C1(G68), .C2(G77), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n340), .A2(G50), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT50), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1074), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1109), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n878), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n824), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G322), .A2(new_n833), .B1(new_n844), .B2(G303), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n1095), .B2(new_n914), .C1(new_n902), .C2(new_n906), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT48), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n855), .A2(G283), .B1(new_n839), .B2(G294), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT49), .ZN(new_n1125));
  OR2_X1    g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n847), .A2(new_n240), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n295), .B(new_n1128), .C1(G326), .C2(new_n862), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1126), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n214), .A2(new_n838), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n295), .B1(new_n850), .B2(new_n916), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1131), .B(new_n1132), .C1(new_n848), .C2(G97), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT113), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n828), .A2(new_n472), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n832), .A2(new_n851), .B1(new_n843), .B2(new_n246), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n250), .A2(new_n914), .B1(new_n915), .B2(new_n340), .ZN(new_n1137));
  NOR4_X1   g0937(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT114), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1130), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1117), .B1(new_n1140), .B2(new_n866), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1107), .B1(new_n1108), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1106), .A2(new_n1142), .ZN(G393));
  AOI22_X1  g0943(.A1(new_n841), .A2(G311), .B1(new_n833), .B2(G317), .ZN(new_n1144));
  XOR2_X1   g0944(.A(new_n1144), .B(KEYINPUT52), .Z(new_n1145));
  NAND2_X1  g0945(.A1(new_n903), .A2(G303), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n295), .B1(new_n862), .B2(G322), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n844), .A2(G294), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1147), .B(new_n1148), .C1(new_n1094), .C2(new_n838), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G116), .B2(new_n855), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1145), .A2(new_n1146), .A3(new_n849), .A4(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n841), .A2(G159), .B1(new_n833), .B2(G150), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT51), .Z(new_n1153));
  NAND2_X1  g0953(.A1(new_n903), .A2(G50), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n246), .A2(new_n838), .B1(new_n843), .B2(new_n340), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n828), .A2(new_n202), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n295), .B1(new_n850), .B2(new_n913), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1153), .A2(new_n1154), .A3(new_n910), .A4(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n897), .B1(new_n1151), .B2(new_n1159), .ZN(new_n1160));
  OR2_X1    g0960(.A1(new_n241), .A2(new_n1074), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1116), .B1(G97), .B2(new_n762), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n868), .B(new_n1160), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1048), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1163), .B1(new_n1164), .B2(new_n880), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1063), .A2(new_n1068), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n1071), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1069), .A2(new_n763), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1104), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(G390));
  NAND3_X1  g0971(.A1(new_n967), .A2(new_n979), .A3(new_n875), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n340), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n824), .B1(new_n1173), .B2(new_n898), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n832), .A2(new_n1094), .B1(new_n843), .B2(new_n523), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n914), .A2(new_n240), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(G294), .C2(new_n862), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n295), .B(new_n1156), .C1(G87), .C2(new_n839), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n903), .A2(G107), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n920), .A4(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n841), .A2(G132), .B1(new_n833), .B2(G128), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(KEYINPUT54), .B(G143), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n844), .A2(new_n1183), .B1(new_n862), .B2(G125), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1181), .B(new_n1184), .C1(new_n851), .C2(new_n828), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n295), .B1(new_n847), .B2(new_n250), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT118), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n838), .A2(new_n916), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT53), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1187), .B(new_n1189), .C1(new_n902), .C2(new_n1078), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1180), .B1(new_n1185), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1174), .B1(new_n1191), .B2(new_n866), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1172), .A2(new_n1192), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n999), .A2(new_n1000), .A3(G330), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n987), .B1(new_n988), .B2(new_n990), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n980), .B1(new_n1195), .B2(new_n981), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n981), .B(KEYINPUT115), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1004), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n989), .B1(new_n788), .B2(new_n888), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n1200), .B2(new_n987), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1194), .B1(new_n1196), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n974), .B1(new_n691), .B2(new_n692), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n700), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n970), .B1(new_n1204), .B2(new_n975), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n959), .B1(new_n1205), .B2(new_n972), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1197), .B1(new_n1206), .B2(new_n958), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n781), .A2(new_n783), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n775), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n729), .B1(new_n732), .B2(new_n733), .ZN(new_n1210));
  NOR4_X1   g1010(.A1(new_n549), .A2(KEYINPUT26), .A3(new_n667), .A4(new_n553), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1210), .A2(new_n1211), .A3(new_n773), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n743), .B1(new_n1209), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n990), .B1(new_n1213), .B2(new_n890), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n987), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1207), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n816), .A2(new_n1000), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n989), .B1(new_n736), .B2(new_n892), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n982), .B1(new_n1218), .B2(new_n987), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1216), .B(new_n1217), .C1(new_n1219), .C2(new_n980), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1202), .A2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1193), .B1(new_n1221), .B2(new_n1071), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n987), .B1(new_n816), .B2(new_n890), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1218), .B1(new_n1194), .B2(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(G330), .B(new_n890), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1225), .A2(new_n1215), .B1(new_n816), .B2(new_n1000), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT116), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1226), .A2(new_n1214), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1227), .B1(new_n1226), .B2(new_n1214), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1224), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1015), .A2(G330), .A3(new_n999), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n994), .A2(new_n1231), .A3(new_n703), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1230), .A2(new_n1202), .A3(new_n1220), .A4(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n763), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT117), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1234), .A2(new_n1235), .B1(new_n1221), .B2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1233), .A2(KEYINPUT117), .A3(new_n763), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1222), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(G378));
  NAND3_X1  g1040(.A1(new_n983), .A2(new_n991), .A3(new_n992), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n434), .A2(new_n741), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n451), .A2(new_n1245), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n432), .B(new_n1244), .C1(new_n449), .C2(new_n450), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1243), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n451), .A2(new_n1245), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n431), .B1(new_n488), .B2(new_n489), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1244), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(new_n1251), .A3(new_n1242), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1248), .A2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n1012), .B2(G330), .ZN(new_n1254));
  AND4_X1   g1054(.A1(G330), .A2(new_n1003), .A3(new_n1253), .A4(new_n1005), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1241), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1253), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n1006), .B2(new_n792), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1012), .A2(G330), .A3(new_n1253), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n993), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1256), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1257), .A2(new_n875), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n824), .B1(G50), .B2(new_n898), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n843), .A2(new_n472), .B1(new_n850), .B2(new_n1094), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n359), .A2(new_n277), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1264), .A2(new_n1131), .A3(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n847), .A2(new_n348), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(new_n841), .B2(G107), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n836), .A2(G97), .B1(new_n833), .B2(G116), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1266), .A2(new_n1081), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT58), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1265), .B(new_n250), .C1(G33), .C2(G41), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(G125), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n832), .A2(new_n1275), .B1(new_n843), .B2(new_n1078), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n841), .A2(G128), .B1(new_n839), .B2(new_n1183), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n916), .B2(new_n828), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1276), .B(new_n1278), .C1(G132), .C2(new_n836), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(KEYINPUT59), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1090), .A2(G159), .ZN(new_n1282));
  AOI211_X1 g1082(.A(G33), .B(G41), .C1(new_n862), .C2(G124), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1280), .A2(KEYINPUT59), .ZN(new_n1285));
  OAI221_X1 g1085(.A(new_n1274), .B1(new_n1271), .B2(new_n1270), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1263), .B1(new_n1286), .B2(new_n866), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1261), .A2(new_n1072), .B1(new_n1262), .B2(new_n1287), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(new_n1233), .A2(new_n1232), .B1(new_n1260), .B2(new_n1256), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n763), .B1(new_n1289), .B2(KEYINPUT57), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1224), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1229), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1226), .A2(new_n1214), .A3(new_n1227), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1291), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1232), .B1(new_n1221), .B2(new_n1294), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1295), .A2(KEYINPUT57), .A3(new_n1261), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1288), .B1(new_n1290), .B2(new_n1296), .ZN(G375));
  OR2_X1    g1097(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1052), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1236), .ZN(new_n1300));
  XOR2_X1   g1100(.A(new_n1300), .B(KEYINPUT119), .Z(new_n1301));
  AOI22_X1  g1101(.A1(G294), .A2(new_n833), .B1(new_n844), .B2(G107), .ZN(new_n1302));
  OAI221_X1 g1102(.A(new_n1302), .B1(new_n623), .B2(new_n850), .C1(new_n1094), .C2(new_n914), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n359), .B1(new_n838), .B2(new_n523), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(new_n1303), .A2(new_n1135), .A3(new_n1304), .ZN(new_n1305));
  AOI22_X1  g1105(.A1(new_n903), .A2(G116), .B1(G77), .B2(new_n848), .ZN(new_n1306));
  AOI22_X1  g1106(.A1(new_n841), .A2(G137), .B1(G150), .B2(new_n844), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1307), .B1(new_n923), .B2(new_n832), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1308), .B1(new_n903), .B2(new_n1183), .ZN(new_n1309));
  INV_X1    g1109(.A(G128), .ZN(new_n1310));
  OAI22_X1  g1110(.A1(new_n838), .A2(new_n851), .B1(new_n850), .B2(new_n1310), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n828), .A2(new_n250), .ZN(new_n1312));
  NOR4_X1   g1112(.A1(new_n1311), .A2(new_n1312), .A3(new_n1267), .A4(new_n359), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(new_n1305), .A2(new_n1306), .B1(new_n1309), .B2(new_n1313), .ZN(new_n1314));
  OAI221_X1 g1114(.A(new_n824), .B1(G68), .B2(new_n898), .C1(new_n1314), .C2(new_n897), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1315), .B1(new_n1215), .B2(new_n875), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1316), .B1(new_n1230), .B2(new_n1072), .ZN(new_n1317));
  AND2_X1   g1117(.A1(new_n1301), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(G381));
  INV_X1    g1119(.A(G396), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1106), .A2(new_n1142), .A3(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n896), .A2(new_n930), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(new_n1324), .B(KEYINPUT120), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1073), .A2(new_n1102), .A3(new_n1170), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1325), .A2(new_n1318), .A3(new_n1239), .A4(new_n1327), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1328), .A2(G375), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT121), .ZN(new_n1330));
  XNOR2_X1  g1130(.A(new_n1329), .B(new_n1330), .ZN(G407));
  NAND3_X1  g1131(.A1(new_n1239), .A2(G213), .A3(new_n742), .ZN(new_n1332));
  OAI211_X1 g1132(.A(G407), .B(G213), .C1(G375), .C2(new_n1332), .ZN(G409));
  INV_X1    g1133(.A(KEYINPUT125), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(G387), .A2(G390), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1320), .B1(new_n1106), .B2(new_n1142), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1322), .A2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  AND3_X1   g1138(.A1(new_n1335), .A2(new_n1338), .A3(new_n1326), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1338), .B1(new_n1335), .B2(new_n1326), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1334), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1335), .A2(new_n1326), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1337), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1335), .A2(new_n1338), .A3(new_n1326), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1343), .A2(KEYINPUT125), .A3(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1341), .A2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n742), .A2(G213), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT60), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1348), .B1(new_n1298), .B2(new_n1236), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1348), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1350), .A2(new_n763), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1317), .B1(new_n1349), .B2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1352), .A2(new_n1323), .ZN(new_n1353));
  OAI211_X1 g1153(.A(G384), .B(new_n1317), .C1(new_n1349), .C2(new_n1351), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1236), .A2(new_n1221), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1357), .A2(new_n1238), .A3(new_n1358), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1295), .A2(new_n1299), .A3(new_n1261), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1360), .A2(new_n1288), .ZN(new_n1361));
  INV_X1    g1161(.A(KEYINPUT122), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1222), .ZN(new_n1363));
  NAND4_X1  g1163(.A1(new_n1359), .A2(new_n1361), .A3(new_n1362), .A4(new_n1363), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1364), .B1(G375), .B2(new_n1239), .ZN(new_n1365));
  AOI21_X1  g1165(.A(new_n1362), .B1(new_n1239), .B2(new_n1361), .ZN(new_n1366));
  OAI211_X1 g1166(.A(new_n1347), .B(new_n1356), .C1(new_n1365), .C2(new_n1366), .ZN(new_n1367));
  XOR2_X1   g1167(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n1368));
  NAND2_X1  g1168(.A1(new_n1367), .A2(new_n1368), .ZN(new_n1369));
  AND3_X1   g1169(.A1(new_n1353), .A2(new_n1354), .A3(KEYINPUT62), .ZN(new_n1370));
  OAI211_X1 g1170(.A(new_n1347), .B(new_n1370), .C1(new_n1365), .C2(new_n1366), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1371), .A2(KEYINPUT124), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(new_n1359), .A2(new_n1361), .A3(new_n1363), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1373), .A2(KEYINPUT122), .ZN(new_n1374));
  OAI211_X1 g1174(.A(new_n1374), .B(new_n1364), .C1(new_n1239), .C2(G375), .ZN(new_n1375));
  INV_X1    g1175(.A(KEYINPUT124), .ZN(new_n1376));
  NAND4_X1  g1176(.A1(new_n1375), .A2(new_n1376), .A3(new_n1347), .A4(new_n1370), .ZN(new_n1377));
  NAND3_X1  g1177(.A1(new_n1369), .A2(new_n1372), .A3(new_n1377), .ZN(new_n1378));
  OAI21_X1  g1178(.A(new_n1347), .B1(new_n1365), .B2(new_n1366), .ZN(new_n1379));
  NAND3_X1  g1179(.A1(new_n742), .A2(G213), .A3(G2897), .ZN(new_n1380));
  AND3_X1   g1180(.A1(new_n1353), .A2(new_n1354), .A3(new_n1380), .ZN(new_n1381));
  AOI21_X1  g1181(.A(new_n1380), .B1(new_n1353), .B2(new_n1354), .ZN(new_n1382));
  NOR2_X1   g1182(.A1(new_n1381), .A2(new_n1382), .ZN(new_n1383));
  AOI21_X1  g1183(.A(KEYINPUT61), .B1(new_n1379), .B2(new_n1383), .ZN(new_n1384));
  AOI21_X1  g1184(.A(new_n1346), .B1(new_n1378), .B2(new_n1384), .ZN(new_n1385));
  INV_X1    g1185(.A(KEYINPUT63), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1367), .A2(new_n1386), .ZN(new_n1387));
  NOR2_X1   g1187(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1388));
  NAND4_X1  g1188(.A1(new_n1375), .A2(KEYINPUT63), .A3(new_n1347), .A4(new_n1356), .ZN(new_n1389));
  NAND4_X1  g1189(.A1(new_n1384), .A2(new_n1387), .A3(new_n1388), .A4(new_n1389), .ZN(new_n1390));
  INV_X1    g1190(.A(new_n1390), .ZN(new_n1391));
  OAI21_X1  g1191(.A(KEYINPUT126), .B1(new_n1385), .B2(new_n1391), .ZN(new_n1392));
  INV_X1    g1192(.A(KEYINPUT126), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(new_n1379), .A2(new_n1383), .ZN(new_n1394));
  INV_X1    g1194(.A(KEYINPUT61), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1394), .A2(new_n1395), .ZN(new_n1396));
  AOI22_X1  g1196(.A1(KEYINPUT124), .A2(new_n1371), .B1(new_n1367), .B2(new_n1368), .ZN(new_n1397));
  AOI21_X1  g1197(.A(new_n1396), .B1(new_n1397), .B2(new_n1377), .ZN(new_n1398));
  OAI211_X1 g1198(.A(new_n1393), .B(new_n1390), .C1(new_n1398), .C2(new_n1346), .ZN(new_n1399));
  NAND2_X1  g1199(.A1(new_n1392), .A2(new_n1399), .ZN(G405));
  INV_X1    g1200(.A(KEYINPUT127), .ZN(new_n1401));
  NAND3_X1  g1201(.A1(new_n1346), .A2(new_n1401), .A3(new_n1356), .ZN(new_n1402));
  XNOR2_X1  g1202(.A(G378), .B(G375), .ZN(new_n1403));
  OAI211_X1 g1203(.A(new_n1341), .B(new_n1345), .C1(KEYINPUT127), .C2(new_n1355), .ZN(new_n1404));
  AND3_X1   g1204(.A1(new_n1402), .A2(new_n1403), .A3(new_n1404), .ZN(new_n1405));
  AOI21_X1  g1205(.A(new_n1403), .B1(new_n1402), .B2(new_n1404), .ZN(new_n1406));
  NOR2_X1   g1206(.A1(new_n1405), .A2(new_n1406), .ZN(G402));
endmodule


