//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(KEYINPUT1), .B2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G120gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G113gat), .ZN(new_n206));
  INV_X1    g005(.A(G113gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G120gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G127gat), .B(G134gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n204), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(KEYINPUT24), .ZN(new_n215));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n214), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G183gat), .ZN(new_n219));
  INV_X1    g018(.A(G190gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(KEYINPUT24), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT24), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(KEYINPUT65), .ZN(new_n228));
  OAI211_X1 g027(.A(KEYINPUT66), .B(new_n216), .C1(new_n226), .C2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n218), .A2(new_n224), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n231));
  INV_X1    g030(.A(G169gat), .ZN(new_n232));
  INV_X1    g031(.A(G176gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT64), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(G169gat), .A3(G176gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n236), .A2(new_n241), .A3(KEYINPUT25), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n221), .B(new_n222), .C1(new_n217), .C2(KEYINPUT24), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(new_n241), .A3(new_n236), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT25), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n230), .A2(new_n243), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n241), .ZN(new_n248));
  NOR2_X1   g047(.A1(G169gat), .A2(G176gat), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT26), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n216), .B1(new_n248), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n219), .A2(KEYINPUT27), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT27), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G183gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n257), .A3(new_n220), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n258), .A2(new_n259), .A3(KEYINPUT28), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT28), .B1(new_n258), .B2(new_n259), .ZN(new_n261));
  NOR3_X1   g060(.A1(new_n254), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n213), .B1(new_n247), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n251), .A2(new_n252), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n217), .B1(new_n264), .B2(new_n241), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n258), .A2(new_n259), .A3(KEYINPUT28), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n258), .A2(new_n259), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT28), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n265), .A2(new_n266), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n213), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n216), .B1(new_n226), .B2(new_n228), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n223), .B1(new_n272), .B2(new_n214), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n242), .B1(new_n273), .B2(new_n229), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n245), .A2(new_n246), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n270), .B(new_n271), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n263), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G227gat), .A2(G233gat), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT32), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT33), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(G15gat), .B(G43gat), .Z(new_n284));
  XNOR2_X1  g083(.A(G71gat), .B(G99gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n281), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT34), .B1(new_n277), .B2(new_n279), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT34), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n263), .A2(new_n289), .A3(new_n276), .A4(new_n278), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT68), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n278), .B1(new_n263), .B2(new_n276), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n286), .B1(new_n294), .B2(KEYINPUT33), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT32), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n290), .A2(new_n291), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n287), .A2(new_n293), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(new_n288), .A3(new_n292), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n295), .A2(new_n297), .ZN(new_n302));
  AOI221_X4 g101(.A(new_n296), .B1(KEYINPUT33), .B2(new_n286), .C1(new_n277), .C2(new_n279), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n300), .A2(new_n304), .A3(KEYINPUT82), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT82), .B1(new_n300), .B2(new_n304), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G228gat), .A2(G233gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(G211gat), .B(G218gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G218gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT70), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT70), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G218gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT22), .B1(new_n316), .B2(G211gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(G197gat), .B(G204gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n311), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G211gat), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n321), .B1(new_n313), .B2(new_n315), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n318), .B(new_n310), .C1(new_n322), .C2(KEYINPUT22), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G141gat), .B(G148gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT2), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n329), .B1(G155gat), .B2(G162gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n327), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G141gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G148gat), .ZN(new_n333));
  INV_X1    g132(.A(G148gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(G141gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G155gat), .B(G162gat), .ZN(new_n337));
  INV_X1    g136(.A(G155gat), .ZN(new_n338));
  INV_X1    g137(.A(G162gat), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT2), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n336), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n331), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT73), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n331), .A2(new_n341), .A3(KEYINPUT73), .A4(new_n342), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT29), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n324), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n341), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n323), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT22), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT70), .B(G218gat), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n353), .B1(new_n354), .B2(new_n321), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n310), .B1(new_n355), .B2(new_n318), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n348), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n351), .B1(new_n357), .B2(new_n342), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n309), .B1(new_n349), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G22gat), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n331), .A2(new_n341), .A3(KEYINPUT72), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT72), .B1(new_n331), .B2(new_n341), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT29), .B1(new_n320), .B2(new_n323), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n363), .B1(new_n364), .B2(KEYINPUT3), .ZN(new_n365));
  INV_X1    g164(.A(new_n309), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT29), .B1(new_n345), .B2(new_n346), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n365), .B(new_n366), .C1(new_n324), .C2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n359), .A2(new_n360), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n359), .A2(new_n368), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G22gat), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n359), .A2(new_n368), .A3(KEYINPUT79), .A4(new_n360), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n371), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G78gat), .B(G106gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT31), .B(G50gat), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n376), .B(new_n377), .Z(new_n378));
  XOR2_X1   g177(.A(new_n378), .B(KEYINPUT78), .Z(new_n379));
  NAND2_X1  g178(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n378), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n373), .A2(new_n369), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n324), .ZN(new_n385));
  INV_X1    g184(.A(G226gat), .ZN(new_n386));
  INV_X1    g185(.A(G233gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n270), .B1(new_n274), .B2(new_n275), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n388), .B1(new_n389), .B2(new_n348), .ZN(new_n390));
  INV_X1    g189(.A(new_n388), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n230), .A2(new_n243), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n245), .A2(new_n246), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n391), .B1(new_n394), .B2(new_n270), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n385), .B1(new_n390), .B2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G8gat), .B(G36gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(G64gat), .B(G92gat), .ZN(new_n398));
  XOR2_X1   g197(.A(new_n397), .B(new_n398), .Z(new_n399));
  NAND2_X1  g198(.A1(new_n389), .A2(new_n388), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT29), .B1(new_n394), .B2(new_n270), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n400), .B(new_n324), .C1(new_n401), .C2(new_n388), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n396), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT71), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT30), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n396), .A2(new_n402), .A3(KEYINPUT71), .A4(new_n399), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n399), .B1(new_n396), .B2(new_n402), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n396), .A2(new_n399), .A3(new_n402), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n409), .B1(new_n410), .B2(KEYINPUT30), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n384), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT72), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n350), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n331), .A2(new_n341), .A3(KEYINPUT72), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(KEYINPUT3), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n347), .A2(new_n418), .A3(new_n213), .ZN(new_n419));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n204), .A2(new_n331), .A3(new_n341), .A4(new_n212), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(KEYINPUT4), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n419), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT75), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n416), .A2(new_n213), .A3(new_n417), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n421), .ZN(new_n428));
  INV_X1    g227(.A(new_n420), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n426), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  XOR2_X1   g230(.A(G1gat), .B(G29gat), .Z(new_n432));
  XNOR2_X1  g231(.A(G57gat), .B(G85gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n435));
  XOR2_X1   g234(.A(new_n434), .B(new_n435), .Z(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n427), .A2(new_n421), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n425), .B1(new_n438), .B2(new_n420), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n439), .A2(new_n423), .A3(KEYINPUT75), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT77), .B(KEYINPUT6), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n431), .A2(new_n437), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n431), .A2(new_n437), .A3(new_n440), .ZN(new_n444));
  INV_X1    g243(.A(new_n441), .ZN(new_n445));
  AND2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n440), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n439), .B1(KEYINPUT75), .B2(new_n423), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n436), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n443), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n450), .A2(KEYINPUT35), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n308), .A2(new_n413), .A3(new_n414), .A4(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n412), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n449), .A2(new_n444), .A3(new_n445), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n442), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT35), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n453), .A2(new_n455), .A3(new_n383), .A4(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT83), .B1(new_n457), .B2(new_n307), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n301), .B(KEYINPUT69), .C1(new_n302), .C2(new_n303), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT69), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n300), .A2(new_n304), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n384), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n450), .A2(new_n412), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT35), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT36), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n468), .B1(new_n462), .B2(new_n460), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT36), .B1(new_n300), .B2(new_n304), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n453), .A2(new_n455), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n470), .A2(new_n472), .B1(new_n384), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n420), .B1(new_n419), .B2(new_n422), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT39), .B1(new_n428), .B2(new_n429), .ZN(new_n476));
  OR2_X1    g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT39), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n477), .A2(KEYINPUT40), .A3(new_n436), .A4(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT40), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n436), .B1(new_n475), .B2(new_n476), .ZN(new_n482));
  AOI211_X1 g281(.A(KEYINPUT39), .B(new_n420), .C1(new_n419), .C2(new_n422), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n480), .A2(new_n444), .A3(new_n484), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n412), .A2(new_n485), .B1(new_n380), .B2(new_n382), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT81), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT80), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT37), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n396), .A2(new_n489), .A3(new_n402), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n489), .B1(new_n396), .B2(new_n402), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n490), .A2(new_n491), .A3(new_n399), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT38), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n488), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n491), .ZN(new_n495));
  INV_X1    g294(.A(new_n399), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n396), .A2(new_n489), .A3(new_n402), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n498), .A2(KEYINPUT80), .A3(KEYINPUT38), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n405), .A2(new_n407), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n495), .A2(new_n493), .A3(new_n496), .A4(new_n497), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n454), .A2(new_n502), .A3(new_n503), .A4(new_n442), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n486), .B(new_n487), .C1(new_n500), .C2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n501), .B1(new_n492), .B2(new_n493), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n450), .A2(new_n507), .A3(new_n494), .A4(new_n499), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n487), .B1(new_n508), .B2(new_n486), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n474), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n467), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G15gat), .B(G22gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT88), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(G8gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT16), .ZN(new_n517));
  AOI21_X1  g316(.A(G1gat), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n516), .B(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G43gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(G50gat), .ZN(new_n521));
  INV_X1    g320(.A(G50gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(G43gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT85), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT15), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n525), .B(new_n526), .C1(new_n524), .C2(new_n523), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT86), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n521), .A2(new_n523), .A3(KEYINPUT15), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G29gat), .ZN(new_n531));
  INV_X1    g330(.A(G36gat), .ZN(new_n532));
  OR3_X1    g331(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT84), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT84), .B1(new_n531), .B2(new_n532), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n535));
  OR3_X1    g334(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n533), .A2(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n530), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n537), .B1(new_n527), .B2(KEYINPUT86), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n529), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n519), .B1(KEYINPUT17), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT87), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n538), .A2(new_n540), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT17), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n541), .A2(KEYINPUT87), .A3(KEYINPUT17), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n542), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G229gat), .A2(G233gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n544), .A2(new_n519), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n548), .A2(KEYINPUT18), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n519), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n541), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n550), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n549), .B(KEYINPUT13), .Z(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n544), .A2(new_n543), .A3(new_n545), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT87), .B1(new_n541), .B2(KEYINPUT17), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n560), .A2(new_n542), .B1(new_n544), .B2(new_n519), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT18), .B1(new_n561), .B2(new_n549), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT89), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n551), .A2(new_n564), .A3(new_n556), .ZN(new_n565));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566));
  INV_X1    g365(.A(G197gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT11), .B(G169gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n570), .B(KEYINPUT12), .Z(new_n571));
  NAND2_X1  g370(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n563), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n565), .B(new_n571), .C1(new_n557), .C2(new_n562), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT99), .ZN(new_n577));
  NAND2_X1  g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578));
  INV_X1    g377(.A(G85gat), .ZN(new_n579));
  INV_X1    g378(.A(G92gat), .ZN(new_n580));
  AOI22_X1  g379(.A1(KEYINPUT8), .A2(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT97), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n584), .A2(G85gat), .A3(G92gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT7), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G99gat), .B(G106gat), .Z(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n588), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n583), .A2(new_n590), .A3(new_n586), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(G57gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n594), .A2(G64gat), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n594), .A2(G64gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT92), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n598), .B1(new_n597), .B2(new_n596), .ZN(new_n599));
  NAND2_X1  g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  OR2_X1    g399(.A1(G71gat), .A2(G78gat), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT9), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n600), .A2(new_n602), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n605), .B1(new_n596), .B2(new_n595), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n600), .B(KEYINPUT90), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n606), .A2(new_n607), .A3(new_n601), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n608), .A2(KEYINPUT91), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(KEYINPUT91), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n604), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n593), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT98), .B1(new_n592), .B2(new_n611), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n593), .A2(KEYINPUT98), .A3(new_n612), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G230gat), .A2(G233gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n613), .A2(KEYINPUT10), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n615), .A2(G230gat), .A3(G233gat), .A4(new_n616), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n624), .B(new_n625), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n577), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n621), .A2(KEYINPUT99), .A3(new_n622), .A4(new_n626), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n623), .A2(new_n627), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n634));
  NOR2_X1   g433(.A1(new_n612), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G127gat), .B(G155gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n519), .B1(new_n612), .B2(KEYINPUT21), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n637), .B(new_n638), .Z(new_n639));
  NAND2_X1  g438(.A1(G231gat), .A2(G233gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT94), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G183gat), .B(G211gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n639), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G232gat), .A2(G233gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n648), .A2(KEYINPUT41), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT95), .ZN(new_n650));
  XNOR2_X1  g449(.A(G134gat), .B(G162gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n593), .B1(KEYINPUT17), .B2(new_n541), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n560), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(G190gat), .B(G218gat), .Z(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AOI22_X1  g456(.A1(new_n544), .A2(new_n593), .B1(KEYINPUT41), .B2(new_n648), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n655), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n657), .B1(new_n655), .B2(new_n658), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n653), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n661), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n664), .A2(new_n652), .A3(new_n659), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n633), .A2(new_n646), .A3(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n512), .A2(new_n576), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n450), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G1gat), .ZN(G1324gat));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n669), .A2(new_n412), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT16), .B(G8gat), .Z(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n672), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n669), .A2(KEYINPUT42), .A3(new_n412), .A4(new_n674), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n673), .A2(G8gat), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(G1325gat));
  INV_X1    g478(.A(G15gat), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n669), .A2(new_n680), .A3(new_n308), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n470), .A2(new_n472), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT100), .Z(new_n683));
  NAND2_X1  g482(.A1(new_n669), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n681), .B1(new_n685), .B2(new_n680), .ZN(G1326gat));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n384), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT43), .B(G22gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  INV_X1    g488(.A(new_n667), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n576), .A2(new_n646), .A3(new_n632), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n511), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(G29gat), .A3(new_n455), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT45), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n691), .B(KEYINPUT101), .Z(new_n695));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n696));
  OAI22_X1  g495(.A1(new_n464), .A2(new_n383), .B1(new_n469), .B2(new_n471), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n486), .B1(new_n500), .B2(new_n504), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT81), .ZN(new_n699));
  AOI211_X1 g498(.A(new_n696), .B(new_n697), .C1(new_n699), .C2(new_n505), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n505), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT102), .B1(new_n701), .B2(new_n474), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n467), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n662), .A2(new_n665), .A3(KEYINPUT103), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT103), .B1(new_n662), .B2(new_n665), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n703), .A2(new_n704), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n704), .B1(new_n511), .B2(new_n690), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n695), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n531), .B1(new_n712), .B2(new_n450), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n694), .A2(new_n713), .ZN(G1328gat));
  NOR3_X1   g513(.A1(new_n692), .A2(G36gat), .A3(new_n453), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT46), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n712), .A2(new_n412), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n717), .B2(new_n532), .ZN(G1329gat));
  NOR3_X1   g517(.A1(new_n692), .A2(G43gat), .A3(new_n307), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n712), .A2(new_n683), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n719), .B1(new_n720), .B2(G43gat), .ZN(new_n721));
  INV_X1    g520(.A(new_n682), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n520), .B1(new_n712), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT47), .ZN(new_n724));
  OR2_X1    g523(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  OAI22_X1  g524(.A1(new_n721), .A2(KEYINPUT47), .B1(new_n723), .B2(new_n725), .ZN(G1330gat));
  NOR3_X1   g525(.A1(new_n692), .A2(G50gat), .A3(new_n383), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n384), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n727), .B1(new_n728), .B2(G50gat), .ZN(new_n729));
  XNOR2_X1  g528(.A(KEYINPUT104), .B(KEYINPUT48), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n729), .B(new_n730), .Z(G1331gat));
  AOI22_X1  g530(.A1(new_n452), .A2(new_n458), .B1(new_n465), .B2(KEYINPUT35), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n510), .A2(new_n696), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n701), .A2(KEYINPUT102), .A3(new_n474), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n576), .A2(new_n646), .A3(new_n667), .A4(new_n632), .ZN(new_n736));
  OR3_X1    g535(.A1(new_n735), .A2(KEYINPUT105), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT105), .B1(new_n735), .B2(new_n736), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n455), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(new_n594), .ZN(G1332gat));
  NOR2_X1   g540(.A1(new_n739), .A2(new_n453), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  AND2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n742), .B2(new_n743), .ZN(G1333gat));
  INV_X1    g545(.A(G71gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(new_n739), .B2(new_n307), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT106), .ZN(new_n749));
  INV_X1    g548(.A(new_n739), .ZN(new_n750));
  INV_X1    g549(.A(new_n683), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n747), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n749), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n752), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n739), .A2(KEYINPUT106), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n748), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g556(.A1(new_n750), .A2(new_n384), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G78gat), .ZN(G1335gat));
  OAI21_X1  g558(.A(KEYINPUT107), .B1(new_n735), .B2(new_n667), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT107), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n703), .A2(new_n761), .A3(new_n690), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n646), .A2(new_n575), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n760), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n760), .A2(new_n762), .A3(KEYINPUT51), .A4(new_n763), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n633), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(new_n579), .A3(new_n450), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n763), .A2(new_n632), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n707), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n705), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n735), .A2(KEYINPUT44), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n771), .B1(new_n774), .B2(new_n710), .ZN(new_n775));
  OAI21_X1  g574(.A(G85gat), .B1(new_n775), .B2(new_n455), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n769), .A2(new_n776), .ZN(G1336gat));
  NOR3_X1   g576(.A1(new_n633), .A2(G92gat), .A3(new_n453), .ZN(new_n778));
  INV_X1    g577(.A(new_n763), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n703), .A2(new_n690), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n779), .B1(new_n780), .B2(KEYINPUT107), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT51), .B1(new_n781), .B2(new_n762), .ZN(new_n782));
  INV_X1    g581(.A(new_n767), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n778), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n785));
  OAI21_X1  g584(.A(G92gat), .B1(new_n775), .B2(new_n453), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n778), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n788), .B1(new_n766), .B2(new_n767), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n770), .B1(new_n711), .B2(new_n709), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n580), .B1(new_n790), .B2(new_n412), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT109), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT52), .B1(new_n786), .B2(new_n793), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n787), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n794), .B1(new_n787), .B2(new_n792), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(G1337gat));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n798));
  XOR2_X1   g597(.A(KEYINPUT110), .B(G99gat), .Z(new_n799));
  NOR3_X1   g598(.A1(new_n775), .A2(new_n751), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n768), .A2(new_n308), .ZN(new_n802));
  INV_X1    g601(.A(new_n799), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n798), .B(new_n801), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n768), .B2(new_n308), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT111), .B1(new_n805), .B2(new_n800), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(G1338gat));
  OAI211_X1 g606(.A(new_n384), .B(new_n771), .C1(new_n774), .C2(new_n710), .ZN(new_n808));
  XOR2_X1   g607(.A(KEYINPUT112), .B(G106gat), .Z(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(KEYINPUT113), .A2(KEYINPUT53), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n383), .A2(G106gat), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n812), .B1(new_n768), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(KEYINPUT113), .A2(KEYINPUT53), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n814), .B(new_n815), .ZN(G1339gat));
  INV_X1    g615(.A(new_n646), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n618), .A2(new_n818), .A3(new_n619), .A4(new_n620), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n621), .A2(KEYINPUT54), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n619), .B1(new_n618), .B2(new_n620), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n627), .B(new_n819), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n822), .A2(new_n823), .B1(new_n628), .B2(new_n629), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n825), .B1(new_n822), .B2(new_n823), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n820), .A2(new_n821), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n819), .A2(new_n627), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n827), .A2(KEYINPUT114), .A3(KEYINPUT55), .A4(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n824), .A2(new_n575), .A3(new_n826), .A4(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n571), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n561), .A2(new_n549), .B1(new_n554), .B2(new_n555), .ZN(new_n832));
  AOI22_X1  g631(.A1(new_n563), .A2(new_n831), .B1(new_n570), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n632), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n708), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n824), .A2(new_n826), .A3(new_n829), .A4(new_n833), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(new_n773), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n817), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n668), .A2(new_n575), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n839), .B1(new_n838), .B2(new_n841), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n842), .A2(new_n843), .A3(new_n384), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n450), .A2(new_n453), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n307), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(G113gat), .A3(new_n575), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n842), .A2(new_n843), .A3(new_n455), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(KEYINPUT116), .A3(new_n463), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n838), .A2(new_n841), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT115), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n853), .A2(new_n450), .A3(new_n463), .A4(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI211_X1 g656(.A(new_n412), .B(new_n576), .C1(new_n851), .C2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n849), .B1(new_n858), .B2(G113gat), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g660(.A(KEYINPUT117), .B(new_n849), .C1(new_n858), .C2(G113gat), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1340gat));
  NAND3_X1  g662(.A1(new_n848), .A2(G120gat), .A3(new_n632), .ZN(new_n864));
  AOI211_X1 g663(.A(new_n412), .B(new_n633), .C1(new_n851), .C2(new_n857), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n865), .B2(G120gat), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT118), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n868), .B(new_n864), .C1(new_n865), .C2(G120gat), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(G1341gat));
  NOR2_X1   g669(.A1(new_n817), .A2(G127gat), .ZN(new_n871));
  INV_X1    g670(.A(new_n857), .ZN(new_n872));
  INV_X1    g671(.A(new_n851), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n453), .B(new_n871), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(G127gat), .B1(new_n847), .B2(new_n817), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n874), .A2(new_n875), .A3(KEYINPUT119), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1342gat));
  NOR3_X1   g679(.A1(new_n667), .A2(G134gat), .A3(new_n412), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n881), .B1(new_n873), .B2(new_n872), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n882), .A2(KEYINPUT56), .ZN(new_n883));
  OAI21_X1  g682(.A(G134gat), .B1(new_n847), .B2(new_n667), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(KEYINPUT56), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(G1343gat));
  NOR2_X1   g685(.A1(new_n683), .A2(new_n383), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n853), .A2(new_n450), .A3(new_n854), .A4(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n576), .A2(G141gat), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n888), .A2(new_n412), .A3(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT58), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT122), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n830), .A2(new_n834), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT120), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n830), .A2(new_n897), .A3(new_n834), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n896), .A2(new_n667), .A3(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n837), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n646), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n384), .B1(new_n901), .B2(new_n840), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT57), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n853), .A2(new_n904), .A3(new_n384), .A4(new_n854), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n722), .A2(new_n845), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n903), .A2(new_n575), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n891), .B1(new_n907), .B2(G141gat), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n850), .A2(new_n453), .A3(new_n887), .A4(new_n889), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT121), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT58), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n894), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n908), .B1(new_n894), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(G1344gat));
  NOR2_X1   g714(.A1(new_n888), .A2(new_n412), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n334), .A3(new_n632), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n918), .A2(new_n633), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n919), .A2(KEYINPUT59), .A3(new_n334), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n842), .A2(new_n843), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n384), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(KEYINPUT57), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n836), .A2(new_n667), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n899), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n841), .B1(new_n926), .B2(new_n646), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n904), .A3(new_n384), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n924), .A2(new_n928), .A3(new_n632), .A4(new_n906), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n921), .B1(new_n929), .B2(G148gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n917), .B1(new_n920), .B2(new_n930), .ZN(G1345gat));
  OAI21_X1  g730(.A(G155gat), .B1(new_n918), .B2(new_n817), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n916), .A2(new_n338), .A3(new_n646), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1346gat));
  OAI21_X1  g733(.A(G162gat), .B1(new_n918), .B2(new_n773), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n690), .A2(new_n339), .A3(new_n453), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n888), .B2(new_n936), .ZN(G1347gat));
  NOR2_X1   g736(.A1(new_n450), .A2(new_n453), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n844), .A2(new_n308), .A3(new_n938), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n939), .A2(new_n232), .A3(new_n576), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n922), .A2(new_n463), .A3(new_n938), .ZN(new_n941));
  AOI21_X1  g740(.A(G169gat), .B1(new_n941), .B2(new_n575), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n940), .A2(new_n942), .ZN(G1348gat));
  OAI21_X1  g742(.A(G176gat), .B1(new_n939), .B2(new_n633), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n941), .A2(new_n233), .A3(new_n632), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1349gat));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n947), .A2(KEYINPUT60), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n941), .A2(new_n255), .A3(new_n257), .A4(new_n646), .ZN(new_n949));
  OAI21_X1  g748(.A(G183gat), .B1(new_n939), .B2(new_n817), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n947), .A2(KEYINPUT60), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n951), .B(new_n952), .ZN(G1350gat));
  OAI21_X1  g752(.A(G190gat), .B1(new_n939), .B2(new_n667), .ZN(new_n954));
  NOR2_X1   g753(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n941), .A2(new_n220), .A3(new_n708), .ZN(new_n957));
  XNOR2_X1  g756(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n958));
  OAI211_X1 g757(.A(new_n956), .B(new_n957), .C1(new_n954), .C2(new_n958), .ZN(G1351gat));
  NAND2_X1  g758(.A1(new_n751), .A2(new_n938), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n924), .A2(new_n928), .A3(new_n575), .A4(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n567), .B1(new_n962), .B2(KEYINPUT125), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n963), .B1(KEYINPUT125), .B2(new_n962), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n923), .A2(new_n960), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n965), .A2(new_n567), .A3(new_n575), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(G1352gat));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n968));
  INV_X1    g767(.A(new_n965), .ZN(new_n969));
  AOI211_X1 g768(.A(G204gat), .B(new_n633), .C1(new_n968), .C2(KEYINPUT62), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  OR4_X1    g770(.A1(new_n968), .A2(new_n969), .A3(KEYINPUT62), .A4(new_n971), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n924), .A2(new_n928), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n973), .A2(new_n632), .A3(new_n961), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(G204gat), .ZN(new_n975));
  OAI22_X1  g774(.A1(new_n969), .A2(new_n971), .B1(new_n968), .B2(KEYINPUT62), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n972), .A2(new_n975), .A3(new_n976), .ZN(G1353gat));
  NAND3_X1  g776(.A1(new_n965), .A2(new_n321), .A3(new_n646), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n924), .A2(new_n928), .A3(new_n646), .A4(new_n961), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n979), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n980));
  AOI21_X1  g779(.A(KEYINPUT63), .B1(new_n979), .B2(G211gat), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(G1354gat));
  AOI21_X1  g781(.A(G218gat), .B1(new_n965), .B2(new_n708), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT127), .ZN(new_n984));
  OR2_X1    g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n983), .A2(new_n984), .ZN(new_n986));
  AND2_X1   g785(.A1(new_n973), .A2(new_n961), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n667), .A2(new_n354), .ZN(new_n988));
  AOI22_X1  g787(.A1(new_n985), .A2(new_n986), .B1(new_n987), .B2(new_n988), .ZN(G1355gat));
endmodule


