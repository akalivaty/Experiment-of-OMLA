//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n616, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160,
    new_n1161;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n454), .A2(new_n458), .B1(new_n449), .B2(new_n455), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT68), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  XOR2_X1   g036(.A(KEYINPUT3), .B(G2104), .Z(new_n462));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT69), .B(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n464), .A2(G2105), .B1(G101), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT71), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT71), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT3), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n469), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n476), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n469), .A2(KEYINPUT69), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2104), .ZN(new_n480));
  AND4_X1   g055(.A1(new_n476), .A2(new_n478), .A3(new_n480), .A4(KEYINPUT3), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n468), .B(new_n475), .C1(new_n477), .C2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G137), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n467), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  INV_X1    g060(.A(new_n482), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  OAI211_X1 g062(.A(G2105), .B(new_n475), .C1(new_n477), .C2(new_n481), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  AND2_X1   g065(.A1(G112), .A2(G2105), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(G100), .B2(new_n468), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n487), .B(new_n490), .C1(new_n469), .C2(new_n492), .ZN(new_n493));
  XOR2_X1   g068(.A(new_n493), .B(KEYINPUT72), .Z(G162));
  NAND3_X1  g069(.A1(new_n478), .A2(new_n480), .A3(KEYINPUT3), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT70), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n465), .A2(new_n476), .A3(KEYINPUT3), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n498), .A2(G138), .A3(new_n468), .A4(new_n475), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR4_X1   g076(.A1(new_n462), .A2(KEYINPUT4), .A3(new_n501), .A4(G2105), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  MUX2_X1   g079(.A(G102), .B(G114), .S(G2105), .Z(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G2104), .ZN(new_n506));
  INV_X1    g081(.A(G126), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n488), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g085(.A(KEYINPUT73), .B(new_n506), .C1(new_n488), .C2(new_n507), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n504), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n515), .B2(KEYINPUT75), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT75), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n517), .A2(KEYINPUT5), .A3(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT74), .B(G651), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  OAI211_X1 g098(.A(G88), .B(new_n519), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  OAI211_X1 g099(.A(G50), .B(G543), .C1(new_n522), .C2(new_n523), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n519), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n524), .B(new_n525), .C1(new_n520), .C2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT76), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n526), .A2(new_n520), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n530), .A2(KEYINPUT76), .A3(new_n524), .A4(new_n525), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(G166));
  NOR2_X1   g107(.A1(new_n522), .A2(new_n523), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n514), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  INV_X1    g110(.A(new_n519), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT77), .B(G89), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g114(.A1(G63), .A2(G651), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(KEYINPUT7), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(KEYINPUT7), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n519), .A2(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n535), .A2(new_n539), .A3(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  NAND2_X1  g121(.A1(new_n537), .A2(G90), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n534), .A2(G52), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n520), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  NAND2_X1  g127(.A1(new_n537), .A2(G81), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n534), .A2(G43), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(new_n520), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(new_n534), .A2(G53), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n536), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n537), .A2(G91), .B1(G651), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G166), .ZN(G303));
  NAND2_X1  g147(.A1(new_n537), .A2(G87), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n534), .A2(G49), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n536), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n520), .ZN(new_n580));
  AOI21_X1  g155(.A(KEYINPUT78), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  OAI211_X1 g157(.A(G86), .B(new_n519), .C1(new_n522), .C2(new_n523), .ZN(new_n583));
  OAI211_X1 g158(.A(G48), .B(G543), .C1(new_n522), .C2(new_n523), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n579), .A2(KEYINPUT78), .A3(new_n580), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n582), .A2(new_n585), .A3(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(new_n537), .A2(G85), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n534), .A2(G47), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n588), .B(new_n589), .C1(new_n520), .C2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT79), .Z(new_n593));
  NAND2_X1  g168(.A1(new_n537), .A2(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XOR2_X1   g171(.A(KEYINPUT80), .B(G66), .Z(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(new_n519), .B1(G79), .B2(G543), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(KEYINPUT81), .ZN(new_n599));
  INV_X1    g174(.A(G651), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(new_n598), .B2(KEYINPUT81), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n599), .A2(new_n601), .B1(new_n534), .B2(G54), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT82), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT83), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT82), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n603), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(KEYINPUT83), .ZN(new_n609));
  AND2_X1   g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n593), .B1(new_n610), .B2(G868), .ZN(G284));
  OAI21_X1  g186(.A(new_n593), .B1(new_n610), .B2(G868), .ZN(G321));
  NOR2_X1   g187(.A1(G299), .A2(G868), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g189(.A(new_n613), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n610), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND3_X1  g192(.A1(new_n606), .A2(new_n609), .A3(new_n616), .ZN(new_n618));
  MUX2_X1   g193(.A(new_n557), .B(new_n618), .S(G868), .Z(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g195(.A(new_n466), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n621), .A2(new_n462), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT13), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2100), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n486), .A2(G135), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n489), .A2(G123), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT84), .ZN(new_n628));
  OR3_X1    g203(.A1(new_n628), .A2(new_n468), .A3(G111), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n468), .B2(G111), .ZN(new_n630));
  OR2_X1    g205(.A1(G99), .A2(G2105), .ZN(new_n631));
  NAND4_X1  g206(.A1(new_n629), .A2(G2104), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  AND3_X1   g207(.A1(new_n626), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT85), .B(G2096), .Z(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n625), .A2(new_n636), .A3(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(KEYINPUT86), .B(KEYINPUT16), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n643), .B(new_n644), .Z(new_n645));
  XOR2_X1   g220(.A(KEYINPUT15), .B(G2435), .Z(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT87), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2430), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT14), .ZN(new_n652));
  INV_X1    g227(.A(new_n650), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n652), .B1(new_n648), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(G14), .B1(new_n645), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n654), .B2(new_n645), .ZN(G401));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  INV_X1    g238(.A(new_n659), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n660), .B1(new_n666), .B2(new_n657), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(new_n658), .B2(new_n665), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n658), .A2(new_n661), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n664), .B1(new_n669), .B2(KEYINPUT17), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n663), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(G2096), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2100), .ZN(G227));
  XNOR2_X1  g248(.A(G1956), .B(G2474), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1961), .B(G1966), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n674), .A2(new_n675), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n676), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  OR3_X1    g256(.A1(new_n681), .A2(KEYINPUT88), .A3(new_n678), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT20), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n681), .B1(KEYINPUT88), .B2(new_n678), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT89), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n689), .B(new_n692), .ZN(G229));
  MUX2_X1   g268(.A(G5), .B(G301), .S(G16), .Z(new_n694));
  NOR2_X1   g269(.A1(new_n694), .A2(G1961), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT90), .B(G16), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n697), .A2(G19), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n558), .B2(new_n697), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G1341), .ZN(new_n700));
  INV_X1    g275(.A(G2084), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  AND2_X1   g277(.A1(KEYINPUT24), .A2(G34), .ZN(new_n703));
  NOR2_X1   g278(.A1(KEYINPUT24), .A2(G34), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n484), .B2(new_n702), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT97), .Z(new_n707));
  AOI211_X1 g282(.A(new_n695), .B(new_n700), .C1(new_n701), .C2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(G27), .A2(G29), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G164), .B2(G29), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n708), .B1(G2078), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n702), .A2(G32), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n489), .A2(G129), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT98), .ZN(new_n714));
  NAND3_X1  g289(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT26), .Z(new_n716));
  INV_X1    g291(.A(G105), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n621), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n486), .B2(G141), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n712), .B1(new_n721), .B2(new_n702), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT27), .B(G1996), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n702), .A2(G26), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT28), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n486), .A2(G140), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n489), .A2(G128), .ZN(new_n728));
  AND2_X1   g303(.A1(G116), .A2(G2105), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G104), .B2(new_n468), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n727), .B(new_n728), .C1(new_n469), .C2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n726), .B1(new_n731), .B2(G29), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2067), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n724), .B(new_n733), .C1(new_n701), .C2(new_n707), .ZN(new_n734));
  NOR2_X1   g309(.A1(G29), .A2(G33), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n486), .A2(G139), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT94), .ZN(new_n737));
  NAND2_X1  g312(.A1(G115), .A2(G2104), .ZN(new_n738));
  INV_X1    g313(.A(G127), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n462), .B2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT25), .ZN(new_n741));
  NAND2_X1  g316(.A1(G103), .A2(G2104), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(G2105), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n468), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n740), .A2(G2105), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n737), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n735), .B1(new_n746), .B2(G29), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT95), .ZN(new_n748));
  INV_X1    g323(.A(G2072), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR3_X1   g325(.A1(new_n711), .A2(new_n734), .A3(new_n750), .ZN(new_n751));
  MUX2_X1   g326(.A(G21), .B(G286), .S(G16), .Z(new_n752));
  INV_X1    g327(.A(G1966), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n633), .A2(G29), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT99), .ZN(new_n756));
  OR2_X1    g331(.A1(KEYINPUT30), .A2(G28), .ZN(new_n757));
  NAND2_X1  g332(.A1(KEYINPUT30), .A2(G28), .ZN(new_n758));
  AOI21_X1  g333(.A(G29), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT31), .B(G11), .Z(new_n760));
  AOI211_X1 g335(.A(new_n759), .B(new_n760), .C1(new_n694), .C2(G1961), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n754), .A2(new_n756), .A3(new_n761), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT100), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n702), .A2(G35), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G162), .B2(new_n702), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT29), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n766), .A2(G2090), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n710), .A2(G2078), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n763), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G4), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n770), .A2(G16), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n606), .A2(new_n609), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1348), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n748), .A2(new_n749), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT96), .ZN(new_n776));
  AND4_X1   g351(.A1(new_n751), .A2(new_n769), .A3(new_n774), .A4(new_n776), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n585), .A2(new_n582), .A3(G16), .A4(new_n586), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G6), .B2(G16), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT91), .Z(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT32), .B(G1981), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT34), .ZN(new_n783));
  MUX2_X1   g358(.A(G23), .B(G288), .S(G16), .Z(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT33), .B(G1976), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n784), .B(new_n785), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n696), .A2(G22), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G166), .B2(new_n696), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1971), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n782), .A2(new_n783), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G25), .A2(G29), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n486), .A2(G131), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n489), .A2(G119), .ZN(new_n794));
  MUX2_X1   g369(.A(G95), .B(G107), .S(G2105), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(G2104), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n792), .B1(new_n798), .B2(G29), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT35), .B(G1991), .Z(new_n800));
  XOR2_X1   g375(.A(new_n799), .B(new_n800), .Z(new_n801));
  MUX2_X1   g376(.A(G24), .B(G290), .S(new_n697), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1986), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n791), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n783), .B1(new_n782), .B2(new_n790), .ZN(new_n806));
  OR3_X1    g381(.A1(new_n805), .A2(KEYINPUT93), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(KEYINPUT93), .B1(new_n805), .B2(new_n806), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT92), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(KEYINPUT36), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n777), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n807), .A2(new_n808), .B1(new_n810), .B2(KEYINPUT36), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n766), .A2(G2090), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT101), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n766), .A2(KEYINPUT101), .A3(G2090), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n696), .A2(G20), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT23), .Z(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G299), .B2(G16), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G1956), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n816), .A2(new_n817), .A3(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT102), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n812), .A2(new_n813), .A3(new_n823), .ZN(G311));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n813), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n809), .A2(new_n811), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n825), .A2(new_n826), .A3(new_n777), .ZN(G150));
  NAND2_X1  g402(.A1(new_n610), .A2(G559), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n537), .A2(G93), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n534), .A2(G55), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n829), .B(new_n830), .C1(new_n520), .C2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n557), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n828), .B(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n828), .B(new_n833), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(new_n836), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(G860), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n838), .A2(new_n840), .A3(KEYINPUT39), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n832), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT104), .B(KEYINPUT37), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n846), .A2(new_n849), .ZN(G145));
  INV_X1    g425(.A(new_n508), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n504), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n746), .B(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n720), .B(new_n731), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n797), .B(new_n623), .ZN(new_n856));
  MUX2_X1   g431(.A(G106), .B(G118), .S(G2105), .Z(new_n857));
  AOI22_X1  g432(.A1(new_n489), .A2(G130), .B1(G2104), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(G142), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n858), .B1(new_n859), .B2(new_n482), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n856), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(G162), .B(G160), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n633), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n855), .A2(new_n861), .ZN(new_n866));
  AOI21_X1  g441(.A(G37), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n862), .A2(KEYINPUT105), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(new_n866), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n862), .A2(KEYINPUT105), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n867), .B1(new_n871), .B2(new_n864), .ZN(new_n872));
  XOR2_X1   g447(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(G395));
  NOR2_X1   g449(.A1(new_n832), .A2(G868), .ZN(new_n875));
  XOR2_X1   g450(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n876));
  NAND3_X1  g451(.A1(new_n610), .A2(new_n616), .A3(new_n833), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n618), .A2(new_n834), .ZN(new_n878));
  XNOR2_X1  g453(.A(G299), .B(new_n603), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(G288), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(G290), .ZN(new_n884));
  XNOR2_X1  g459(.A(G166), .B(G305), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n886), .B(KEYINPUT107), .Z(new_n887));
  NOR2_X1   g462(.A1(new_n884), .A2(new_n885), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n879), .B(KEYINPUT41), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n891), .B1(new_n877), .B2(new_n878), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n882), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n889), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n877), .A2(new_n878), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n890), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n894), .B1(new_n896), .B2(new_n881), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n876), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n889), .B1(new_n882), .B2(new_n892), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n896), .A2(new_n894), .A3(new_n881), .ZN(new_n900));
  INV_X1    g475(.A(new_n876), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n875), .B1(new_n903), .B2(G868), .ZN(G295));
  AOI21_X1  g479(.A(new_n875), .B1(new_n903), .B2(G868), .ZN(G331));
  XNOR2_X1  g480(.A(G286), .B(G301), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n833), .B(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n907), .A2(new_n879), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n908), .B1(new_n890), .B2(new_n907), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n894), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(G37), .B1(new_n894), .B2(new_n909), .ZN(new_n912));
  XNOR2_X1  g487(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT110), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT110), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n911), .A2(new_n912), .A3(new_n916), .A4(new_n913), .ZN(new_n917));
  INV_X1    g492(.A(new_n912), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT43), .B1(new_n918), .B2(new_n910), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n915), .A2(KEYINPUT44), .A3(new_n917), .A4(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n913), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(new_n918), .B2(new_n910), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n922), .A2(new_n914), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n920), .B1(KEYINPUT44), .B2(new_n923), .ZN(G397));
  INV_X1    g499(.A(G1996), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n721), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(G2067), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n731), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n720), .A2(G1996), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n798), .A2(new_n800), .ZN(new_n932));
  OAI22_X1  g507(.A1(new_n931), .A2(new_n932), .B1(G2067), .B2(new_n731), .ZN(new_n933));
  INV_X1    g508(.A(G1384), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n502), .B1(new_n499), .B2(KEYINPUT4), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n934), .B1(new_n935), .B2(new_n508), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g513(.A(KEYINPUT111), .B(new_n934), .C1(new_n935), .C2(new_n508), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT45), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n467), .B(G40), .C1(new_n483), .C2(new_n482), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n933), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n928), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n944), .B1(new_n720), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT46), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n948), .B1(new_n944), .B2(new_n925), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n943), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n951), .B(KEYINPUT47), .Z(new_n952));
  OR2_X1    g527(.A1(new_n798), .A2(new_n800), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n930), .A2(new_n932), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n944), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT127), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n943), .A2(G1986), .A3(G290), .ZN(new_n957));
  XOR2_X1   g532(.A(new_n957), .B(KEYINPUT48), .Z(new_n958));
  AOI211_X1 g533(.A(new_n945), .B(new_n952), .C1(new_n956), .C2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT51), .ZN(new_n960));
  AOI211_X1 g535(.A(KEYINPUT123), .B(new_n960), .C1(G286), .C2(G8), .ZN(new_n961));
  NAND2_X1  g536(.A1(G286), .A2(G8), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n961), .B1(new_n963), .B2(KEYINPUT123), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n512), .A2(KEYINPUT50), .A3(new_n934), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n936), .A2(new_n967), .ZN(new_n968));
  AOI211_X1 g543(.A(G2084), .B(new_n941), .C1(new_n966), .C2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n941), .B1(new_n936), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT116), .ZN(new_n972));
  AOI22_X1  g547(.A1(new_n500), .A2(new_n503), .B1(new_n508), .B2(new_n509), .ZN(new_n973));
  AOI21_X1  g548(.A(G1384), .B1(new_n973), .B2(new_n511), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n972), .B1(new_n974), .B2(KEYINPUT45), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n512), .A2(new_n972), .A3(KEYINPUT45), .A4(new_n934), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n971), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n969), .B1(new_n978), .B2(new_n753), .ZN(new_n979));
  INV_X1    g554(.A(G8), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n965), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n941), .B1(new_n966), .B2(new_n968), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n701), .ZN(new_n983));
  INV_X1    g558(.A(new_n971), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n512), .A2(KEYINPUT45), .A3(new_n934), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT116), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n984), .B1(new_n986), .B2(new_n976), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n983), .B1(new_n987), .B2(G1966), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n960), .B(G8), .C1(new_n988), .C2(G286), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(G8), .A3(G286), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n981), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n991), .A2(KEYINPUT62), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n529), .A2(G8), .A3(new_n531), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n529), .A2(KEYINPUT55), .A3(G8), .A4(new_n531), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G2090), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT50), .B1(new_n512), .B2(new_n934), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT50), .B(new_n934), .C1(new_n935), .C2(new_n508), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n999), .B(new_n942), .C1(new_n1000), .C2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n1004));
  INV_X1    g579(.A(G1971), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT45), .B1(new_n512), .B2(new_n934), .ZN(new_n1006));
  OAI211_X1 g581(.A(KEYINPUT45), .B(new_n934), .C1(new_n935), .C2(new_n508), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n942), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1005), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1003), .A2(new_n1004), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(G8), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1004), .B1(new_n1003), .B2(new_n1009), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n998), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n982), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT124), .B(G1961), .Z(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n512), .A2(new_n934), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n970), .ZN(new_n1018));
  INV_X1    g593(.A(G2078), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1008), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1014), .A2(new_n1016), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(G2078), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n987), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(G301), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(G1384), .B1(new_n504), .B2(new_n851), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n942), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n883), .A2(G1976), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(G8), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT52), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT49), .ZN(new_n1032));
  NOR2_X1   g607(.A1(G305), .A2(G1981), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n579), .A2(new_n580), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n585), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(G1981), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1032), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1036), .B(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1038), .A2(G8), .A3(new_n1028), .A4(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G1976), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT52), .B1(G288), .B2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1028), .A2(G8), .A3(new_n1029), .A4(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1031), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n982), .A2(new_n999), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n980), .B1(new_n1045), .B2(new_n1009), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n997), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n995), .A2(KEYINPUT113), .A3(new_n996), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1044), .B1(new_n1046), .B2(new_n1050), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n1013), .A2(new_n1026), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT62), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n981), .A2(new_n989), .A3(new_n1053), .A4(new_n990), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT126), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1052), .A2(new_n1054), .A3(KEYINPUT126), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n992), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n938), .A2(new_n939), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n970), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1007), .A2(new_n942), .A3(new_n1024), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1062), .A2(KEYINPUT125), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT125), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1066), .B1(new_n940), .B2(new_n1063), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1006), .A2(G2078), .A3(new_n1008), .ZN(new_n1069));
  OAI22_X1  g644(.A1(new_n1069), .A2(KEYINPUT53), .B1(new_n982), .B2(new_n1015), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1068), .A2(G171), .A3(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1060), .B1(new_n1071), .B2(new_n1026), .ZN(new_n1072));
  AOI211_X1 g647(.A(G2090), .B(new_n941), .C1(new_n966), .C2(new_n968), .ZN(new_n1073));
  AOI21_X1  g648(.A(G1971), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1074));
  OAI211_X1 g649(.A(G8), .B(new_n1050), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1031), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1012), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1078), .A2(G8), .A3(new_n1010), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1077), .B1(new_n1079), .B2(new_n998), .ZN(new_n1080));
  OAI21_X1  g655(.A(G171), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1023), .A2(G301), .A3(new_n1025), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(KEYINPUT54), .A3(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1072), .A2(new_n991), .A3(new_n1080), .A4(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n1085));
  NAND3_X1  g660(.A1(G299), .A2(new_n1085), .A3(KEYINPUT57), .ZN(new_n1086));
  OR2_X1    g661(.A1(new_n1085), .A2(KEYINPUT57), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(KEYINPUT57), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n566), .A2(new_n570), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1001), .B1(new_n974), .B2(KEYINPUT50), .ZN(new_n1091));
  AOI21_X1  g666(.A(G1956), .B1(new_n1091), .B2(new_n942), .ZN(new_n1092));
  XOR2_X1   g667(.A(KEYINPUT56), .B(G2072), .Z(new_n1093));
  NOR3_X1   g668(.A1(new_n1006), .A2(new_n1008), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1090), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT118), .ZN(new_n1096));
  NOR4_X1   g671(.A1(new_n1092), .A2(new_n1090), .A3(new_n1094), .A4(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n942), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1098));
  INV_X1    g673(.A(G1956), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1008), .B1(new_n970), .B2(new_n1017), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1093), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1098), .A2(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1090), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT118), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1095), .B1(new_n1097), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT61), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT61), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1092), .A2(new_n1090), .A3(new_n1094), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1108), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1112), .A2(new_n1095), .A3(KEYINPUT121), .A4(KEYINPUT61), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n982), .A2(G1348), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT119), .B1(new_n1027), .B2(new_n942), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n936), .A2(new_n1117), .A3(new_n941), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n927), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT60), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1119), .B(KEYINPUT60), .C1(new_n982), .C2(G1348), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(new_n1124), .A3(new_n604), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1115), .A2(KEYINPUT60), .A3(new_n608), .A4(new_n1119), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1124), .B1(new_n1123), .B2(new_n604), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1122), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT58), .B(G1341), .ZN(new_n1130));
  OR3_X1    g705(.A1(new_n1116), .A2(new_n1118), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1100), .A2(new_n925), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n557), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n1133), .B(KEYINPUT59), .Z(new_n1134));
  NAND4_X1  g709(.A1(new_n1107), .A2(new_n1114), .A3(new_n1129), .A4(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1120), .A2(KEYINPUT120), .A3(new_n604), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n1095), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT120), .B1(new_n1120), .B2(new_n604), .ZN(new_n1138));
  OAI22_X1  g713(.A1(new_n1137), .A2(new_n1138), .B1(new_n1104), .B2(new_n1097), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1084), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1028), .A2(G8), .ZN(new_n1141));
  XOR2_X1   g716(.A(new_n1141), .B(KEYINPUT114), .Z(new_n1142));
  INV_X1    g717(.A(new_n1033), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1040), .A2(new_n1041), .A3(new_n883), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1075), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1145), .B1(new_n1146), .B2(new_n1076), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n979), .A2(new_n980), .A3(G286), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT63), .B1(new_n1080), .B2(new_n1148), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n1046), .A2(new_n997), .ZN(new_n1150));
  AND4_X1   g725(.A1(KEYINPUT63), .A2(new_n1148), .A3(new_n1051), .A4(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1147), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1059), .A2(new_n1140), .A3(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(G290), .B(G1986), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n944), .B1(new_n954), .B2(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT112), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n959), .B1(new_n1153), .B2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g732(.A1(new_n922), .A2(new_n914), .ZN(new_n1159));
  INV_X1    g733(.A(G319), .ZN(new_n1160));
  NOR4_X1   g734(.A1(G229), .A2(G227), .A3(new_n1160), .A4(G401), .ZN(new_n1161));
  NAND3_X1  g735(.A1(new_n1159), .A2(new_n872), .A3(new_n1161), .ZN(G225));
  INV_X1    g736(.A(G225), .ZN(G308));
endmodule


