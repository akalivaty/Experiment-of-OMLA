

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588;

  NOR2_X1 U322 ( .A1(n418), .A2(n524), .ZN(n420) );
  XNOR2_X1 U323 ( .A(n300), .B(n299), .ZN(n304) );
  NOR2_X1 U324 ( .A1(n456), .A2(n473), .ZN(n457) );
  XOR2_X1 U325 ( .A(n327), .B(n326), .Z(n561) );
  XOR2_X1 U326 ( .A(KEYINPUT38), .B(n481), .Z(n509) );
  XNOR2_X1 U327 ( .A(n393), .B(n433), .ZN(n526) );
  XOR2_X1 U328 ( .A(n297), .B(n296), .Z(n290) );
  XOR2_X1 U329 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n291) );
  XOR2_X1 U330 ( .A(KEYINPUT37), .B(KEYINPUT102), .Z(n292) );
  NOR2_X1 U331 ( .A1(n570), .A2(n471), .ZN(n293) );
  INV_X1 U332 ( .A(KEYINPUT110), .ZN(n365) );
  XOR2_X1 U333 ( .A(KEYINPUT13), .B(G57GAT), .Z(n317) );
  INV_X1 U334 ( .A(n317), .ZN(n318) );
  NOR2_X1 U335 ( .A1(n524), .A2(n469), .ZN(n470) );
  XNOR2_X1 U336 ( .A(n298), .B(n290), .ZN(n299) );
  INV_X1 U337 ( .A(KEYINPUT64), .ZN(n419) );
  XOR2_X1 U338 ( .A(n368), .B(KEYINPUT36), .Z(n584) );
  XNOR2_X1 U339 ( .A(n309), .B(n308), .ZN(n577) );
  XNOR2_X1 U340 ( .A(n480), .B(n292), .ZN(n522) );
  XOR2_X1 U341 ( .A(KEYINPUT119), .B(n457), .Z(n566) );
  XOR2_X1 U342 ( .A(n455), .B(n454), .Z(n537) );
  XNOR2_X1 U343 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U344 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n482) );
  XNOR2_X1 U345 ( .A(n489), .B(n488), .ZN(G1351GAT) );
  XNOR2_X1 U346 ( .A(n483), .B(n482), .ZN(G1330GAT) );
  XNOR2_X1 U347 ( .A(KEYINPUT55), .B(KEYINPUT118), .ZN(n437) );
  XOR2_X1 U348 ( .A(KEYINPUT31), .B(n317), .Z(n295) );
  XOR2_X1 U349 ( .A(G176GAT), .B(G64GAT), .Z(n375) );
  XNOR2_X1 U350 ( .A(G204GAT), .B(n375), .ZN(n294) );
  XNOR2_X1 U351 ( .A(n295), .B(n294), .ZN(n300) );
  XOR2_X1 U352 ( .A(G120GAT), .B(G71GAT), .Z(n445) );
  XNOR2_X1 U353 ( .A(n445), .B(KEYINPUT76), .ZN(n298) );
  XOR2_X1 U354 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n297) );
  NAND2_X1 U355 ( .A1(G230GAT), .A2(G233GAT), .ZN(n296) );
  XOR2_X1 U356 ( .A(KEYINPUT32), .B(KEYINPUT72), .Z(n302) );
  XNOR2_X1 U357 ( .A(KEYINPUT71), .B(KEYINPUT75), .ZN(n301) );
  XOR2_X1 U358 ( .A(n302), .B(n301), .Z(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n309) );
  XNOR2_X1 U360 ( .A(G106GAT), .B(G78GAT), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n305), .B(G148GAT), .ZN(n427) );
  XOR2_X1 U362 ( .A(G85GAT), .B(KEYINPUT74), .Z(n307) );
  XNOR2_X1 U363 ( .A(G99GAT), .B(G92GAT), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n335) );
  XNOR2_X1 U365 ( .A(n427), .B(n335), .ZN(n308) );
  XOR2_X1 U366 ( .A(G64GAT), .B(G71GAT), .Z(n311) );
  XNOR2_X1 U367 ( .A(G8GAT), .B(G183GAT), .ZN(n310) );
  XNOR2_X1 U368 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U369 ( .A(KEYINPUT12), .B(KEYINPUT80), .Z(n313) );
  XNOR2_X1 U370 ( .A(G1GAT), .B(KEYINPUT15), .ZN(n312) );
  XNOR2_X1 U371 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n315), .B(n314), .ZN(n327) );
  XOR2_X1 U373 ( .A(G22GAT), .B(G155GAT), .Z(n424) );
  XNOR2_X1 U374 ( .A(G211GAT), .B(G78GAT), .ZN(n316) );
  XNOR2_X1 U375 ( .A(n424), .B(n316), .ZN(n319) );
  XNOR2_X1 U376 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U377 ( .A(KEYINPUT14), .B(KEYINPUT82), .Z(n321) );
  NAND2_X1 U378 ( .A1(G231GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U380 ( .A(n323), .B(n322), .Z(n325) );
  XOR2_X1 U381 ( .A(G15GAT), .B(G127GAT), .Z(n441) );
  XNOR2_X1 U382 ( .A(n441), .B(KEYINPUT81), .ZN(n324) );
  XNOR2_X1 U383 ( .A(n325), .B(n324), .ZN(n326) );
  INV_X1 U384 ( .A(n561), .ZN(n581) );
  XOR2_X1 U385 ( .A(G50GAT), .B(G162GAT), .Z(n428) );
  XOR2_X1 U386 ( .A(KEYINPUT9), .B(G106GAT), .Z(n329) );
  XNOR2_X1 U387 ( .A(G134GAT), .B(G218GAT), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U389 ( .A(n428), .B(n330), .Z(n332) );
  NAND2_X1 U390 ( .A1(G232GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U391 ( .A(n332), .B(n331), .ZN(n343) );
  XOR2_X1 U392 ( .A(KEYINPUT77), .B(KEYINPUT79), .Z(n334) );
  XNOR2_X1 U393 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n333) );
  XNOR2_X1 U394 ( .A(n334), .B(n333), .ZN(n336) );
  XOR2_X1 U395 ( .A(n336), .B(n335), .Z(n341) );
  XNOR2_X1 U396 ( .A(G43GAT), .B(G29GAT), .ZN(n337) );
  XNOR2_X1 U397 ( .A(n291), .B(n337), .ZN(n338) );
  XOR2_X1 U398 ( .A(KEYINPUT69), .B(n338), .Z(n358) );
  XNOR2_X1 U399 ( .A(G36GAT), .B(G190GAT), .ZN(n339) );
  XNOR2_X1 U400 ( .A(n339), .B(KEYINPUT78), .ZN(n376) );
  XNOR2_X1 U401 ( .A(n358), .B(n376), .ZN(n340) );
  XNOR2_X1 U402 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n343), .B(n342), .ZN(n368) );
  NAND2_X1 U404 ( .A1(n581), .A2(n584), .ZN(n346) );
  XOR2_X1 U405 ( .A(KEYINPUT109), .B(KEYINPUT45), .Z(n344) );
  XNOR2_X1 U406 ( .A(KEYINPUT65), .B(n344), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n346), .B(n345), .ZN(n363) );
  XOR2_X1 U408 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n348) );
  XNOR2_X1 U409 ( .A(KEYINPUT66), .B(KEYINPUT67), .ZN(n347) );
  XNOR2_X1 U410 ( .A(n348), .B(n347), .ZN(n362) );
  XOR2_X1 U411 ( .A(G15GAT), .B(G22GAT), .Z(n350) );
  XNOR2_X1 U412 ( .A(G141GAT), .B(G197GAT), .ZN(n349) );
  XNOR2_X1 U413 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U414 ( .A(n351), .B(G36GAT), .Z(n353) );
  XOR2_X1 U415 ( .A(G113GAT), .B(G1GAT), .Z(n399) );
  XNOR2_X1 U416 ( .A(n399), .B(G50GAT), .ZN(n352) );
  XNOR2_X1 U417 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U418 ( .A(KEYINPUT70), .B(KEYINPUT29), .Z(n355) );
  NAND2_X1 U419 ( .A1(G229GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U420 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U421 ( .A(n357), .B(n356), .Z(n360) );
  XOR2_X1 U422 ( .A(G169GAT), .B(G8GAT), .Z(n383) );
  XNOR2_X1 U423 ( .A(n358), .B(n383), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n362), .B(n361), .ZN(n571) );
  INV_X1 U426 ( .A(n571), .ZN(n553) );
  NAND2_X1 U427 ( .A1(n363), .A2(n553), .ZN(n364) );
  NOR2_X1 U428 ( .A1(n577), .A2(n364), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n366), .B(n365), .ZN(n373) );
  XOR2_X1 U430 ( .A(KEYINPUT41), .B(n577), .Z(n555) );
  AND2_X1 U431 ( .A1(n555), .A2(n571), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n367), .B(KEYINPUT46), .ZN(n370) );
  NAND2_X1 U433 ( .A1(n368), .A2(n561), .ZN(n369) );
  NOR2_X1 U434 ( .A1(n370), .A2(n369), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n371), .B(KEYINPUT47), .ZN(n372) );
  NAND2_X1 U436 ( .A1(n373), .A2(n372), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n374), .B(KEYINPUT48), .ZN(n533) );
  XNOR2_X1 U438 ( .A(n376), .B(n375), .ZN(n378) );
  AND2_X1 U439 ( .A1(G226GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U440 ( .A(n378), .B(n377), .ZN(n380) );
  INV_X1 U441 ( .A(KEYINPUT95), .ZN(n379) );
  NAND2_X1 U442 ( .A1(n380), .A2(n379), .ZN(n382) );
  OR2_X1 U443 ( .A1(n380), .A2(n379), .ZN(n381) );
  NAND2_X1 U444 ( .A1(n382), .A2(n381), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n383), .B(G92GAT), .ZN(n384) );
  XNOR2_X1 U446 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U447 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n387) );
  XNOR2_X1 U448 ( .A(KEYINPUT86), .B(G183GAT), .ZN(n386) );
  XNOR2_X1 U449 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U450 ( .A(KEYINPUT19), .B(n388), .Z(n453) );
  XNOR2_X1 U451 ( .A(n389), .B(n453), .ZN(n393) );
  XOR2_X1 U452 ( .A(G211GAT), .B(G218GAT), .Z(n391) );
  XNOR2_X1 U453 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n390) );
  XNOR2_X1 U454 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U455 ( .A(G197GAT), .B(n392), .ZN(n433) );
  NAND2_X1 U456 ( .A1(n533), .A2(n526), .ZN(n395) );
  XOR2_X1 U457 ( .A(KEYINPUT117), .B(KEYINPUT54), .Z(n394) );
  XNOR2_X1 U458 ( .A(n395), .B(n394), .ZN(n418) );
  XOR2_X1 U459 ( .A(G85GAT), .B(G148GAT), .Z(n397) );
  XNOR2_X1 U460 ( .A(G29GAT), .B(G162GAT), .ZN(n396) );
  XNOR2_X1 U461 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U462 ( .A(n399), .B(n398), .Z(n401) );
  NAND2_X1 U463 ( .A1(G225GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U464 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U465 ( .A(n402), .B(KEYINPUT5), .Z(n405) );
  XNOR2_X1 U466 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n403) );
  XNOR2_X1 U467 ( .A(n403), .B(KEYINPUT83), .ZN(n444) );
  XNOR2_X1 U468 ( .A(n444), .B(KEYINPUT93), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U470 ( .A(G57GAT), .B(G155GAT), .Z(n407) );
  XNOR2_X1 U471 ( .A(G120GAT), .B(G127GAT), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U473 ( .A(n409), .B(n408), .Z(n417) );
  XOR2_X1 U474 ( .A(KEYINPUT2), .B(KEYINPUT90), .Z(n411) );
  XNOR2_X1 U475 ( .A(KEYINPUT91), .B(KEYINPUT3), .ZN(n410) );
  XNOR2_X1 U476 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U477 ( .A(G141GAT), .B(n412), .Z(n434) );
  XOR2_X1 U478 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n414) );
  XNOR2_X1 U479 ( .A(KEYINPUT1), .B(KEYINPUT94), .ZN(n413) );
  XNOR2_X1 U480 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U481 ( .A(n434), .B(n415), .ZN(n416) );
  XNOR2_X1 U482 ( .A(n417), .B(n416), .ZN(n524) );
  XNOR2_X1 U483 ( .A(n420), .B(n419), .ZN(n570) );
  XOR2_X1 U484 ( .A(KEYINPUT92), .B(KEYINPUT22), .Z(n422) );
  XNOR2_X1 U485 ( .A(KEYINPUT23), .B(KEYINPUT88), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U487 ( .A(n423), .B(KEYINPUT24), .Z(n426) );
  XNOR2_X1 U488 ( .A(n424), .B(KEYINPUT89), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n432) );
  XOR2_X1 U490 ( .A(n428), .B(n427), .Z(n430) );
  NAND2_X1 U491 ( .A1(G228GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U492 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U493 ( .A(n432), .B(n431), .Z(n436) );
  XOR2_X1 U494 ( .A(n434), .B(n433), .Z(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n471) );
  XNOR2_X1 U496 ( .A(n437), .B(n293), .ZN(n456) );
  XOR2_X1 U497 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n439) );
  XNOR2_X1 U498 ( .A(G113GAT), .B(G99GAT), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U500 ( .A(n440), .B(G190GAT), .Z(n443) );
  XNOR2_X1 U501 ( .A(G43GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U502 ( .A(n443), .B(n442), .ZN(n449) );
  XOR2_X1 U503 ( .A(n445), .B(n444), .Z(n447) );
  NAND2_X1 U504 ( .A1(G227GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U506 ( .A(n449), .B(n448), .Z(n455) );
  XOR2_X1 U507 ( .A(G176GAT), .B(KEYINPUT87), .Z(n451) );
  XNOR2_X1 U508 ( .A(G169GAT), .B(KEYINPUT85), .ZN(n450) );
  XNOR2_X1 U509 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U510 ( .A(n453), .B(n452), .ZN(n454) );
  INV_X1 U511 ( .A(n537), .ZN(n473) );
  NAND2_X1 U512 ( .A1(n566), .A2(n555), .ZN(n461) );
  XOR2_X1 U513 ( .A(G176GAT), .B(KEYINPUT56), .Z(n459) );
  XOR2_X1 U514 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n458) );
  XNOR2_X1 U515 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U516 ( .A(n461), .B(n460), .ZN(G1349GAT) );
  INV_X1 U517 ( .A(n526), .ZN(n462) );
  XOR2_X1 U518 ( .A(KEYINPUT27), .B(n462), .Z(n472) );
  NAND2_X1 U519 ( .A1(n471), .A2(n473), .ZN(n463) );
  XOR2_X1 U520 ( .A(n463), .B(KEYINPUT26), .Z(n568) );
  AND2_X1 U521 ( .A1(n472), .A2(n568), .ZN(n468) );
  AND2_X1 U522 ( .A1(n537), .A2(n526), .ZN(n464) );
  NOR2_X1 U523 ( .A1(n471), .A2(n464), .ZN(n465) );
  XOR2_X1 U524 ( .A(n465), .B(KEYINPUT96), .Z(n466) );
  XNOR2_X1 U525 ( .A(n466), .B(KEYINPUT25), .ZN(n467) );
  NOR2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U527 ( .A(n470), .B(KEYINPUT97), .ZN(n476) );
  XNOR2_X1 U528 ( .A(n471), .B(KEYINPUT28), .ZN(n539) );
  NAND2_X1 U529 ( .A1(n524), .A2(n472), .ZN(n534) );
  NOR2_X1 U530 ( .A1(n539), .A2(n534), .ZN(n474) );
  NAND2_X1 U531 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND2_X1 U532 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U533 ( .A(KEYINPUT98), .B(n477), .ZN(n497) );
  NAND2_X1 U534 ( .A1(n497), .A2(n561), .ZN(n478) );
  XNOR2_X1 U535 ( .A(n478), .B(KEYINPUT101), .ZN(n479) );
  NAND2_X1 U536 ( .A1(n479), .A2(n584), .ZN(n480) );
  OR2_X1 U537 ( .A1(n553), .A2(n577), .ZN(n499) );
  OR2_X1 U538 ( .A1(n522), .A2(n499), .ZN(n481) );
  NAND2_X1 U539 ( .A1(n509), .A2(n537), .ZN(n483) );
  NAND2_X1 U540 ( .A1(n509), .A2(n526), .ZN(n485) );
  XNOR2_X1 U541 ( .A(G36GAT), .B(KEYINPUT104), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n485), .B(n484), .ZN(G1329GAT) );
  INV_X1 U543 ( .A(n368), .ZN(n548) );
  NAND2_X1 U544 ( .A1(n566), .A2(n548), .ZN(n489) );
  XOR2_X1 U545 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n487) );
  INV_X1 U546 ( .A(G190GAT), .ZN(n486) );
  NAND2_X1 U547 ( .A1(n571), .A2(n566), .ZN(n491) );
  XNOR2_X1 U548 ( .A(KEYINPUT120), .B(G169GAT), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n491), .B(n490), .ZN(G1348GAT) );
  NAND2_X1 U550 ( .A1(n524), .A2(n509), .ZN(n495) );
  XOR2_X1 U551 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n493) );
  INV_X1 U552 ( .A(G29GAT), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n495), .B(n494), .ZN(G1328GAT) );
  NOR2_X1 U555 ( .A1(n548), .A2(n561), .ZN(n496) );
  XNOR2_X1 U556 ( .A(KEYINPUT16), .B(n496), .ZN(n498) );
  NAND2_X1 U557 ( .A1(n498), .A2(n497), .ZN(n512) );
  NOR2_X1 U558 ( .A1(n499), .A2(n512), .ZN(n506) );
  NAND2_X1 U559 ( .A1(n506), .A2(n524), .ZN(n500) );
  XNOR2_X1 U560 ( .A(n500), .B(KEYINPUT34), .ZN(n501) );
  XNOR2_X1 U561 ( .A(G1GAT), .B(n501), .ZN(G1324GAT) );
  NAND2_X1 U562 ( .A1(n526), .A2(n506), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n502), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n504) );
  NAND2_X1 U565 ( .A1(n506), .A2(n537), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U567 ( .A(G15GAT), .B(n505), .Z(G1326GAT) );
  NAND2_X1 U568 ( .A1(n539), .A2(n506), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n507), .B(KEYINPUT100), .ZN(n508) );
  XNOR2_X1 U570 ( .A(G22GAT), .B(n508), .ZN(G1327GAT) );
  NAND2_X1 U571 ( .A1(n509), .A2(n539), .ZN(n510) );
  XNOR2_X1 U572 ( .A(n510), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 U573 ( .A1(n555), .A2(n553), .ZN(n511) );
  XOR2_X1 U574 ( .A(n511), .B(KEYINPUT105), .Z(n523) );
  NOR2_X1 U575 ( .A1(n523), .A2(n512), .ZN(n519) );
  NAND2_X1 U576 ( .A1(n524), .A2(n519), .ZN(n513) );
  XNOR2_X1 U577 ( .A(KEYINPUT42), .B(n513), .ZN(n514) );
  XNOR2_X1 U578 ( .A(G57GAT), .B(n514), .ZN(G1332GAT) );
  NAND2_X1 U579 ( .A1(n526), .A2(n519), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n517) );
  NAND2_X1 U582 ( .A1(n519), .A2(n537), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U584 ( .A(G71GAT), .B(n518), .ZN(G1334GAT) );
  XOR2_X1 U585 ( .A(G78GAT), .B(KEYINPUT43), .Z(n521) );
  NAND2_X1 U586 ( .A1(n519), .A2(n539), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(G1335GAT) );
  NOR2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n530) );
  NAND2_X1 U589 ( .A1(n530), .A2(n524), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U591 ( .A1(n526), .A2(n530), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n527), .B(KEYINPUT108), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G92GAT), .B(n528), .ZN(G1337GAT) );
  NAND2_X1 U594 ( .A1(n537), .A2(n530), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n529), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U596 ( .A1(n539), .A2(n530), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n531), .B(KEYINPUT44), .ZN(n532) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  INV_X1 U599 ( .A(n534), .ZN(n535) );
  NAND2_X1 U600 ( .A1(n533), .A2(n535), .ZN(n536) );
  XNOR2_X1 U601 ( .A(KEYINPUT111), .B(n536), .ZN(n552) );
  NAND2_X1 U602 ( .A1(n552), .A2(n537), .ZN(n538) );
  NOR2_X1 U603 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U604 ( .A(KEYINPUT112), .B(n540), .ZN(n547) );
  NAND2_X1 U605 ( .A1(n547), .A2(n571), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n541), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n543) );
  NAND2_X1 U608 ( .A1(n555), .A2(n547), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U610 ( .A(G120GAT), .B(n544), .Z(G1341GAT) );
  NAND2_X1 U611 ( .A1(n547), .A2(n581), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n545), .B(KEYINPUT50), .ZN(n546) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U615 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G134GAT), .B(n551), .ZN(G1343GAT) );
  NAND2_X1 U618 ( .A1(n552), .A2(n568), .ZN(n564) );
  NOR2_X1 U619 ( .A1(n553), .A2(n564), .ZN(n554) );
  XOR2_X1 U620 ( .A(G141GAT), .B(n554), .Z(G1344GAT) );
  INV_X1 U621 ( .A(n555), .ZN(n556) );
  NOR2_X1 U622 ( .A1(n564), .A2(n556), .ZN(n560) );
  XOR2_X1 U623 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n558) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(KEYINPUT115), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1345GAT) );
  NOR2_X1 U627 ( .A1(n561), .A2(n564), .ZN(n562) );
  XOR2_X1 U628 ( .A(KEYINPUT116), .B(n562), .Z(n563) );
  XNOR2_X1 U629 ( .A(G155GAT), .B(n563), .ZN(G1346GAT) );
  NOR2_X1 U630 ( .A1(n368), .A2(n564), .ZN(n565) );
  XOR2_X1 U631 ( .A(G162GAT), .B(n565), .Z(G1347GAT) );
  NAND2_X1 U632 ( .A1(n566), .A2(n581), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n573) );
  INV_X1 U635 ( .A(n568), .ZN(n569) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n585) );
  NAND2_X1 U637 ( .A1(n585), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(n574), .B(KEYINPUT59), .Z(n576) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n579) );
  NAND2_X1 U643 ( .A1(n585), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XOR2_X1 U645 ( .A(G204GAT), .B(n580), .Z(G1353GAT) );
  NAND2_X1 U646 ( .A1(n585), .A2(n581), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(KEYINPUT126), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G211GAT), .B(n583), .ZN(G1354GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n587) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

