

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856;

  XNOR2_X1 U379 ( .A(n362), .B(KEYINPUT41), .ZN(n808) );
  INV_X1 U380 ( .A(n709), .ZN(n358) );
  NOR2_X1 U381 ( .A1(n505), .A2(n793), .ZN(n504) );
  AND2_X2 U382 ( .A1(n700), .A2(n701), .ZN(n426) );
  BUF_X2 U383 ( .A(n845), .Z(n460) );
  NOR2_X2 U384 ( .A1(n797), .A2(n657), .ZN(n658) );
  XNOR2_X2 U385 ( .A(KEYINPUT77), .B(KEYINPUT22), .ZN(n640) );
  AND2_X2 U386 ( .A1(n426), .A2(n702), .ZN(n703) );
  AND2_X2 U387 ( .A1(n410), .A2(n406), .ZN(n405) );
  NAND2_X2 U388 ( .A1(n405), .A2(n403), .ZN(n412) );
  NOR2_X1 U389 ( .A1(n471), .A2(KEYINPUT47), .ZN(n433) );
  XNOR2_X1 U390 ( .A(n488), .B(n486), .ZN(n617) );
  BUF_X1 U391 ( .A(G107), .Z(n455) );
  BUF_X1 U392 ( .A(G128), .Z(n461) );
  BUF_X1 U393 ( .A(G101), .Z(n459) );
  BUF_X2 U394 ( .A(n620), .Z(n793) );
  NOR2_X2 U395 ( .A1(n855), .A2(n856), .ZN(n710) );
  NAND2_X2 U396 ( .A1(n365), .A2(n369), .ZN(n855) );
  AND2_X2 U397 ( .A1(n501), .A2(n499), .ZN(n498) );
  AND2_X1 U398 ( .A1(n731), .A2(n730), .ZN(n420) );
  XNOR2_X2 U399 ( .A(n538), .B(n537), .ZN(n448) );
  NAND2_X2 U400 ( .A1(n830), .A2(n735), .ZN(n737) );
  XNOR2_X2 U401 ( .A(n617), .B(KEYINPUT1), .ZN(n690) );
  XNOR2_X1 U402 ( .A(G122), .B(G104), .ZN(n581) );
  NOR2_X1 U403 ( .A1(n361), .A2(n381), .ZN(n380) );
  NOR2_X1 U404 ( .A1(n360), .A2(n373), .ZN(n372) );
  AND2_X1 U405 ( .A1(n435), .A2(n635), .ZN(n434) );
  INV_X1 U406 ( .A(n390), .ZN(n782) );
  AND2_X1 U407 ( .A1(n358), .A2(n707), .ZN(n456) );
  NOR2_X1 U408 ( .A1(n427), .A2(n606), .ZN(n708) );
  NOR2_X1 U409 ( .A1(n638), .A2(n637), .ZN(n635) );
  AND2_X1 U410 ( .A1(n464), .A2(n494), .ZN(n463) );
  XNOR2_X1 U411 ( .A(n599), .B(n705), .ZN(n709) );
  NAND2_X1 U412 ( .A1(n380), .A2(n379), .ZN(n385) );
  NAND2_X1 U413 ( .A1(n372), .A2(n371), .ZN(n377) );
  NAND2_X1 U414 ( .A1(n404), .A2(n409), .ZN(n403) );
  XNOR2_X1 U415 ( .A(n364), .B(n363), .ZN(n762) );
  XNOR2_X1 U416 ( .A(n737), .B(n736), .ZN(n776) );
  XNOR2_X1 U417 ( .A(n737), .B(n736), .ZN(n393) );
  XNOR2_X1 U418 ( .A(n737), .B(n736), .ZN(n392) );
  XNOR2_X1 U419 ( .A(n647), .B(n469), .ZN(n672) );
  AND2_X1 U420 ( .A1(n437), .A2(n429), .ZN(n425) );
  AND2_X1 U421 ( .A1(n445), .A2(n400), .ZN(n443) );
  XNOR2_X1 U422 ( .A(n367), .B(n479), .ZN(n856) );
  NAND2_X1 U423 ( .A1(n456), .A2(n708), .ZN(n451) );
  NAND2_X1 U424 ( .A1(n370), .A2(n358), .ZN(n362) );
  AND2_X1 U425 ( .A1(n431), .A2(n778), .ZN(n370) );
  NAND2_X1 U426 ( .A1(n374), .A2(n761), .ZN(n373) );
  NAND2_X1 U427 ( .A1(n637), .A2(n638), .ZN(n781) );
  NAND2_X1 U428 ( .A1(n463), .A2(n462), .ZN(n687) );
  NOR2_X1 U429 ( .A1(n378), .A2(n376), .ZN(n375) );
  NAND2_X1 U430 ( .A1(n378), .A2(n376), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n536), .B(G478), .ZN(n615) );
  NAND2_X1 U432 ( .A1(n382), .A2(n761), .ZN(n381) );
  NAND2_X1 U433 ( .A1(n386), .A2(n384), .ZN(n382) );
  NOR2_X1 U434 ( .A1(n386), .A2(n384), .ZN(n383) );
  INV_X1 U435 ( .A(n760), .ZN(n363) );
  XNOR2_X1 U436 ( .A(n535), .B(n534), .ZN(n760) );
  XNOR2_X1 U437 ( .A(n522), .B(n473), .ZN(n638) );
  NAND2_X1 U438 ( .A1(n743), .A2(n742), .ZN(n761) );
  XNOR2_X1 U439 ( .A(G122), .B(G104), .ZN(n391) );
  XNOR2_X1 U440 ( .A(KEYINPUT68), .B(KEYINPUT19), .ZN(n604) );
  XNOR2_X1 U441 ( .A(G113), .B(G143), .ZN(n518) );
  INV_X2 U442 ( .A(KEYINPUT64), .ZN(n531) );
  XNOR2_X1 U443 ( .A(KEYINPUT71), .B(KEYINPUT48), .ZN(n713) );
  AND2_X1 U444 ( .A1(n423), .A2(n375), .ZN(n360) );
  AND2_X1 U445 ( .A1(n763), .A2(n383), .ZN(n361) );
  NAND2_X1 U446 ( .A1(n359), .A2(n761), .ZN(n454) );
  XNOR2_X1 U447 ( .A(n748), .B(n470), .ZN(n359) );
  INV_X1 U448 ( .A(n781), .ZN(n431) );
  NAND2_X1 U449 ( .A1(n422), .A2(G478), .ZN(n364) );
  AND2_X2 U450 ( .A1(n366), .A2(n477), .ZN(n365) );
  NAND2_X1 U451 ( .A1(n368), .A2(n476), .ZN(n366) );
  NAND2_X1 U452 ( .A1(n808), .A2(n480), .ZN(n367) );
  XNOR2_X1 U453 ( .A(n451), .B(KEYINPUT39), .ZN(n368) );
  NAND2_X1 U454 ( .A1(n716), .A2(n478), .ZN(n369) );
  NAND2_X1 U455 ( .A1(n703), .A2(n747), .ZN(n449) );
  OR2_X1 U456 ( .A1(n423), .A2(n752), .ZN(n371) );
  INV_X1 U457 ( .A(G210), .ZN(n376) );
  XNOR2_X1 U458 ( .A(n377), .B(n753), .ZN(G51) );
  INV_X1 U459 ( .A(n752), .ZN(n378) );
  OR2_X1 U460 ( .A1(n763), .A2(n741), .ZN(n379) );
  INV_X1 U461 ( .A(G475), .ZN(n384) );
  XNOR2_X1 U462 ( .A(n385), .B(n744), .ZN(G60) );
  INV_X1 U463 ( .A(n741), .ZN(n386) );
  BUF_X1 U464 ( .A(n556), .Z(n387) );
  BUF_X1 U465 ( .A(n605), .Z(n388) );
  BUF_X1 U466 ( .A(n693), .Z(n389) );
  NAND2_X1 U467 ( .A1(n715), .A2(n823), .ZN(n390) );
  NOR2_X1 U468 ( .A1(n420), .A2(n776), .ZN(n423) );
  NOR2_X4 U469 ( .A1(n738), .A2(n393), .ZN(n422) );
  AND2_X2 U470 ( .A1(n480), .A2(n390), .ZN(n394) );
  XNOR2_X2 U471 ( .A(n608), .B(KEYINPUT73), .ZN(n621) );
  XNOR2_X1 U472 ( .A(n451), .B(n450), .ZN(n716) );
  XNOR2_X1 U473 ( .A(KEYINPUT15), .B(G902), .ZN(n723) );
  NOR2_X1 U474 ( .A1(n672), .A2(n402), .ZN(n484) );
  INV_X1 U475 ( .A(n723), .ZN(n724) );
  INV_X1 U476 ( .A(KEYINPUT106), .ZN(n507) );
  INV_X1 U477 ( .A(KEYINPUT39), .ZN(n450) );
  XNOR2_X1 U478 ( .A(n546), .B(n487), .ZN(n486) );
  NAND2_X1 U479 ( .A1(n430), .A2(n572), .ZN(n488) );
  INV_X1 U480 ( .A(G469), .ZN(n487) );
  INV_X1 U481 ( .A(G472), .ZN(n408) );
  INV_X1 U482 ( .A(KEYINPUT40), .ZN(n478) );
  NAND2_X1 U483 ( .A1(n823), .A2(n478), .ZN(n477) );
  OR2_X1 U484 ( .A1(n688), .A2(n689), .ZN(n444) );
  INV_X1 U485 ( .A(n689), .ZN(n441) );
  XNOR2_X1 U486 ( .A(n574), .B(n573), .ZN(n427) );
  XNOR2_X1 U487 ( .A(n523), .B(G475), .ZN(n473) );
  INV_X1 U488 ( .A(n756), .ZN(n409) );
  INV_X1 U489 ( .A(G217), .ZN(n491) );
  XNOR2_X1 U490 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U491 ( .A(G146), .B(G137), .ZN(n564) );
  XOR2_X1 U492 ( .A(KEYINPUT5), .B(G116), .Z(n565) );
  NOR2_X1 U493 ( .A1(G953), .A2(G237), .ZN(n568) );
  INV_X1 U494 ( .A(G237), .ZN(n571) );
  XNOR2_X1 U495 ( .A(G113), .B(KEYINPUT76), .ZN(n465) );
  XNOR2_X1 U496 ( .A(G119), .B(KEYINPUT24), .ZN(n489) );
  XOR2_X1 U497 ( .A(KEYINPUT23), .B(G110), .Z(n551) );
  XOR2_X1 U498 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n513) );
  XNOR2_X1 U499 ( .A(G140), .B(G131), .ZN(n514) );
  XOR2_X1 U500 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n515) );
  NOR2_X1 U501 ( .A1(n770), .A2(n721), .ZN(n722) );
  XNOR2_X1 U502 ( .A(KEYINPUT4), .B(G131), .ZN(n537) );
  XNOR2_X1 U503 ( .A(n687), .B(n604), .ZN(n605) );
  NOR2_X1 U504 ( .A1(n790), .A2(n507), .ZN(n505) );
  XNOR2_X1 U505 ( .A(n755), .B(n754), .ZN(n756) );
  XNOR2_X1 U506 ( .A(KEYINPUT9), .B(KEYINPUT100), .ZN(n524) );
  XOR2_X1 U507 ( .A(KEYINPUT7), .B(KEYINPUT101), .Z(n525) );
  INV_X1 U508 ( .A(KEYINPUT102), .ZN(n472) );
  XOR2_X1 U509 ( .A(n455), .B(G110), .Z(n541) );
  XNOR2_X1 U510 ( .A(G146), .B(n459), .ZN(n542) );
  INV_X1 U511 ( .A(G953), .ZN(n829) );
  INV_X1 U512 ( .A(n823), .ZN(n508) );
  INV_X1 U513 ( .A(KEYINPUT108), .ZN(n510) );
  AND2_X1 U514 ( .A1(n407), .A2(n761), .ZN(n406) );
  NAND2_X1 U515 ( .A1(n409), .A2(n408), .ZN(n407) );
  XNOR2_X1 U516 ( .A(n740), .B(n739), .ZN(n741) );
  XNOR2_X1 U517 ( .A(n750), .B(n751), .ZN(n752) );
  NAND2_X1 U518 ( .A1(n442), .A2(n441), .ZN(n440) );
  INV_X1 U519 ( .A(KEYINPUT32), .ZN(n469) );
  INV_X1 U520 ( .A(n599), .ZN(n600) );
  INV_X1 U521 ( .A(KEYINPUT122), .ZN(n453) );
  XNOR2_X1 U522 ( .A(n672), .B(n468), .ZN(G21) );
  INV_X1 U523 ( .A(G119), .ZN(n468) );
  AND2_X1 U524 ( .A1(n568), .A2(G210), .ZN(n395) );
  AND2_X1 U525 ( .A1(n809), .A2(n483), .ZN(n396) );
  INV_X1 U526 ( .A(n612), .ZN(n471) );
  AND2_X1 U527 ( .A1(n646), .A2(n790), .ZN(n397) );
  AND2_X1 U528 ( .A1(n790), .A2(n507), .ZN(n398) );
  NAND2_X1 U529 ( .A1(n778), .A2(KEYINPUT92), .ZN(n399) );
  AND2_X1 U530 ( .A1(n444), .A2(n690), .ZN(n400) );
  INV_X1 U531 ( .A(G902), .ZN(n572) );
  INV_X1 U532 ( .A(n634), .ZN(n483) );
  XOR2_X1 U533 ( .A(KEYINPUT82), .B(KEYINPUT35), .Z(n401) );
  AND2_X1 U534 ( .A1(n676), .A2(KEYINPUT44), .ZN(n402) );
  OR2_X2 U535 ( .A1(n605), .A2(n631), .ZN(n633) );
  INV_X1 U536 ( .A(n422), .ZN(n404) );
  NAND2_X1 U537 ( .A1(n422), .A2(n411), .ZN(n410) );
  AND2_X1 U538 ( .A1(n756), .A2(G472), .ZN(n411) );
  XNOR2_X1 U539 ( .A(n412), .B(n757), .ZN(G57) );
  XNOR2_X1 U540 ( .A(n532), .B(n533), .ZN(n556) );
  XNOR2_X1 U541 ( .A(n530), .B(KEYINPUT89), .ZN(n533) );
  INV_X1 U542 ( .A(n677), .ZN(n413) );
  INV_X1 U543 ( .A(n722), .ZN(n414) );
  NAND2_X1 U544 ( .A1(n448), .A2(n566), .ZN(n417) );
  NAND2_X1 U545 ( .A1(n415), .A2(n416), .ZN(n418) );
  NAND2_X1 U546 ( .A1(n417), .A2(n418), .ZN(n452) );
  INV_X1 U547 ( .A(n448), .ZN(n415) );
  INV_X1 U548 ( .A(n566), .ZN(n416) );
  INV_X1 U549 ( .A(n773), .ZN(n419) );
  INV_X1 U550 ( .A(n770), .ZN(n830) );
  XNOR2_X1 U551 ( .A(n686), .B(n685), .ZN(n421) );
  XNOR2_X1 U552 ( .A(n686), .B(n685), .ZN(n447) );
  BUF_X2 U553 ( .A(n655), .Z(n656) );
  OR2_X1 U554 ( .A1(n706), .A2(n399), .ZN(n462) );
  XNOR2_X1 U555 ( .A(n493), .B(n560), .ZN(n424) );
  NOR2_X1 U556 ( .A1(n420), .A2(n776), .ZN(n763) );
  XNOR2_X1 U557 ( .A(n493), .B(n560), .ZN(n642) );
  NAND2_X1 U558 ( .A1(n470), .A2(n572), .ZN(n493) );
  NOR2_X1 U559 ( .A1(n392), .A2(n491), .ZN(n490) );
  INV_X1 U560 ( .A(n648), .ZN(n502) );
  NAND2_X1 U561 ( .A1(n425), .A2(n434), .ZN(n439) );
  NAND2_X2 U562 ( .A1(n443), .A2(n440), .ZN(n747) );
  NAND2_X1 U563 ( .A1(n414), .A2(n733), .ZN(n725) );
  NOR2_X1 U564 ( .A1(n758), .A2(n428), .ZN(n671) );
  NAND2_X1 U565 ( .A1(n485), .A2(n484), .ZN(n428) );
  XNOR2_X2 U566 ( .A(n652), .B(KEYINPUT107), .ZN(n758) );
  NAND2_X1 U567 ( .A1(n396), .A2(n656), .ZN(n429) );
  INV_X1 U568 ( .A(n765), .ZN(n430) );
  XNOR2_X1 U569 ( .A(n545), .B(n844), .ZN(n765) );
  NAND2_X1 U570 ( .A1(n358), .A2(n778), .ZN(n432) );
  NOR2_X1 U571 ( .A1(n782), .A2(n432), .ZN(n783) );
  NAND2_X1 U572 ( .A1(n394), .A2(n612), .ZN(n698) );
  NAND2_X1 U573 ( .A1(n433), .A2(n394), .ZN(n692) );
  NAND2_X1 U574 ( .A1(n436), .A2(n634), .ZN(n435) );
  INV_X1 U575 ( .A(n809), .ZN(n436) );
  NAND2_X1 U576 ( .A1(n438), .A2(n634), .ZN(n437) );
  INV_X1 U577 ( .A(n656), .ZN(n438) );
  XNOR2_X2 U578 ( .A(n439), .B(n401), .ZN(n854) );
  INV_X1 U579 ( .A(n447), .ZN(n442) );
  NAND2_X1 U580 ( .A1(n421), .A2(n446), .ZN(n445) );
  AND2_X1 U581 ( .A1(n688), .A2(n689), .ZN(n446) );
  XNOR2_X1 U582 ( .A(n448), .B(n539), .ZN(n844) );
  XNOR2_X1 U583 ( .A(n449), .B(n704), .ZN(n712) );
  XNOR2_X2 U584 ( .A(n452), .B(n569), .ZN(n755) );
  NAND2_X1 U585 ( .A1(n492), .A2(n490), .ZN(n748) );
  XNOR2_X1 U586 ( .A(n454), .B(n453), .ZN(G66) );
  NAND2_X1 U587 ( .A1(n506), .A2(n504), .ZN(n503) );
  NAND2_X1 U588 ( .A1(n503), .A2(n649), .ZN(n501) );
  NAND2_X1 U589 ( .A1(n457), .A2(n497), .ZN(n495) );
  INV_X1 U590 ( .A(n458), .ZN(n457) );
  NAND2_X1 U591 ( .A1(n496), .A2(KEYINPUT66), .ZN(n458) );
  BUF_X2 U592 ( .A(n706), .Z(n599) );
  NAND2_X1 U593 ( .A1(n556), .A2(G221), .ZN(n482) );
  XNOR2_X2 U594 ( .A(n620), .B(n619), .ZN(n665) );
  NAND2_X1 U595 ( .A1(n706), .A2(n603), .ZN(n464) );
  XNOR2_X2 U596 ( .A(n474), .B(n598), .ZN(n706) );
  XNOR2_X2 U597 ( .A(n466), .B(n465), .ZN(n586) );
  XNOR2_X2 U598 ( .A(n467), .B(n567), .ZN(n466) );
  XNOR2_X2 U599 ( .A(G119), .B(G101), .ZN(n467) );
  XNOR2_X2 U600 ( .A(n481), .B(n555), .ZN(n470) );
  NAND2_X1 U601 ( .A1(n480), .A2(n612), .ZN(n693) );
  XNOR2_X1 U602 ( .A(n538), .B(n472), .ZN(n529) );
  XNOR2_X2 U603 ( .A(n593), .B(G134), .ZN(n538) );
  XNOR2_X2 U604 ( .A(G143), .B(G128), .ZN(n593) );
  INV_X1 U605 ( .A(n615), .ZN(n637) );
  XNOR2_X1 U606 ( .A(n826), .B(n661), .ZN(n715) );
  NAND2_X1 U607 ( .A1(n615), .A2(n638), .ZN(n826) );
  OR2_X2 U608 ( .A1(n749), .A2(n724), .ZN(n474) );
  XNOR2_X1 U609 ( .A(n836), .B(n475), .ZN(n749) );
  XNOR2_X1 U610 ( .A(n595), .B(n596), .ZN(n475) );
  XNOR2_X1 U611 ( .A(n586), .B(n587), .ZN(n836) );
  NOR2_X1 U612 ( .A1(n823), .A2(n478), .ZN(n476) );
  XNOR2_X1 U613 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n479) );
  AND2_X2 U614 ( .A1(n611), .A2(n617), .ZN(n480) );
  XNOR2_X2 U615 ( .A(n482), .B(n843), .ZN(n481) );
  NAND2_X1 U616 ( .A1(n636), .A2(n676), .ZN(n485) );
  XNOR2_X1 U617 ( .A(n489), .B(n461), .ZN(n548) );
  INV_X1 U618 ( .A(n738), .ZN(n492) );
  NAND2_X1 U619 ( .A1(n618), .A2(n603), .ZN(n494) );
  NAND2_X1 U620 ( .A1(n495), .A2(n498), .ZN(n651) );
  NAND2_X1 U621 ( .A1(n502), .A2(KEYINPUT106), .ZN(n496) );
  INV_X1 U622 ( .A(n503), .ZN(n497) );
  NAND2_X1 U623 ( .A1(n502), .A2(n500), .ZN(n499) );
  AND2_X1 U624 ( .A1(n649), .A2(KEYINPUT106), .ZN(n500) );
  NAND2_X1 U625 ( .A1(n648), .A2(n398), .ZN(n506) );
  XNOR2_X2 U626 ( .A(G146), .B(G125), .ZN(n589) );
  NAND2_X2 U627 ( .A1(n509), .A2(n508), .ZN(n686) );
  XNOR2_X2 U628 ( .A(n511), .B(n510), .ZN(n509) );
  NAND2_X1 U629 ( .A1(n621), .A2(n665), .ZN(n511) );
  INV_X1 U630 ( .A(KEYINPUT80), .ZN(n736) );
  AND2_X1 U631 ( .A1(n708), .A2(n600), .ZN(n601) );
  NAND2_X1 U632 ( .A1(n602), .A2(n601), .ZN(n699) );
  XNOR2_X1 U633 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n523) );
  NAND2_X1 U634 ( .A1(n568), .A2(G214), .ZN(n512) );
  XNOR2_X1 U635 ( .A(n513), .B(n512), .ZN(n517) );
  XNOR2_X1 U636 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U637 ( .A(n517), .B(n516), .ZN(n521) );
  XNOR2_X1 U638 ( .A(n589), .B(KEYINPUT10), .ZN(n843) );
  XNOR2_X1 U639 ( .A(n391), .B(n518), .ZN(n519) );
  XNOR2_X1 U640 ( .A(n843), .B(n519), .ZN(n520) );
  XNOR2_X1 U641 ( .A(n521), .B(n520), .ZN(n740) );
  NOR2_X1 U642 ( .A1(G902), .A2(n740), .ZN(n522) );
  XNOR2_X1 U643 ( .A(n525), .B(n524), .ZN(n527) );
  XNOR2_X2 U644 ( .A(G116), .B(G107), .ZN(n582) );
  XNOR2_X1 U645 ( .A(n582), .B(G122), .ZN(n526) );
  XNOR2_X1 U646 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U647 ( .A(n529), .B(n528), .ZN(n535) );
  XNOR2_X2 U648 ( .A(KEYINPUT8), .B(KEYINPUT70), .ZN(n530) );
  XNOR2_X2 U649 ( .A(n531), .B(G953), .ZN(n845) );
  NAND2_X1 U650 ( .A1(n845), .A2(G234), .ZN(n532) );
  NAND2_X1 U651 ( .A1(n387), .A2(G217), .ZN(n534) );
  NAND2_X1 U652 ( .A1(n760), .A2(n572), .ZN(n536) );
  XNOR2_X1 U653 ( .A(KEYINPUT75), .B(KEYINPUT74), .ZN(n546) );
  XNOR2_X1 U654 ( .A(G140), .B(G137), .ZN(n547) );
  INV_X1 U655 ( .A(n547), .ZN(n539) );
  NAND2_X1 U656 ( .A1(n460), .A2(G227), .ZN(n540) );
  XOR2_X1 U657 ( .A(n541), .B(n540), .Z(n544) );
  XNOR2_X1 U658 ( .A(n542), .B(G104), .ZN(n543) );
  XNOR2_X1 U659 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U660 ( .A(n548), .B(n547), .ZN(n552) );
  INV_X1 U661 ( .A(n552), .ZN(n550) );
  INV_X1 U662 ( .A(n551), .ZN(n549) );
  NAND2_X1 U663 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U664 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U665 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U666 ( .A1(n723), .A2(G234), .ZN(n557) );
  XNOR2_X1 U667 ( .A(n557), .B(KEYINPUT20), .ZN(n558) );
  XNOR2_X1 U668 ( .A(n558), .B(KEYINPUT96), .ZN(n561) );
  NAND2_X1 U669 ( .A1(n561), .A2(G217), .ZN(n559) );
  XNOR2_X1 U670 ( .A(n559), .B(KEYINPUT25), .ZN(n560) );
  NAND2_X1 U671 ( .A1(n561), .A2(G221), .ZN(n562) );
  XNOR2_X1 U672 ( .A(n562), .B(KEYINPUT21), .ZN(n786) );
  OR2_X2 U673 ( .A1(n424), .A2(n786), .ZN(n789) );
  INV_X1 U674 ( .A(n789), .ZN(n563) );
  AND2_X2 U675 ( .A1(n617), .A2(n563), .ZN(n707) );
  AND2_X1 U676 ( .A1(n635), .A2(n707), .ZN(n602) );
  XNOR2_X2 U677 ( .A(KEYINPUT93), .B(KEYINPUT3), .ZN(n567) );
  XNOR2_X1 U678 ( .A(n586), .B(n395), .ZN(n569) );
  NAND2_X1 U679 ( .A1(n755), .A2(n572), .ZN(n570) );
  XNOR2_X2 U680 ( .A(n570), .B(G472), .ZN(n620) );
  NAND2_X1 U681 ( .A1(n572), .A2(n571), .ZN(n597) );
  NAND2_X1 U682 ( .A1(n597), .A2(G214), .ZN(n778) );
  NAND2_X1 U683 ( .A1(n620), .A2(n778), .ZN(n574) );
  XOR2_X1 U684 ( .A(KEYINPUT109), .B(KEYINPUT30), .Z(n573) );
  NAND2_X1 U685 ( .A1(G237), .A2(G234), .ZN(n575) );
  XNOR2_X1 U686 ( .A(n575), .B(KEYINPUT14), .ZN(n577) );
  NAND2_X1 U687 ( .A1(G952), .A2(n577), .ZN(n576) );
  XNOR2_X1 U688 ( .A(KEYINPUT95), .B(n576), .ZN(n806) );
  NAND2_X1 U689 ( .A1(n806), .A2(n829), .ZN(n630) );
  AND2_X1 U690 ( .A1(G902), .A2(n577), .ZN(n628) );
  NOR2_X1 U691 ( .A1(n460), .A2(G900), .ZN(n578) );
  NAND2_X1 U692 ( .A1(n628), .A2(n578), .ZN(n579) );
  NAND2_X1 U693 ( .A1(n630), .A2(n579), .ZN(n580) );
  XNOR2_X1 U694 ( .A(n580), .B(KEYINPUT85), .ZN(n606) );
  XNOR2_X1 U695 ( .A(n582), .B(n581), .ZN(n585) );
  XNOR2_X1 U696 ( .A(KEYINPUT78), .B(KEYINPUT16), .ZN(n583) );
  XNOR2_X1 U697 ( .A(n583), .B(G110), .ZN(n584) );
  XNOR2_X1 U698 ( .A(n585), .B(n584), .ZN(n587) );
  XNOR2_X1 U699 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n588) );
  XNOR2_X1 U700 ( .A(n589), .B(n588), .ZN(n592) );
  XNOR2_X1 U701 ( .A(KEYINPUT94), .B(KEYINPUT4), .ZN(n590) );
  XNOR2_X1 U702 ( .A(n590), .B(KEYINPUT81), .ZN(n591) );
  XNOR2_X1 U703 ( .A(n592), .B(n591), .ZN(n596) );
  NAND2_X1 U704 ( .A1(n845), .A2(G224), .ZN(n594) );
  XNOR2_X1 U705 ( .A(n593), .B(n594), .ZN(n595) );
  NAND2_X1 U706 ( .A1(n597), .A2(G210), .ZN(n598) );
  XNOR2_X1 U707 ( .A(n699), .B(G143), .ZN(G45) );
  INV_X1 U708 ( .A(n778), .ZN(n618) );
  INV_X1 U709 ( .A(KEYINPUT92), .ZN(n603) );
  INV_X1 U710 ( .A(n388), .ZN(n612) );
  NOR2_X1 U711 ( .A1(n786), .A2(n606), .ZN(n607) );
  NAND2_X1 U712 ( .A1(n642), .A2(n607), .ZN(n608) );
  NAND2_X1 U713 ( .A1(n621), .A2(n793), .ZN(n610) );
  XOR2_X1 U714 ( .A(KEYINPUT28), .B(KEYINPUT110), .Z(n609) );
  XNOR2_X1 U715 ( .A(n610), .B(n609), .ZN(n611) );
  NOR2_X1 U716 ( .A1(n389), .A2(n826), .ZN(n614) );
  XNOR2_X1 U717 ( .A(n461), .B(KEYINPUT29), .ZN(n613) );
  XNOR2_X1 U718 ( .A(n614), .B(n613), .ZN(G30) );
  OR2_X1 U719 ( .A1(n638), .A2(n615), .ZN(n823) );
  NOR2_X1 U720 ( .A1(n389), .A2(n823), .ZN(n616) );
  XOR2_X1 U721 ( .A(G146), .B(n616), .Z(G48) );
  OR2_X1 U722 ( .A1(n690), .A2(n618), .ZN(n622) );
  INV_X1 U723 ( .A(KEYINPUT6), .ZN(n619) );
  NOR2_X1 U724 ( .A1(n622), .A2(n686), .ZN(n624) );
  INV_X1 U725 ( .A(KEYINPUT43), .ZN(n623) );
  XNOR2_X1 U726 ( .A(n624), .B(n623), .ZN(n625) );
  AND2_X1 U727 ( .A1(n599), .A2(n625), .ZN(n717) );
  XOR2_X1 U728 ( .A(G140), .B(n717), .Z(G42) );
  INV_X1 U729 ( .A(n789), .ZN(n653) );
  AND2_X1 U730 ( .A1(n665), .A2(n653), .ZN(n626) );
  NAND2_X1 U731 ( .A1(n626), .A2(n690), .ZN(n627) );
  XNOR2_X2 U732 ( .A(n627), .B(KEYINPUT33), .ZN(n809) );
  NOR2_X1 U733 ( .A1(G898), .A2(n829), .ZN(n840) );
  NAND2_X1 U734 ( .A1(n840), .A2(n628), .ZN(n629) );
  AND2_X1 U735 ( .A1(n630), .A2(n629), .ZN(n631) );
  INV_X1 U736 ( .A(KEYINPUT0), .ZN(n632) );
  XNOR2_X2 U737 ( .A(n633), .B(n632), .ZN(n655) );
  XOR2_X1 U738 ( .A(KEYINPUT34), .B(KEYINPUT83), .Z(n634) );
  XNOR2_X1 U739 ( .A(n854), .B(KEYINPUT69), .ZN(n636) );
  INV_X1 U740 ( .A(KEYINPUT65), .ZN(n676) );
  NOR2_X1 U741 ( .A1(n781), .A2(n786), .ZN(n639) );
  NAND2_X1 U742 ( .A1(n655), .A2(n639), .ZN(n641) );
  XNOR2_X2 U743 ( .A(n641), .B(n640), .ZN(n648) );
  BUF_X1 U744 ( .A(n648), .Z(n646) );
  BUF_X1 U745 ( .A(n424), .Z(n650) );
  XOR2_X1 U746 ( .A(KEYINPUT105), .B(n650), .Z(n787) );
  NAND2_X1 U747 ( .A1(n690), .A2(n787), .ZN(n644) );
  XNOR2_X1 U748 ( .A(n665), .B(KEYINPUT84), .ZN(n643) );
  NOR2_X1 U749 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U750 ( .A1(n646), .A2(n645), .ZN(n647) );
  INV_X1 U751 ( .A(n690), .ZN(n790) );
  INV_X1 U752 ( .A(KEYINPUT66), .ZN(n649) );
  NAND2_X1 U753 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U754 ( .A1(n690), .A2(n653), .ZN(n654) );
  NAND2_X1 U755 ( .A1(n654), .A2(n793), .ZN(n797) );
  INV_X1 U756 ( .A(n656), .ZN(n657) );
  XNOR2_X1 U757 ( .A(n658), .B(KEYINPUT31), .ZN(n825) );
  INV_X1 U758 ( .A(n707), .ZN(n659) );
  NOR2_X1 U759 ( .A1(n659), .A2(n793), .ZN(n660) );
  NAND2_X1 U760 ( .A1(n656), .A2(n660), .ZN(n820) );
  NAND2_X1 U761 ( .A1(n825), .A2(n820), .ZN(n663) );
  INV_X1 U762 ( .A(KEYINPUT103), .ZN(n661) );
  XNOR2_X1 U763 ( .A(KEYINPUT87), .B(n782), .ZN(n662) );
  NAND2_X1 U764 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U765 ( .A(n664), .B(KEYINPUT104), .ZN(n669) );
  NOR2_X1 U766 ( .A1(n665), .A2(n787), .ZN(n666) );
  AND2_X1 U767 ( .A1(n397), .A2(n666), .ZN(n816) );
  NOR2_X1 U768 ( .A1(KEYINPUT44), .A2(n676), .ZN(n667) );
  NOR2_X1 U769 ( .A1(n816), .A2(n667), .ZN(n668) );
  NAND2_X1 U770 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U771 ( .A1(n671), .A2(n670), .ZN(n682) );
  INV_X1 U772 ( .A(n758), .ZN(n675) );
  NOR2_X1 U773 ( .A1(n672), .A2(KEYINPUT69), .ZN(n673) );
  AND2_X1 U774 ( .A1(n413), .A2(n673), .ZN(n674) );
  NAND2_X1 U775 ( .A1(n675), .A2(n674), .ZN(n680) );
  INV_X1 U776 ( .A(n854), .ZN(n677) );
  OR2_X1 U777 ( .A1(n677), .A2(n676), .ZN(n678) );
  AND2_X1 U778 ( .A1(n678), .A2(KEYINPUT44), .ZN(n679) );
  NAND2_X1 U779 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U780 ( .A1(n682), .A2(n681), .ZN(n684) );
  INV_X1 U781 ( .A(KEYINPUT45), .ZN(n683) );
  XNOR2_X2 U782 ( .A(n684), .B(n683), .ZN(n770) );
  INV_X1 U783 ( .A(KEYINPUT112), .ZN(n685) );
  BUF_X1 U784 ( .A(n687), .Z(n688) );
  XNOR2_X1 U785 ( .A(KEYINPUT113), .B(KEYINPUT36), .ZN(n689) );
  INV_X1 U786 ( .A(KEYINPUT87), .ZN(n691) );
  NAND2_X1 U787 ( .A1(n692), .A2(n691), .ZN(n697) );
  INV_X1 U788 ( .A(n693), .ZN(n694) );
  NAND2_X1 U789 ( .A1(n694), .A2(n782), .ZN(n695) );
  NAND2_X1 U790 ( .A1(n695), .A2(KEYINPUT87), .ZN(n696) );
  NAND2_X1 U791 ( .A1(n697), .A2(n696), .ZN(n702) );
  NAND2_X1 U792 ( .A1(n698), .A2(KEYINPUT47), .ZN(n701) );
  XNOR2_X1 U793 ( .A(n699), .B(KEYINPUT88), .ZN(n700) );
  INV_X1 U794 ( .A(KEYINPUT72), .ZN(n704) );
  INV_X1 U795 ( .A(KEYINPUT38), .ZN(n705) );
  XNOR2_X1 U796 ( .A(n710), .B(KEYINPUT46), .ZN(n711) );
  NAND2_X1 U797 ( .A1(n712), .A2(n711), .ZN(n714) );
  XNOR2_X1 U798 ( .A(n714), .B(n713), .ZN(n719) );
  NOR2_X1 U799 ( .A1(n716), .A2(n715), .ZN(n828) );
  NOR2_X1 U800 ( .A1(n828), .A2(n717), .ZN(n718) );
  NAND2_X2 U801 ( .A1(n719), .A2(n718), .ZN(n732) );
  INV_X1 U802 ( .A(KEYINPUT91), .ZN(n720) );
  XNOR2_X2 U803 ( .A(n732), .B(n720), .ZN(n771) );
  XNOR2_X1 U804 ( .A(n771), .B(KEYINPUT79), .ZN(n726) );
  NAND2_X1 U805 ( .A1(n726), .A2(KEYINPUT90), .ZN(n721) );
  NAND2_X1 U806 ( .A1(n725), .A2(n724), .ZN(n731) );
  NAND2_X1 U807 ( .A1(n726), .A2(n724), .ZN(n727) );
  NOR2_X1 U808 ( .A1(n770), .A2(n727), .ZN(n728) );
  NOR2_X1 U809 ( .A1(n728), .A2(KEYINPUT90), .ZN(n729) );
  INV_X1 U810 ( .A(n729), .ZN(n730) );
  AND2_X2 U811 ( .A1(n731), .A2(n730), .ZN(n738) );
  BUF_X1 U812 ( .A(n732), .Z(n734) );
  INV_X1 U813 ( .A(KEYINPUT2), .ZN(n733) );
  NOR2_X1 U814 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U815 ( .A(KEYINPUT67), .B(KEYINPUT59), .Z(n739) );
  INV_X1 U816 ( .A(n460), .ZN(n743) );
  INV_X1 U817 ( .A(G952), .ZN(n742) );
  INV_X1 U818 ( .A(KEYINPUT60), .ZN(n744) );
  XOR2_X1 U819 ( .A(KEYINPUT37), .B(KEYINPUT117), .Z(n745) );
  XOR2_X1 U820 ( .A(n745), .B(G125), .Z(n746) );
  XNOR2_X1 U821 ( .A(n747), .B(n746), .ZN(G27) );
  BUF_X1 U822 ( .A(n749), .Z(n750) );
  XNOR2_X1 U823 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n751) );
  INV_X1 U824 ( .A(KEYINPUT56), .ZN(n753) );
  XNOR2_X1 U825 ( .A(KEYINPUT114), .B(KEYINPUT62), .ZN(n754) );
  XOR2_X1 U826 ( .A(KEYINPUT115), .B(KEYINPUT63), .Z(n757) );
  BUF_X1 U827 ( .A(n758), .Z(n759) );
  XOR2_X1 U828 ( .A(n759), .B(G110), .Z(G12) );
  INV_X1 U829 ( .A(n761), .ZN(n768) );
  NOR2_X1 U830 ( .A1(n762), .A2(n768), .ZN(G63) );
  NAND2_X1 U831 ( .A1(n422), .A2(G469), .ZN(n767) );
  XOR2_X1 U832 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n764) );
  XNOR2_X1 U833 ( .A(n765), .B(n764), .ZN(n766) );
  XNOR2_X1 U834 ( .A(n767), .B(n766), .ZN(n769) );
  NOR2_X1 U835 ( .A1(n769), .A2(n768), .ZN(G54) );
  BUF_X1 U836 ( .A(n770), .Z(n773) );
  BUF_X1 U837 ( .A(n771), .Z(n772) );
  NOR2_X1 U838 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U839 ( .A1(n774), .A2(KEYINPUT2), .ZN(n775) );
  XNOR2_X1 U840 ( .A(n775), .B(KEYINPUT86), .ZN(n777) );
  NOR2_X1 U841 ( .A1(n777), .A2(n392), .ZN(n814) );
  NOR2_X1 U842 ( .A1(n358), .A2(n778), .ZN(n779) );
  XOR2_X1 U843 ( .A(KEYINPUT121), .B(n779), .Z(n780) );
  NOR2_X1 U844 ( .A1(n781), .A2(n780), .ZN(n784) );
  NOR2_X1 U845 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U846 ( .A1(n436), .A2(n785), .ZN(n804) );
  AND2_X1 U847 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U848 ( .A(KEYINPUT49), .B(n788), .ZN(n795) );
  NAND2_X1 U849 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U850 ( .A(KEYINPUT50), .B(n791), .Z(n792) );
  NOR2_X1 U851 ( .A1(n793), .A2(n792), .ZN(n794) );
  NAND2_X1 U852 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U853 ( .A(n796), .B(KEYINPUT118), .ZN(n798) );
  NAND2_X1 U854 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U855 ( .A(n799), .B(KEYINPUT51), .ZN(n800) );
  XNOR2_X1 U856 ( .A(n800), .B(KEYINPUT119), .ZN(n801) );
  NAND2_X1 U857 ( .A1(n801), .A2(n808), .ZN(n802) );
  XOR2_X1 U858 ( .A(KEYINPUT120), .B(n802), .Z(n803) );
  NOR2_X1 U859 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U860 ( .A(KEYINPUT52), .B(n805), .Z(n807) );
  NAND2_X1 U861 ( .A1(n807), .A2(n806), .ZN(n812) );
  NAND2_X1 U862 ( .A1(n809), .A2(n808), .ZN(n810) );
  AND2_X1 U863 ( .A1(n810), .A2(n829), .ZN(n811) );
  NAND2_X1 U864 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U865 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U866 ( .A(n815), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U867 ( .A(n459), .B(n816), .Z(G3) );
  NOR2_X1 U868 ( .A1(n820), .A2(n823), .ZN(n817) );
  XOR2_X1 U869 ( .A(G104), .B(n817), .Z(G6) );
  XOR2_X1 U870 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n819) );
  XNOR2_X1 U871 ( .A(n455), .B(KEYINPUT116), .ZN(n818) );
  XNOR2_X1 U872 ( .A(n819), .B(n818), .ZN(n822) );
  NOR2_X1 U873 ( .A1(n820), .A2(n826), .ZN(n821) );
  XOR2_X1 U874 ( .A(n822), .B(n821), .Z(G9) );
  NOR2_X1 U875 ( .A1(n823), .A2(n825), .ZN(n824) );
  XOR2_X1 U876 ( .A(G113), .B(n824), .Z(G15) );
  NOR2_X1 U877 ( .A1(n826), .A2(n825), .ZN(n827) );
  XOR2_X1 U878 ( .A(G116), .B(n827), .Z(G18) );
  XOR2_X1 U879 ( .A(G134), .B(n828), .Z(G36) );
  NAND2_X1 U880 ( .A1(n419), .A2(n829), .ZN(n834) );
  NAND2_X1 U881 ( .A1(G953), .A2(G224), .ZN(n831) );
  XNOR2_X1 U882 ( .A(KEYINPUT61), .B(n831), .ZN(n832) );
  NAND2_X1 U883 ( .A1(n832), .A2(G898), .ZN(n833) );
  NAND2_X1 U884 ( .A1(n834), .A2(n833), .ZN(n835) );
  XNOR2_X1 U885 ( .A(n835), .B(KEYINPUT125), .ZN(n842) );
  BUF_X1 U886 ( .A(n836), .Z(n837) );
  XNOR2_X1 U887 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n838) );
  XNOR2_X1 U888 ( .A(n837), .B(n838), .ZN(n839) );
  NOR2_X1 U889 ( .A1(n840), .A2(n839), .ZN(n841) );
  XOR2_X1 U890 ( .A(n842), .B(n841), .Z(G69) );
  XNOR2_X1 U891 ( .A(n844), .B(n843), .ZN(n847) );
  XNOR2_X1 U892 ( .A(n772), .B(n847), .ZN(n846) );
  NAND2_X1 U893 ( .A1(n846), .A2(n460), .ZN(n852) );
  XNOR2_X1 U894 ( .A(n847), .B(G227), .ZN(n848) );
  NAND2_X1 U895 ( .A1(n848), .A2(G900), .ZN(n849) );
  XNOR2_X1 U896 ( .A(n849), .B(KEYINPUT126), .ZN(n850) );
  NAND2_X1 U897 ( .A1(n850), .A2(G953), .ZN(n851) );
  NAND2_X1 U898 ( .A1(n852), .A2(n851), .ZN(n853) );
  XOR2_X1 U899 ( .A(KEYINPUT127), .B(n853), .Z(G72) );
  XNOR2_X1 U900 ( .A(n413), .B(G122), .ZN(G24) );
  XOR2_X1 U901 ( .A(n855), .B(G131), .Z(G33) );
  XOR2_X1 U902 ( .A(n856), .B(G137), .Z(G39) );
endmodule

