//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT71), .B(G237), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G210), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n190), .B(KEYINPUT27), .Z(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT72), .ZN(new_n192));
  XOR2_X1   g006(.A(KEYINPUT26), .B(G101), .Z(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT73), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n192), .B(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(G143), .B(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  OR2_X1    g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n199), .A2(new_n197), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n198), .B1(new_n200), .B2(new_n196), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G137), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT11), .B1(new_n203), .B2(G134), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(G134), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT64), .A2(G137), .ZN(new_n208));
  NOR2_X1   g022(.A1(KEYINPUT64), .A2(G137), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT11), .A2(G134), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n207), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  NOR4_X1   g027(.A1(new_n208), .A2(new_n209), .A3(new_n211), .A4(KEYINPUT65), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n206), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G131), .ZN(new_n216));
  XOR2_X1   g030(.A(KEYINPUT66), .B(G131), .Z(new_n217));
  OAI211_X1 g031(.A(new_n206), .B(new_n217), .C1(new_n213), .C2(new_n214), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n202), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G143), .ZN(new_n221));
  INV_X1    g035(.A(G143), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n225), .A3(G128), .ZN(new_n226));
  INV_X1    g040(.A(G128), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n221), .B(new_n223), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G131), .ZN(new_n230));
  INV_X1    g044(.A(G134), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(new_n208), .B2(new_n209), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n230), .B1(new_n232), .B2(new_n205), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n218), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n219), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT2), .B(G113), .ZN(new_n238));
  INV_X1    g052(.A(G116), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(G119), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT70), .B(G116), .ZN(new_n242));
  INV_X1    g056(.A(G119), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n238), .B1(new_n245), .B2(KEYINPUT69), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n247));
  INV_X1    g061(.A(new_n238), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n244), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n237), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT28), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n235), .B1(new_n219), .B2(KEYINPUT67), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n256));
  AOI211_X1 g070(.A(new_n256), .B(new_n202), .C1(new_n216), .C2(new_n218), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n250), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n258), .A2(new_n252), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n195), .B(new_n254), .C1(new_n259), .C2(new_n253), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT29), .B1(new_n260), .B2(KEYINPUT75), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT30), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n262), .B1(new_n255), .B2(new_n257), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT68), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n265), .B(new_n262), .C1(new_n255), .C2(new_n257), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n237), .A2(KEYINPUT30), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n264), .A2(new_n250), .A3(new_n266), .A4(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n252), .ZN(new_n269));
  INV_X1    g083(.A(new_n195), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n261), .B(new_n271), .C1(KEYINPUT75), .C2(new_n260), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n250), .B1(new_n219), .B2(new_n236), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n252), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT28), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n195), .A2(KEYINPUT29), .A3(new_n254), .A4(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT76), .ZN(new_n277));
  INV_X1    g091(.A(G902), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n277), .B1(new_n276), .B2(new_n278), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n187), .B1(new_n272), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT32), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n268), .A2(new_n195), .A3(new_n252), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(KEYINPUT74), .A3(KEYINPUT31), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n254), .B1(new_n259), .B2(new_n253), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n270), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT31), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n268), .A2(new_n291), .A3(new_n195), .A4(new_n252), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT74), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n285), .A2(KEYINPUT31), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(G902), .B1(new_n290), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n284), .B1(new_n296), .B2(new_n187), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n288), .A3(new_n286), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n298), .A2(new_n284), .A3(new_n187), .A4(new_n278), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n283), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT77), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT16), .ZN(new_n303));
  INV_X1    g117(.A(G140), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(G125), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n305), .B(KEYINPUT80), .ZN(new_n306));
  NAND2_X1  g120(.A1(KEYINPUT79), .A2(G125), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(new_n304), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT16), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(new_n309), .A3(G146), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT81), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n306), .A2(new_n309), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n220), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT81), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n306), .A2(new_n309), .A3(new_n314), .A4(G146), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n311), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n317), .B1(new_n243), .B2(G128), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n227), .A2(KEYINPUT23), .A3(G119), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n318), .B(new_n319), .C1(G119), .C2(new_n227), .ZN(new_n320));
  XNOR2_X1  g134(.A(G119), .B(G128), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT24), .B(G110), .Z(new_n322));
  AOI22_X1  g136(.A1(new_n320), .A2(G110), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n316), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(G125), .B(G140), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n220), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(KEYINPUT82), .ZN(new_n327));
  OAI22_X1  g141(.A1(new_n320), .A2(G110), .B1(new_n321), .B2(new_n322), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n310), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  XOR2_X1   g144(.A(KEYINPUT22), .B(G137), .Z(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT83), .ZN(new_n332));
  INV_X1    g146(.A(G953), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n333), .A2(G221), .A3(G234), .ZN(new_n334));
  XOR2_X1   g148(.A(new_n332), .B(new_n334), .Z(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n330), .B(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n278), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n339), .A2(KEYINPUT25), .ZN(new_n340));
  INV_X1    g154(.A(G217), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n341), .B1(G234), .B2(new_n278), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT78), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n343), .B1(new_n339), .B2(KEYINPUT25), .ZN(new_n344));
  OR2_X1    g158(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n343), .A2(G902), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n338), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n293), .A2(new_n294), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n187), .B(new_n278), .C1(new_n350), .C2(new_n289), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT32), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n299), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n283), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n189), .A2(G214), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n222), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n189), .A2(G143), .A3(G214), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(KEYINPUT18), .A2(G131), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n357), .A2(KEYINPUT18), .A3(G131), .A4(new_n358), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n327), .B1(new_n220), .B2(new_n308), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(G113), .B(G122), .ZN(new_n366));
  INV_X1    g180(.A(G104), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n366), .B(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(KEYINPUT95), .ZN(new_n369));
  INV_X1    g183(.A(new_n217), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n359), .A2(KEYINPUT17), .A3(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n371), .A2(new_n311), .A3(new_n315), .A4(new_n313), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n357), .A2(new_n217), .A3(new_n358), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n217), .B1(new_n357), .B2(new_n358), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n374), .A2(KEYINPUT17), .A3(new_n375), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n365), .B(new_n369), .C1(new_n372), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n278), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n316), .B1(KEYINPUT17), .B2(new_n375), .ZN(new_n379));
  INV_X1    g193(.A(new_n375), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT17), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(new_n373), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n369), .B1(new_n383), .B2(new_n365), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT96), .B1(new_n378), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n365), .B1(new_n372), .B2(new_n376), .ZN(new_n386));
  INV_X1    g200(.A(new_n369), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT96), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n388), .A2(new_n389), .A3(new_n278), .A4(new_n377), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n385), .A2(G475), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n308), .A2(KEYINPUT19), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(KEYINPUT19), .B2(new_n325), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n220), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n310), .B(new_n394), .C1(new_n374), .C2(new_n375), .ZN(new_n395));
  INV_X1    g209(.A(new_n368), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n365), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(G475), .A2(G902), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n379), .A2(new_n382), .B1(new_n364), .B2(new_n363), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n397), .B(new_n398), .C1(new_n399), .C2(new_n396), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT20), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n386), .A2(new_n368), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT20), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n402), .A2(new_n403), .A3(new_n397), .A4(new_n398), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n391), .A2(new_n405), .ZN(new_n406));
  XOR2_X1   g220(.A(KEYINPUT70), .B(G116), .Z(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G122), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT97), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n239), .A2(G122), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G122), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n242), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT97), .B1(new_n414), .B2(new_n410), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G107), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n408), .A2(KEYINPUT14), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n411), .B1(new_n408), .B2(KEYINPUT14), .ZN(new_n420));
  OAI21_X1  g234(.A(G107), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(G128), .B(G143), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(new_n231), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n418), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT9), .B(G234), .ZN(new_n425));
  NOR3_X1   g239(.A1(new_n425), .A2(new_n341), .A3(G953), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT98), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n412), .A2(new_n415), .A3(G107), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n418), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT13), .B1(new_n227), .B2(G143), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(new_n231), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(new_n422), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n427), .B1(new_n418), .B2(new_n428), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n424), .B(new_n426), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n418), .A2(new_n428), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT98), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n429), .A3(new_n432), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n426), .B1(new_n439), .B2(new_n424), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n278), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G478), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(KEYINPUT15), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  OAI221_X1 g258(.A(new_n278), .B1(KEYINPUT15), .B2(new_n442), .C1(new_n436), .C2(new_n440), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n333), .A2(G952), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(G234), .B2(G237), .ZN(new_n448));
  AOI211_X1 g262(.A(new_n278), .B(new_n333), .C1(G234), .C2(G237), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(G898), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n406), .A2(new_n446), .A3(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G214), .B1(G237), .B2(G902), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(KEYINPUT90), .ZN(new_n454));
  XNOR2_X1  g268(.A(G110), .B(G122), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT91), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n367), .A2(G107), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT3), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT85), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n417), .A2(G104), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT85), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n462), .A3(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  XOR2_X1   g278(.A(KEYINPUT86), .B(G101), .Z(new_n465));
  NAND2_X1  g279(.A1(new_n367), .A2(G107), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n461), .B2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n464), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G101), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n467), .B1(new_n460), .B2(new_n463), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n469), .B(KEYINPUT4), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n470), .B1(new_n464), .B2(new_n468), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT4), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n250), .A2(new_n457), .A3(new_n472), .A4(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT5), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n244), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(G113), .B1(new_n241), .B2(KEYINPUT5), .ZN(new_n479));
  OAI22_X1  g293(.A1(new_n478), .A2(new_n479), .B1(new_n238), .B2(new_n244), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n470), .B1(new_n461), .B2(new_n466), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n469), .A2(new_n482), .ZN(new_n483));
  OR2_X1    g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n476), .A2(new_n484), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n475), .A2(new_n246), .A3(new_n249), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n457), .B1(new_n486), .B2(new_n472), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n456), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n250), .A2(new_n472), .A3(new_n475), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT91), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n490), .A2(new_n476), .A3(new_n484), .A4(new_n455), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT92), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT6), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n488), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  OAI221_X1 g309(.A(new_n456), .B1(new_n492), .B2(new_n493), .C1(new_n485), .C2(new_n487), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n229), .A2(G125), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n201), .A2(G125), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n333), .A2(G224), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n499), .B(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n495), .A2(new_n496), .A3(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n480), .B(new_n483), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n455), .B(KEYINPUT8), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n500), .A2(KEYINPUT7), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n506), .B1(new_n497), .B2(new_n498), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(KEYINPUT94), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n497), .A2(new_n498), .A3(new_n506), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT93), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n505), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(G902), .B1(new_n511), .B2(new_n491), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n502), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(G210), .B1(G237), .B2(G902), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n502), .A2(new_n512), .A3(new_n514), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n454), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(G469), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n483), .A2(new_n229), .ZN(new_n520));
  INV_X1    g334(.A(new_n229), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(new_n469), .A3(new_n482), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n216), .A2(new_n218), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(KEYINPUT12), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT12), .B1(new_n523), .B2(new_n524), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n521), .A2(new_n469), .A3(KEYINPUT10), .A4(new_n482), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT87), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n481), .B1(new_n471), .B2(new_n465), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n532), .A2(KEYINPUT87), .A3(KEYINPUT10), .A4(new_n521), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n202), .B1(new_n473), .B2(new_n474), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT10), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n535), .A2(new_n472), .B1(new_n522), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n524), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n534), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(G110), .B(G140), .ZN(new_n540));
  INV_X1    g354(.A(G227), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(G953), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n540), .B(new_n542), .Z(new_n543));
  NAND2_X1  g357(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n528), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n534), .A2(new_n537), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n524), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n543), .B1(new_n547), .B2(new_n539), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n519), .B(new_n278), .C1(new_n545), .C2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n539), .B1(new_n526), .B2(new_n527), .ZN(new_n550));
  INV_X1    g364(.A(new_n543), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT88), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n539), .A2(new_n553), .A3(new_n543), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n547), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n553), .B1(new_n539), .B2(new_n543), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n552), .B(G469), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n519), .A2(new_n278), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n549), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT89), .ZN(new_n561));
  OAI21_X1  g375(.A(G221), .B1(new_n425), .B2(G902), .ZN(new_n562));
  XOR2_X1   g376(.A(new_n562), .B(KEYINPUT84), .Z(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n560), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n561), .B1(new_n560), .B2(new_n564), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n452), .B(new_n518), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n302), .A2(new_n349), .A3(new_n355), .A4(new_n568), .ZN(new_n569));
  XOR2_X1   g383(.A(new_n569), .B(new_n465), .Z(G3));
  NAND2_X1  g384(.A1(new_n298), .A2(new_n278), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G472), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n565), .A2(new_n566), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(new_n348), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n351), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n451), .ZN(new_n576));
  INV_X1    g390(.A(new_n454), .ZN(new_n577));
  INV_X1    g391(.A(new_n517), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n514), .B1(new_n502), .B2(new_n512), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n576), .B(new_n577), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  OR2_X1    g394(.A1(new_n441), .A2(G478), .ZN(new_n581));
  OR3_X1    g395(.A1(new_n436), .A2(new_n440), .A3(KEYINPUT33), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT33), .B1(new_n436), .B2(new_n440), .ZN(new_n583));
  AOI21_X1  g397(.A(G902), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n406), .B(new_n581), .C1(new_n584), .C2(new_n442), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n575), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(KEYINPUT99), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(KEYINPUT34), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT100), .B(G104), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G6));
  INV_X1    g406(.A(new_n406), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n446), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n580), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT101), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n575), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT35), .B(G107), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G9));
  NOR2_X1   g413(.A1(new_n336), .A2(KEYINPUT36), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(new_n330), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n346), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n602), .B1(new_n340), .B2(new_n344), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT102), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g419(.A(KEYINPUT102), .B(new_n602), .C1(new_n340), .C2(new_n344), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n568), .A2(new_n572), .A3(new_n607), .A4(new_n351), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT37), .B(G110), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G12));
  INV_X1    g424(.A(new_n518), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n573), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n607), .ZN(new_n613));
  INV_X1    g427(.A(G900), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n449), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n448), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n594), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n613), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n302), .A2(new_n355), .A3(new_n612), .A4(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G128), .ZN(G30));
  NAND2_X1  g437(.A1(new_n270), .A2(new_n274), .ZN(new_n624));
  AOI21_X1  g438(.A(G902), .B1(new_n285), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n353), .B1(new_n187), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n617), .B(KEYINPUT39), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n573), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  OR2_X1    g446(.A1(new_n632), .A2(KEYINPUT40), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(KEYINPUT40), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n516), .A2(new_n517), .ZN(new_n635));
  XOR2_X1   g449(.A(new_n635), .B(KEYINPUT38), .Z(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n603), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n406), .A2(new_n446), .ZN(new_n639));
  AND4_X1   g453(.A1(new_n577), .A2(new_n637), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n628), .A2(new_n633), .A3(new_n634), .A4(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G143), .ZN(G45));
  NOR2_X1   g456(.A1(new_n585), .A2(new_n618), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n613), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n302), .A2(new_n355), .A3(new_n612), .A4(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n354), .B1(new_n353), .B2(new_n283), .ZN(new_n649));
  AOI211_X1 g463(.A(KEYINPUT77), .B(new_n282), .C1(new_n352), .C2(new_n299), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n651), .A2(KEYINPUT104), .A3(new_n612), .A4(new_n645), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G146), .ZN(G48));
  OR2_X1    g468(.A1(new_n545), .A2(new_n548), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n278), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(new_n657), .A3(G469), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n655), .B(new_n278), .C1(KEYINPUT105), .C2(new_n519), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n661), .A2(new_n562), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n302), .A2(new_n349), .A3(new_n355), .A4(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n587), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT41), .B(G113), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G15));
  NOR2_X1   g480(.A1(new_n663), .A2(new_n596), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n239), .ZN(G18));
  NAND2_X1  g482(.A1(new_n661), .A2(new_n562), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n611), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n670), .A2(new_n452), .A3(new_n607), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n302), .A2(new_n355), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G119), .ZN(G21));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT106), .B(G472), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n571), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n275), .A2(new_n254), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n294), .B(new_n292), .C1(new_n195), .C2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(G472), .A2(G902), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n676), .A2(new_n349), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n639), .A2(new_n518), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n662), .A2(new_n576), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n674), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n669), .A2(new_n682), .A3(new_n451), .ZN(new_n686));
  AOI22_X1  g500(.A1(new_n571), .A2(new_n675), .B1(new_n678), .B2(new_n679), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n686), .A2(new_n687), .A3(KEYINPUT107), .A4(new_n349), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G122), .ZN(G24));
  AND2_X1   g504(.A1(new_n687), .A2(new_n603), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n643), .A3(new_n670), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G125), .ZN(G27));
  AOI21_X1  g507(.A(new_n348), .B1(new_n353), .B2(new_n283), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n635), .A2(new_n454), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n562), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n549), .A2(new_n559), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n555), .A2(new_n556), .ZN(new_n698));
  OR2_X1    g512(.A1(new_n698), .A2(KEYINPUT108), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(KEYINPUT108), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n699), .A2(new_n552), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n697), .B1(new_n701), .B2(G469), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n644), .A2(new_n696), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n694), .A2(KEYINPUT42), .A3(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT42), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n696), .A2(new_n702), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n302), .A2(new_n349), .A3(new_n355), .A4(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n706), .B1(new_n708), .B2(new_n644), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI211_X1 g525(.A(KEYINPUT109), .B(new_n706), .C1(new_n708), .C2(new_n644), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n705), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n230), .ZN(G33));
  OAI21_X1  g528(.A(KEYINPUT110), .B1(new_n708), .B2(new_n620), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n649), .A2(new_n650), .A3(new_n348), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n716), .A2(new_n717), .A3(new_n619), .A4(new_n707), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G134), .ZN(G36));
  INV_X1    g534(.A(new_n695), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n581), .B1(new_n584), .B2(new_n442), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n406), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(KEYINPUT43), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n724), .A2(new_n603), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n572), .A2(new_n351), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n721), .B1(new_n727), .B2(KEYINPUT44), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n701), .A2(KEYINPUT45), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n552), .B1(new_n555), .B2(new_n556), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n519), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(KEYINPUT46), .A3(new_n559), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n549), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT46), .B1(new_n733), .B2(new_n559), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n562), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n630), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n728), .B(new_n738), .C1(KEYINPUT44), .C2(new_n727), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G137), .ZN(G39));
  XNOR2_X1  g554(.A(new_n737), .B(KEYINPUT47), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n643), .A2(new_n348), .A3(new_n695), .ZN(new_n742));
  OR3_X1    g556(.A1(new_n741), .A2(new_n651), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G140), .ZN(G42));
  NOR2_X1   g558(.A1(G952), .A2(G953), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n622), .A2(new_n692), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n638), .A2(new_n562), .A3(new_n617), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n747), .A2(new_n682), .A3(new_n702), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n628), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n653), .A2(new_n746), .A3(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n653), .A2(KEYINPUT52), .A3(new_n746), .A4(new_n749), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(KEYINPUT114), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n750), .A2(new_n755), .A3(new_n751), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n580), .B1(new_n585), .B2(new_n594), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n574), .A2(new_n572), .A3(new_n351), .A4(new_n758), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n608), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n569), .A2(new_n672), .A3(new_n689), .A4(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n664), .ZN(new_n762));
  INV_X1    g576(.A(new_n667), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n691), .A2(new_n703), .ZN(new_n764));
  OR3_X1    g578(.A1(new_n406), .A2(new_n446), .A3(new_n618), .ZN(new_n765));
  NOR4_X1   g579(.A1(new_n613), .A2(new_n573), .A3(new_n721), .A4(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n302), .A2(new_n766), .A3(new_n355), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT112), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n651), .A2(new_n769), .A3(new_n766), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n764), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n762), .A2(new_n719), .A3(new_n763), .A4(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n713), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n757), .A2(KEYINPUT53), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n622), .A2(new_n692), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(new_n648), .B2(new_n652), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT52), .B1(new_n777), .B2(new_n749), .ZN(new_n778));
  INV_X1    g592(.A(new_n753), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n775), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n752), .A2(KEYINPUT116), .A3(new_n753), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n773), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n774), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n754), .A2(new_n756), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n772), .B2(new_n713), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n719), .A2(new_n771), .ZN(new_n791));
  INV_X1    g605(.A(new_n712), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n651), .A2(new_n349), .A3(new_n643), .A4(new_n707), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT109), .B1(new_n793), .B2(new_n706), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n704), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n761), .A2(new_n664), .A3(new_n667), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n791), .A2(new_n795), .A3(KEYINPUT113), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n788), .B1(new_n790), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT115), .B1(new_n798), .B2(KEYINPUT53), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n797), .A2(new_n790), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n800), .B(new_n783), .C1(new_n801), .C2(new_n788), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n782), .A2(new_n783), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n799), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n787), .B1(new_n804), .B2(KEYINPUT54), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n724), .A2(new_n448), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n806), .A2(new_n349), .A3(new_n687), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n807), .A2(new_n454), .A3(new_n636), .A4(new_n662), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT50), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n696), .A2(new_n660), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n349), .A3(new_n448), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n628), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n813), .A2(new_n593), .A3(new_n722), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n806), .A2(new_n810), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT118), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n809), .B(new_n814), .C1(new_n691), .C2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n661), .A2(new_n563), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n741), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n807), .A2(new_n695), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n818), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n817), .A2(new_n822), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n819), .B(KEYINPUT117), .Z(new_n824));
  NAND2_X1  g638(.A1(new_n741), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n821), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT51), .B1(new_n817), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n812), .A2(new_n585), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n816), .A2(new_n694), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT48), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n447), .B1(new_n807), .B2(new_n670), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n823), .A2(new_n827), .A3(new_n828), .A4(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n745), .B1(new_n805), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n349), .A2(new_n577), .A3(new_n564), .ZN(new_n835));
  XOR2_X1   g649(.A(new_n835), .B(KEYINPUT111), .Z(new_n836));
  XOR2_X1   g650(.A(new_n660), .B(KEYINPUT49), .Z(new_n837));
  NAND3_X1  g651(.A1(new_n836), .A2(new_n723), .A3(new_n837), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n838), .A2(new_n628), .A3(new_n637), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT119), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n841));
  INV_X1    g655(.A(new_n839), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n802), .A2(new_n803), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n797), .A2(new_n790), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n757), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n800), .B1(new_n845), .B2(new_n783), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT54), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n833), .A2(new_n847), .A3(new_n786), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n841), .B(new_n842), .C1(new_n848), .C2(new_n745), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n840), .A2(new_n849), .ZN(G75));
  NOR2_X1   g664(.A1(new_n333), .A2(G952), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n774), .A2(new_n784), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(G902), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT56), .B1(new_n855), .B2(G210), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n495), .A2(new_n496), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(new_n501), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT55), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n852), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(new_n856), .B2(new_n859), .ZN(G51));
  NAND2_X1  g675(.A1(new_n853), .A2(KEYINPUT54), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n786), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n558), .B(KEYINPUT57), .Z(new_n865));
  OAI21_X1  g679(.A(new_n655), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n854), .A2(new_n733), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n851), .B1(new_n866), .B2(new_n867), .ZN(G54));
  NAND3_X1  g682(.A1(new_n855), .A2(KEYINPUT58), .A3(G475), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n402), .A2(new_n397), .ZN(new_n870));
  OR3_X1    g684(.A1(new_n869), .A2(KEYINPUT120), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT120), .B1(new_n869), .B2(new_n870), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n851), .B1(new_n869), .B2(new_n870), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(G60));
  NAND2_X1  g688(.A1(G478), .A2(G902), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT59), .Z(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n582), .B2(new_n583), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n851), .B1(new_n863), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n876), .B1(new_n847), .B2(new_n786), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n582), .A2(new_n583), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g697(.A(KEYINPUT121), .B(new_n878), .C1(new_n879), .C2(new_n880), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(G63));
  NAND2_X1  g699(.A1(G217), .A2(G902), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT60), .Z(new_n887));
  NAND2_X1  g701(.A1(new_n853), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n851), .B1(new_n888), .B2(new_n337), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n853), .A2(new_n601), .A3(new_n887), .ZN(new_n890));
  AOI22_X1  g704(.A1(new_n889), .A2(new_n890), .B1(KEYINPUT122), .B2(KEYINPUT61), .ZN(new_n891));
  NOR2_X1   g705(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n891), .B(new_n892), .ZN(G66));
  NAND2_X1  g707(.A1(G224), .A2(G953), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n450), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n796), .B2(new_n333), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n857), .B1(G898), .B2(new_n333), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n896), .B(new_n897), .ZN(G69));
  XNOR2_X1  g712(.A(new_n777), .B(KEYINPUT124), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n641), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT62), .Z(new_n901));
  AND2_X1   g715(.A1(new_n743), .A2(new_n739), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n594), .A2(new_n585), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n716), .A2(new_n631), .A3(new_n695), .A4(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT123), .Z(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(new_n393), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n908), .A2(G953), .ZN(new_n909));
  OAI21_X1  g723(.A(G953), .B1(new_n541), .B2(new_n614), .ZN(new_n910));
  AOI22_X1  g724(.A1(new_n905), .A2(new_n909), .B1(KEYINPUT126), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n333), .A2(G900), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n738), .A2(new_n683), .A3(new_n694), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n902), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n914), .A2(new_n795), .A3(new_n719), .A4(new_n899), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n912), .B1(new_n915), .B2(new_n333), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n919), .A3(new_n908), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n911), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n910), .A2(KEYINPUT126), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(G72));
  XNOR2_X1  g737(.A(new_n269), .B(KEYINPUT127), .ZN(new_n924));
  OR3_X1    g738(.A1(new_n915), .A2(new_n195), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n195), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n925), .B1(new_n905), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n796), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n924), .B(new_n195), .ZN(new_n929));
  NAND2_X1  g743(.A1(G472), .A2(G902), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT63), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n928), .A2(new_n852), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n931), .B1(new_n271), .B2(new_n285), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(new_n804), .B2(new_n934), .ZN(G57));
endmodule


