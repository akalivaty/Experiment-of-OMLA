

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771;

  XNOR2_X1 U380 ( .A(n385), .B(n546), .ZN(n738) );
  INV_X2 U381 ( .A(G953), .ZN(n759) );
  INV_X1 U382 ( .A(G125), .ZN(n383) );
  XNOR2_X1 U383 ( .A(n568), .B(n421), .ZN(n593) );
  XNOR2_X1 U384 ( .A(n383), .B(G146), .ZN(n528) );
  AND2_X2 U385 ( .A1(n465), .A2(n394), .ZN(n390) );
  OR2_X1 U386 ( .A1(n757), .A2(KEYINPUT2), .ZN(n682) );
  XNOR2_X1 U387 ( .A(n655), .B(KEYINPUT85), .ZN(n757) );
  NAND2_X1 U388 ( .A1(n460), .A2(n458), .ZN(n655) );
  NOR2_X1 U389 ( .A1(n597), .A2(n491), .ZN(n453) );
  AND2_X1 U390 ( .A1(n648), .A2(n365), .ZN(n399) );
  AND2_X1 U391 ( .A1(n450), .A2(n586), .ZN(n475) );
  NOR2_X1 U392 ( .A1(n585), .A2(n593), .ZN(n657) );
  NOR2_X1 U393 ( .A1(n449), .A2(n615), .ZN(n639) );
  OR2_X1 U394 ( .A1(n695), .A2(n700), .ZN(n591) );
  AND2_X1 U395 ( .A1(n609), .A2(n443), .ZN(n576) );
  INV_X1 U396 ( .A(n593), .ZN(n695) );
  XNOR2_X1 U397 ( .A(n474), .B(n552), .ZN(n574) );
  XNOR2_X2 U398 ( .A(n740), .B(n376), .ZN(n391) );
  OR2_X1 U399 ( .A1(n544), .A2(G902), .ZN(n382) );
  NOR2_X1 U400 ( .A1(n666), .A2(n635), .ZN(n636) );
  NOR2_X1 U401 ( .A1(KEYINPUT47), .A2(n686), .ZN(n634) );
  XNOR2_X1 U402 ( .A(n521), .B(n461), .ZN(n581) );
  XNOR2_X1 U403 ( .A(n462), .B(G475), .ZN(n461) );
  NOR2_X1 U404 ( .A1(G902), .A2(n727), .ZN(n521) );
  INV_X1 U405 ( .A(KEYINPUT13), .ZN(n462) );
  NOR2_X1 U406 ( .A1(n655), .A2(n431), .ZN(n430) );
  NAND2_X1 U407 ( .A1(n654), .A2(n653), .ZN(n465) );
  XOR2_X1 U408 ( .A(G140), .B(G131), .Z(n547) );
  XNOR2_X1 U409 ( .A(n530), .B(G110), .ZN(n546) );
  XNOR2_X1 U410 ( .A(G104), .B(KEYINPUT93), .ZN(n530) );
  NOR2_X1 U411 ( .A1(n359), .A2(n368), .ZN(n426) );
  NAND2_X1 U412 ( .A1(n390), .A2(G472), .ZN(n464) );
  XOR2_X1 U413 ( .A(KEYINPUT108), .B(n524), .Z(n686) );
  INV_X1 U414 ( .A(n657), .ZN(n586) );
  XOR2_X1 U415 ( .A(KEYINPUT66), .B(KEYINPUT8), .Z(n507) );
  XNOR2_X1 U416 ( .A(n528), .B(KEYINPUT10), .ZN(n556) );
  NOR2_X1 U417 ( .A1(n769), .A2(n459), .ZN(n458) );
  XNOR2_X1 U418 ( .A(n396), .B(n370), .ZN(n460) );
  INV_X1 U419 ( .A(n767), .ZN(n459) );
  XNOR2_X1 U420 ( .A(n463), .B(n529), .ZN(n387) );
  NAND2_X1 U421 ( .A1(n759), .A2(G224), .ZN(n529) );
  INV_X1 U422 ( .A(n528), .ZN(n463) );
  OR2_X1 U423 ( .A1(n591), .A2(n589), .ZN(n429) );
  OR2_X1 U424 ( .A1(G902), .A2(G237), .ZN(n535) );
  XNOR2_X1 U425 ( .A(n574), .B(KEYINPUT1), .ZN(n609) );
  XNOR2_X1 U426 ( .A(n470), .B(n498), .ZN(n469) );
  XNOR2_X1 U427 ( .A(n500), .B(n471), .ZN(n470) );
  XNOR2_X1 U428 ( .A(n531), .B(n532), .ZN(n385) );
  XOR2_X1 U429 ( .A(KEYINPUT16), .B(KEYINPUT73), .Z(n532) );
  XOR2_X1 U430 ( .A(KEYINPUT78), .B(KEYINPUT98), .Z(n561) );
  XNOR2_X1 U431 ( .A(G110), .B(G140), .ZN(n560) );
  XNOR2_X1 U432 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U433 ( .A(n554), .B(KEYINPUT24), .ZN(n555) );
  INV_X1 U434 ( .A(KEYINPUT23), .ZN(n554) );
  XNOR2_X1 U435 ( .A(n558), .B(n752), .ZN(n454) );
  XOR2_X1 U436 ( .A(G128), .B(G119), .Z(n558) );
  XNOR2_X1 U437 ( .A(n456), .B(n455), .ZN(n517) );
  XNOR2_X1 U438 ( .A(G104), .B(G122), .ZN(n455) );
  XNOR2_X1 U439 ( .A(n457), .B(KEYINPUT103), .ZN(n456) );
  INV_X1 U440 ( .A(KEYINPUT11), .ZN(n457) );
  INV_X1 U441 ( .A(KEYINPUT12), .ZN(n514) );
  NOR2_X1 U442 ( .A1(G237), .A2(G953), .ZN(n499) );
  XNOR2_X1 U443 ( .A(n619), .B(n416), .ZN(n649) );
  INV_X1 U444 ( .A(KEYINPUT39), .ZN(n416) );
  INV_X1 U445 ( .A(n429), .ZN(n425) );
  NAND2_X1 U446 ( .A1(n429), .A2(KEYINPUT32), .ZN(n424) );
  XNOR2_X1 U447 ( .A(n583), .B(n573), .ZN(n578) );
  XNOR2_X1 U448 ( .A(n616), .B(KEYINPUT6), .ZN(n607) );
  XNOR2_X1 U449 ( .A(n567), .B(n363), .ZN(n421) );
  OR2_X2 U450 ( .A1(n583), .A2(n369), .ZN(n392) );
  BUF_X1 U451 ( .A(n609), .Z(n451) );
  INV_X1 U452 ( .A(n684), .ZN(n394) );
  XNOR2_X1 U453 ( .A(n408), .B(n407), .ZN(n725) );
  XNOR2_X1 U454 ( .A(n551), .B(n477), .ZN(n408) );
  XOR2_X1 U455 ( .A(n546), .B(n545), .Z(n477) );
  AND2_X1 U456 ( .A1(n405), .A2(n403), .ZN(n402) );
  INV_X1 U457 ( .A(KEYINPUT109), .ZN(n436) );
  INV_X1 U458 ( .A(n686), .ZN(n445) );
  NAND2_X1 U459 ( .A1(n399), .A2(n397), .ZN(n396) );
  XNOR2_X1 U460 ( .A(n636), .B(n398), .ZN(n397) );
  INV_X1 U461 ( .A(KEYINPUT74), .ZN(n398) );
  NAND2_X1 U462 ( .A1(G234), .A2(G237), .ZN(n536) );
  INV_X1 U463 ( .A(n607), .ZN(n483) );
  XNOR2_X1 U464 ( .A(n576), .B(KEYINPUT111), .ZN(n577) );
  XNOR2_X1 U465 ( .A(n473), .B(n472), .ZN(n471) );
  INV_X1 U466 ( .A(KEYINPUT101), .ZN(n472) );
  XNOR2_X1 U467 ( .A(KEYINPUT5), .B(G137), .ZN(n473) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n491) );
  INV_X1 U469 ( .A(KEYINPUT64), .ZN(n410) );
  XOR2_X1 U470 ( .A(KEYINPUT15), .B(G902), .Z(n600) );
  XOR2_X1 U471 ( .A(G146), .B(G134), .Z(n548) );
  NOR2_X1 U472 ( .A1(n422), .A2(KEYINPUT2), .ZN(n681) );
  AND2_X1 U473 ( .A1(n481), .A2(n484), .ZN(n480) );
  NAND2_X1 U474 ( .A1(n607), .A2(n488), .ZN(n484) );
  OR2_X1 U475 ( .A1(n577), .A2(n482), .ZN(n481) );
  NAND2_X1 U476 ( .A1(n483), .A2(KEYINPUT33), .ZN(n482) );
  XNOR2_X1 U477 ( .A(n512), .B(G478), .ZN(n582) );
  XNOR2_X1 U478 ( .A(n581), .B(n522), .ZN(n523) );
  NOR2_X1 U479 ( .A1(n725), .A2(G902), .ZN(n474) );
  XOR2_X1 U480 ( .A(KEYINPUT105), .B(G134), .Z(n505) );
  XOR2_X1 U481 ( .A(KEYINPUT79), .B(G107), .Z(n545) );
  XNOR2_X1 U482 ( .A(n391), .B(n384), .ZN(n721) );
  XNOR2_X1 U483 ( .A(n386), .B(n738), .ZN(n384) );
  XNOR2_X1 U484 ( .A(n387), .B(n527), .ZN(n386) );
  NOR2_X1 U485 ( .A1(n451), .A2(n418), .ZN(n417) );
  INV_X1 U486 ( .A(n689), .ZN(n418) );
  NAND2_X1 U487 ( .A1(n479), .A2(n480), .ZN(n487) );
  NOR2_X1 U488 ( .A1(n412), .A2(n578), .ZN(n479) );
  INV_X1 U489 ( .A(n485), .ZN(n412) );
  INV_X1 U490 ( .A(KEYINPUT34), .ZN(n486) );
  XNOR2_X1 U491 ( .A(n617), .B(n468), .ZN(n467) );
  XNOR2_X1 U492 ( .A(KEYINPUT30), .B(KEYINPUT115), .ZN(n468) );
  XNOR2_X1 U493 ( .A(n395), .B(KEYINPUT107), .ZN(n659) );
  NOR2_X1 U494 ( .A1(n523), .A2(n582), .ZN(n395) );
  XNOR2_X1 U495 ( .A(n388), .B(n497), .ZN(n740) );
  XNOR2_X1 U496 ( .A(n496), .B(KEYINPUT70), .ZN(n388) );
  XNOR2_X1 U497 ( .A(n557), .B(n454), .ZN(n565) );
  XNOR2_X1 U498 ( .A(n517), .B(n516), .ZN(n518) );
  INV_X1 U499 ( .A(G475), .ZN(n393) );
  NAND2_X1 U500 ( .A1(n415), .A2(n673), .ZN(n622) );
  INV_X1 U501 ( .A(n649), .ZN(n415) );
  NAND2_X1 U502 ( .A1(n361), .A2(n378), .ZN(n770) );
  NAND2_X1 U503 ( .A1(n381), .A2(n380), .ZN(n378) );
  AND2_X1 U504 ( .A1(n425), .A2(n428), .ZN(n380) );
  NAND2_X1 U505 ( .A1(n362), .A2(n379), .ZN(n665) );
  NOR2_X1 U506 ( .A1(n451), .A2(KEYINPUT110), .ZN(n427) );
  NAND2_X1 U507 ( .A1(n414), .A2(n705), .ZN(n413) );
  INV_X1 U508 ( .A(n615), .ZN(n414) );
  NAND2_X1 U509 ( .A1(n438), .A2(n434), .ZN(n432) );
  XNOR2_X1 U510 ( .A(n464), .B(n656), .ZN(n438) );
  XNOR2_X1 U511 ( .A(n723), .B(n441), .ZN(n726) );
  XNOR2_X1 U512 ( .A(n725), .B(n724), .ZN(n441) );
  INV_X1 U513 ( .A(KEYINPUT53), .ZN(n439) );
  NAND2_X1 U514 ( .A1(n402), .A2(n400), .ZN(n440) );
  NAND2_X1 U515 ( .A1(n401), .A2(n685), .ZN(n400) );
  AND2_X1 U516 ( .A1(n451), .A2(KEYINPUT110), .ZN(n359) );
  NOR2_X1 U517 ( .A1(n684), .A2(n685), .ZN(n360) );
  AND2_X1 U518 ( .A1(n377), .A2(n424), .ZN(n361) );
  AND2_X1 U519 ( .A1(n423), .A2(n426), .ZN(n362) );
  XOR2_X1 U520 ( .A(n553), .B(KEYINPUT99), .Z(n363) );
  XOR2_X1 U521 ( .A(n533), .B(KEYINPUT94), .Z(n364) );
  XOR2_X1 U522 ( .A(n630), .B(n629), .Z(n365) );
  NOR2_X1 U523 ( .A1(n684), .A2(n393), .ZN(n366) );
  NAND2_X1 U524 ( .A1(n720), .A2(n759), .ZN(n367) );
  NAND2_X1 U525 ( .A1(n593), .A2(n705), .ZN(n368) );
  OR2_X1 U526 ( .A1(n690), .A2(n601), .ZN(n369) );
  INV_X1 U527 ( .A(KEYINPUT32), .ZN(n428) );
  XOR2_X1 U528 ( .A(KEYINPUT68), .B(KEYINPUT48), .Z(n370) );
  XOR2_X1 U529 ( .A(KEYINPUT86), .B(KEYINPUT35), .Z(n371) );
  XOR2_X1 U530 ( .A(n727), .B(n490), .Z(n372) );
  XOR2_X1 U531 ( .A(n721), .B(n489), .Z(n373) );
  NOR2_X1 U532 ( .A1(G952), .A2(n759), .ZN(n737) );
  INV_X1 U533 ( .A(n737), .ZN(n434) );
  XNOR2_X1 U534 ( .A(KEYINPUT63), .B(KEYINPUT92), .ZN(n374) );
  XNOR2_X1 U535 ( .A(KEYINPUT87), .B(KEYINPUT56), .ZN(n375) );
  INV_X1 U536 ( .A(KEYINPUT2), .ZN(n431) );
  INV_X1 U537 ( .A(KEYINPUT84), .ZN(n685) );
  XNOR2_X1 U538 ( .A(n376), .B(n547), .ZN(n407) );
  XNOR2_X2 U539 ( .A(n755), .B(G101), .ZN(n376) );
  NAND2_X1 U540 ( .A1(n590), .A2(KEYINPUT32), .ZN(n377) );
  NAND2_X1 U541 ( .A1(n665), .A2(n770), .ZN(n596) );
  NAND2_X1 U542 ( .A1(n381), .A2(n427), .ZN(n379) );
  INV_X1 U543 ( .A(n590), .ZN(n381) );
  XNOR2_X2 U544 ( .A(n382), .B(G472), .ZN(n616) );
  XNOR2_X2 U545 ( .A(n478), .B(n503), .ZN(n755) );
  XNOR2_X2 U546 ( .A(n389), .B(KEYINPUT102), .ZN(n660) );
  NOR2_X2 U547 ( .A1(n578), .A2(n413), .ZN(n389) );
  XNOR2_X2 U548 ( .A(n543), .B(KEYINPUT0), .ZN(n583) );
  NAND2_X1 U549 ( .A1(n390), .A2(G210), .ZN(n722) );
  NAND2_X1 U550 ( .A1(n390), .A2(G478), .ZN(n730) );
  NAND2_X1 U551 ( .A1(n390), .A2(G217), .ZN(n734) );
  NAND2_X1 U552 ( .A1(n390), .A2(G469), .ZN(n723) );
  XNOR2_X1 U553 ( .A(n469), .B(n391), .ZN(n544) );
  XNOR2_X2 U554 ( .A(n392), .B(n584), .ZN(n590) );
  AND2_X1 U555 ( .A1(n684), .A2(n685), .ZN(n404) );
  NAND2_X1 U556 ( .A1(n659), .A2(n620), .ZN(n524) );
  INV_X1 U557 ( .A(n406), .ZN(n401) );
  NOR2_X1 U558 ( .A1(n404), .A2(n367), .ZN(n403) );
  NAND2_X1 U559 ( .A1(n406), .A2(n360), .ZN(n405) );
  XNOR2_X2 U560 ( .A(n452), .B(n683), .ZN(n406) );
  NAND2_X1 U561 ( .A1(n409), .A2(n475), .ZN(n587) );
  NAND2_X1 U562 ( .A1(n588), .A2(KEYINPUT44), .ZN(n409) );
  XNOR2_X1 U563 ( .A(n437), .B(n436), .ZN(n450) );
  XNOR2_X1 U564 ( .A(n565), .B(n564), .ZN(n733) );
  NAND2_X1 U565 ( .A1(n596), .A2(KEYINPUT44), .ZN(n411) );
  NAND2_X1 U566 ( .A1(n467), .A2(n614), .ZN(n449) );
  NAND2_X1 U567 ( .A1(n465), .A2(n366), .ZN(n728) );
  NAND2_X1 U568 ( .A1(n419), .A2(n417), .ZN(n610) );
  INV_X1 U569 ( .A(n644), .ZN(n419) );
  NAND2_X1 U570 ( .A1(n420), .A2(n673), .ZN(n644) );
  XNOR2_X1 U571 ( .A(n608), .B(KEYINPUT112), .ZN(n420) );
  AND2_X1 U572 ( .A1(n422), .A2(n430), .ZN(n684) );
  AND2_X1 U573 ( .A1(n422), .A2(n600), .ZN(n651) );
  NAND2_X1 U574 ( .A1(n422), .A2(n759), .ZN(n743) );
  XNOR2_X2 U575 ( .A(n599), .B(KEYINPUT45), .ZN(n422) );
  NAND2_X1 U576 ( .A1(n590), .A2(KEYINPUT110), .ZN(n423) );
  NOR2_X1 U577 ( .A1(n590), .A2(n451), .ZN(n592) );
  AND2_X1 U578 ( .A1(n435), .A2(n434), .ZN(n442) );
  XNOR2_X1 U579 ( .A(n432), .B(n374), .ZN(G57) );
  XNOR2_X1 U580 ( .A(n433), .B(n375), .ZN(G51) );
  NAND2_X1 U581 ( .A1(n444), .A2(n434), .ZN(n433) );
  XNOR2_X1 U582 ( .A(n728), .B(n372), .ZN(n435) );
  XNOR2_X1 U583 ( .A(n595), .B(KEYINPUT71), .ZN(n597) );
  NAND2_X1 U584 ( .A1(n446), .A2(n445), .ZN(n437) );
  XNOR2_X1 U585 ( .A(n440), .B(n439), .ZN(G75) );
  XNOR2_X1 U586 ( .A(n442), .B(KEYINPUT60), .ZN(G60) );
  INV_X2 U587 ( .A(KEYINPUT65), .ZN(n466) );
  XNOR2_X1 U588 ( .A(n487), .B(n486), .ZN(n579) );
  INV_X1 U589 ( .A(n699), .ZN(n443) );
  XNOR2_X1 U590 ( .A(n722), .B(n373), .ZN(n444) );
  NAND2_X1 U591 ( .A1(n448), .A2(n447), .ZN(n446) );
  INV_X1 U592 ( .A(n676), .ZN(n447) );
  INV_X1 U593 ( .A(n660), .ZN(n448) );
  XOR2_X2 U594 ( .A(G122), .B(G107), .Z(n531) );
  NOR2_X1 U595 ( .A1(n706), .A2(n583), .ZN(n572) );
  NAND2_X1 U596 ( .A1(n476), .A2(n682), .ZN(n452) );
  NAND2_X1 U597 ( .A1(n453), .A2(n598), .ZN(n599) );
  INV_X1 U598 ( .A(n768), .ZN(n588) );
  NAND2_X1 U599 ( .A1(n594), .A2(n768), .ZN(n595) );
  XNOR2_X2 U600 ( .A(n580), .B(n371), .ZN(n768) );
  INV_X1 U601 ( .A(n640), .ZN(n618) );
  XNOR2_X2 U602 ( .A(n643), .B(KEYINPUT19), .ZN(n632) );
  NAND2_X2 U603 ( .A1(n640), .A2(n689), .ZN(n643) );
  XNOR2_X2 U604 ( .A(n534), .B(n364), .ZN(n640) );
  XNOR2_X2 U605 ( .A(n466), .B(KEYINPUT4), .ZN(n478) );
  NAND2_X1 U606 ( .A1(n639), .A2(n688), .ZN(n619) );
  NAND2_X1 U607 ( .A1(n575), .A2(n695), .ZN(n615) );
  XNOR2_X1 U608 ( .A(n681), .B(KEYINPUT83), .ZN(n476) );
  NAND2_X1 U609 ( .A1(n577), .A2(n488), .ZN(n485) );
  NAND2_X1 U610 ( .A1(n480), .A2(n485), .ZN(n717) );
  INV_X1 U611 ( .A(KEYINPUT33), .ZN(n488) );
  NAND2_X2 U612 ( .A1(n495), .A2(n494), .ZN(n503) );
  XNOR2_X1 U613 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n489) );
  XNOR2_X1 U614 ( .A(KEYINPUT59), .B(KEYINPUT91), .ZN(n490) );
  INV_X1 U615 ( .A(KEYINPUT46), .ZN(n628) );
  XNOR2_X1 U616 ( .A(n628), .B(KEYINPUT88), .ZN(n629) );
  XNOR2_X1 U617 ( .A(n515), .B(n514), .ZN(n516) );
  INV_X1 U618 ( .A(KEYINPUT82), .ZN(n683) );
  INV_X1 U619 ( .A(KEYINPUT97), .ZN(n573) );
  INV_X1 U620 ( .A(KEYINPUT104), .ZN(n522) );
  XNOR2_X1 U621 ( .A(n563), .B(n562), .ZN(n564) );
  INV_X1 U622 ( .A(G128), .ZN(n492) );
  NAND2_X1 U623 ( .A1(G143), .A2(n492), .ZN(n495) );
  INV_X1 U624 ( .A(G143), .ZN(n493) );
  NAND2_X1 U625 ( .A1(n493), .A2(G128), .ZN(n494) );
  XOR2_X1 U626 ( .A(KEYINPUT3), .B(G119), .Z(n497) );
  XNOR2_X1 U627 ( .A(G116), .B(G113), .ZN(n496) );
  XNOR2_X1 U628 ( .A(G131), .B(n548), .ZN(n498) );
  XNOR2_X1 U629 ( .A(n499), .B(KEYINPUT76), .ZN(n513) );
  AND2_X1 U630 ( .A1(n513), .A2(G210), .ZN(n500) );
  XOR2_X1 U631 ( .A(KEYINPUT62), .B(n544), .Z(n656) );
  XOR2_X1 U632 ( .A(KEYINPUT106), .B(KEYINPUT7), .Z(n502) );
  XNOR2_X1 U633 ( .A(G116), .B(KEYINPUT9), .ZN(n501) );
  XNOR2_X1 U634 ( .A(n502), .B(n501), .ZN(n511) );
  XNOR2_X1 U635 ( .A(n503), .B(n531), .ZN(n504) );
  XNOR2_X1 U636 ( .A(n505), .B(n504), .ZN(n509) );
  NAND2_X1 U637 ( .A1(G234), .A2(n759), .ZN(n506) );
  XNOR2_X1 U638 ( .A(n507), .B(n506), .ZN(n559) );
  NAND2_X1 U639 ( .A1(n559), .A2(G217), .ZN(n508) );
  XOR2_X1 U640 ( .A(n509), .B(n508), .Z(n510) );
  XNOR2_X1 U641 ( .A(n511), .B(n510), .ZN(n729) );
  NOR2_X1 U642 ( .A1(G902), .A2(n729), .ZN(n512) );
  XNOR2_X1 U643 ( .A(n556), .B(n547), .ZN(n751) );
  NAND2_X1 U644 ( .A1(n513), .A2(G214), .ZN(n519) );
  XNOR2_X1 U645 ( .A(G143), .B(G113), .ZN(n515) );
  XNOR2_X1 U646 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U647 ( .A(n751), .B(n520), .ZN(n727) );
  NAND2_X1 U648 ( .A1(n582), .A2(n523), .ZN(n620) );
  INV_X1 U649 ( .A(n600), .ZN(n652) );
  XOR2_X1 U650 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n526) );
  XNOR2_X1 U651 ( .A(KEYINPUT90), .B(KEYINPUT80), .ZN(n525) );
  XNOR2_X1 U652 ( .A(n526), .B(n525), .ZN(n527) );
  NAND2_X1 U653 ( .A1(n652), .A2(n721), .ZN(n534) );
  NAND2_X1 U654 ( .A1(n535), .A2(G210), .ZN(n533) );
  NAND2_X1 U655 ( .A1(G214), .A2(n535), .ZN(n689) );
  XOR2_X1 U656 ( .A(KEYINPUT14), .B(KEYINPUT95), .Z(n537) );
  XNOR2_X1 U657 ( .A(n537), .B(n536), .ZN(n539) );
  NAND2_X1 U658 ( .A1(G952), .A2(n539), .ZN(n538) );
  XNOR2_X1 U659 ( .A(KEYINPUT96), .B(n538), .ZN(n715) );
  OR2_X1 U660 ( .A1(G953), .A2(n715), .ZN(n604) );
  NAND2_X1 U661 ( .A1(G902), .A2(n539), .ZN(n602) );
  INV_X1 U662 ( .A(n602), .ZN(n540) );
  NOR2_X1 U663 ( .A1(G898), .A2(n759), .ZN(n741) );
  NAND2_X1 U664 ( .A1(n540), .A2(n741), .ZN(n541) );
  NAND2_X1 U665 ( .A1(n604), .A2(n541), .ZN(n542) );
  NAND2_X1 U666 ( .A1(n632), .A2(n542), .ZN(n543) );
  XNOR2_X1 U667 ( .A(KEYINPUT69), .B(G469), .ZN(n552) );
  XOR2_X2 U668 ( .A(G137), .B(KEYINPUT67), .Z(n752) );
  XNOR2_X1 U669 ( .A(n548), .B(n752), .ZN(n550) );
  NAND2_X1 U670 ( .A1(G227), .A2(n759), .ZN(n549) );
  XNOR2_X1 U671 ( .A(n550), .B(n549), .ZN(n551) );
  INV_X1 U672 ( .A(n609), .ZN(n700) );
  XNOR2_X1 U673 ( .A(KEYINPUT25), .B(KEYINPUT77), .ZN(n553) );
  NAND2_X1 U674 ( .A1(G221), .A2(n559), .ZN(n563) );
  XNOR2_X1 U675 ( .A(n561), .B(n560), .ZN(n562) );
  NOR2_X1 U676 ( .A1(G902), .A2(n733), .ZN(n568) );
  NAND2_X1 U677 ( .A1(G234), .A2(n652), .ZN(n566) );
  XNOR2_X1 U678 ( .A(KEYINPUT20), .B(n566), .ZN(n569) );
  NAND2_X1 U679 ( .A1(n569), .A2(G217), .ZN(n567) );
  NAND2_X1 U680 ( .A1(n569), .A2(G221), .ZN(n570) );
  XNOR2_X1 U681 ( .A(n570), .B(KEYINPUT21), .ZN(n571) );
  XNOR2_X1 U682 ( .A(KEYINPUT100), .B(n571), .ZN(n601) );
  INV_X1 U683 ( .A(n601), .ZN(n696) );
  NAND2_X1 U684 ( .A1(n695), .A2(n696), .ZN(n699) );
  NAND2_X1 U685 ( .A1(n616), .A2(n576), .ZN(n706) );
  XOR2_X1 U686 ( .A(KEYINPUT31), .B(n572), .Z(n676) );
  INV_X1 U687 ( .A(n616), .ZN(n705) );
  AND2_X1 U688 ( .A1(n574), .A2(n696), .ZN(n575) );
  NOR2_X1 U689 ( .A1(n582), .A2(n581), .ZN(n638) );
  NAND2_X1 U690 ( .A1(n579), .A2(n638), .ZN(n580) );
  NAND2_X1 U691 ( .A1(n582), .A2(n581), .ZN(n690) );
  XNOR2_X1 U692 ( .A(KEYINPUT22), .B(KEYINPUT72), .ZN(n584) );
  NAND2_X1 U693 ( .A1(n592), .A2(n607), .ZN(n585) );
  XNOR2_X1 U694 ( .A(n587), .B(KEYINPUT89), .ZN(n598) );
  XNOR2_X1 U695 ( .A(KEYINPUT81), .B(n607), .ZN(n589) );
  NOR2_X1 U696 ( .A1(n596), .A2(KEYINPUT44), .ZN(n594) );
  XOR2_X1 U697 ( .A(KEYINPUT43), .B(KEYINPUT113), .Z(n611) );
  NOR2_X1 U698 ( .A1(n695), .A2(n601), .ZN(n606) );
  NOR2_X1 U699 ( .A1(G900), .A2(n602), .ZN(n603) );
  NAND2_X1 U700 ( .A1(G953), .A2(n603), .ZN(n605) );
  NAND2_X1 U701 ( .A1(n605), .A2(n604), .ZN(n614) );
  NAND2_X1 U702 ( .A1(n606), .A2(n614), .ZN(n623) );
  NOR2_X1 U703 ( .A1(n623), .A2(n607), .ZN(n608) );
  INV_X1 U704 ( .A(n620), .ZN(n673) );
  XNOR2_X1 U705 ( .A(n611), .B(n610), .ZN(n612) );
  NAND2_X1 U706 ( .A1(n612), .A2(n618), .ZN(n613) );
  XOR2_X1 U707 ( .A(KEYINPUT114), .B(n613), .Z(n769) );
  NAND2_X1 U708 ( .A1(n689), .A2(n616), .ZN(n617) );
  XNOR2_X1 U709 ( .A(n618), .B(KEYINPUT38), .ZN(n688) );
  XOR2_X1 U710 ( .A(KEYINPUT116), .B(KEYINPUT40), .Z(n621) );
  XNOR2_X1 U711 ( .A(n622), .B(n621), .ZN(n766) );
  NOR2_X1 U712 ( .A1(n623), .A2(n705), .ZN(n624) );
  XNOR2_X1 U713 ( .A(KEYINPUT28), .B(n624), .ZN(n625) );
  NAND2_X1 U714 ( .A1(n625), .A2(n574), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n689), .A2(n688), .ZN(n687) );
  NOR2_X1 U716 ( .A1(n687), .A2(n690), .ZN(n626) );
  XNOR2_X1 U717 ( .A(n626), .B(KEYINPUT41), .ZN(n716) );
  NOR2_X1 U718 ( .A1(n631), .A2(n716), .ZN(n627) );
  XNOR2_X1 U719 ( .A(n627), .B(KEYINPUT42), .ZN(n771) );
  NOR2_X1 U720 ( .A1(n766), .A2(n771), .ZN(n630) );
  INV_X1 U721 ( .A(n631), .ZN(n633) );
  NAND2_X1 U722 ( .A1(n633), .A2(n632), .ZN(n666) );
  XNOR2_X1 U723 ( .A(n634), .B(KEYINPUT75), .ZN(n635) );
  OR2_X1 U724 ( .A1(n666), .A2(n686), .ZN(n637) );
  NAND2_X1 U725 ( .A1(n637), .A2(KEYINPUT47), .ZN(n642) );
  AND2_X1 U726 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U727 ( .A1(n641), .A2(n640), .ZN(n670) );
  NAND2_X1 U728 ( .A1(n642), .A2(n670), .ZN(n647) );
  NOR2_X1 U729 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U730 ( .A(KEYINPUT36), .B(n645), .Z(n646) );
  NOR2_X1 U731 ( .A1(n700), .A2(n646), .ZN(n678) );
  NOR2_X1 U732 ( .A1(n647), .A2(n678), .ZN(n648) );
  NOR2_X1 U733 ( .A1(n649), .A2(n659), .ZN(n650) );
  XNOR2_X1 U734 ( .A(n650), .B(KEYINPUT117), .ZN(n767) );
  NAND2_X1 U735 ( .A1(n651), .A2(n757), .ZN(n654) );
  OR2_X1 U736 ( .A1(n652), .A2(n431), .ZN(n653) );
  XOR2_X1 U737 ( .A(n657), .B(G101), .Z(G3) );
  NAND2_X1 U738 ( .A1(n660), .A2(n673), .ZN(n658) );
  XNOR2_X1 U739 ( .A(n658), .B(G104), .ZN(G6) );
  XNOR2_X1 U740 ( .A(KEYINPUT26), .B(KEYINPUT118), .ZN(n664) );
  XOR2_X1 U741 ( .A(G107), .B(KEYINPUT27), .Z(n662) );
  INV_X1 U742 ( .A(n659), .ZN(n675) );
  NAND2_X1 U743 ( .A1(n675), .A2(n660), .ZN(n661) );
  XNOR2_X1 U744 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U745 ( .A(n664), .B(n663), .ZN(G9) );
  XNOR2_X1 U746 ( .A(n665), .B(G110), .ZN(G12) );
  XOR2_X1 U747 ( .A(KEYINPUT29), .B(KEYINPUT119), .Z(n668) );
  INV_X1 U748 ( .A(n666), .ZN(n671) );
  NAND2_X1 U749 ( .A1(n671), .A2(n675), .ZN(n667) );
  XNOR2_X1 U750 ( .A(n668), .B(n667), .ZN(n669) );
  XOR2_X1 U751 ( .A(G128), .B(n669), .Z(G30) );
  XNOR2_X1 U752 ( .A(G143), .B(n670), .ZN(G45) );
  NAND2_X1 U753 ( .A1(n671), .A2(n673), .ZN(n672) );
  XNOR2_X1 U754 ( .A(n672), .B(G146), .ZN(G48) );
  NAND2_X1 U755 ( .A1(n676), .A2(n673), .ZN(n674) );
  XNOR2_X1 U756 ( .A(n674), .B(G113), .ZN(G15) );
  NAND2_X1 U757 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U758 ( .A(n677), .B(G116), .ZN(G18) );
  XNOR2_X1 U759 ( .A(n678), .B(KEYINPUT120), .ZN(n679) );
  XNOR2_X1 U760 ( .A(n679), .B(KEYINPUT37), .ZN(n680) );
  XNOR2_X1 U761 ( .A(G125), .B(n680), .ZN(G27) );
  NOR2_X1 U762 ( .A1(n687), .A2(n686), .ZN(n693) );
  NOR2_X1 U763 ( .A1(n689), .A2(n688), .ZN(n691) );
  NOR2_X1 U764 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U765 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U766 ( .A1(n717), .A2(n694), .ZN(n712) );
  NOR2_X1 U767 ( .A1(n696), .A2(n695), .ZN(n698) );
  XNOR2_X1 U768 ( .A(KEYINPUT121), .B(KEYINPUT49), .ZN(n697) );
  XNOR2_X1 U769 ( .A(n698), .B(n697), .ZN(n703) );
  NAND2_X1 U770 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U771 ( .A(KEYINPUT50), .B(n701), .Z(n702) );
  NOR2_X1 U772 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n707) );
  NAND2_X1 U774 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U775 ( .A(n708), .B(KEYINPUT122), .ZN(n709) );
  XNOR2_X1 U776 ( .A(n709), .B(KEYINPUT51), .ZN(n710) );
  NOR2_X1 U777 ( .A1(n716), .A2(n710), .ZN(n711) );
  NOR2_X1 U778 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U779 ( .A(n713), .B(KEYINPUT52), .ZN(n714) );
  NOR2_X1 U780 ( .A1(n715), .A2(n714), .ZN(n719) );
  NOR2_X1 U781 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U782 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U783 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n724) );
  NOR2_X1 U784 ( .A1(n737), .A2(n726), .ZN(G54) );
  XOR2_X1 U785 ( .A(n729), .B(KEYINPUT123), .Z(n731) );
  XNOR2_X1 U786 ( .A(n731), .B(n730), .ZN(n732) );
  NOR2_X1 U787 ( .A1(n737), .A2(n732), .ZN(G63) );
  XNOR2_X1 U788 ( .A(n733), .B(KEYINPUT124), .ZN(n735) );
  XNOR2_X1 U789 ( .A(n735), .B(n734), .ZN(n736) );
  NOR2_X1 U790 ( .A1(n737), .A2(n736), .ZN(G66) );
  XOR2_X1 U791 ( .A(G101), .B(n738), .Z(n739) );
  XNOR2_X1 U792 ( .A(n740), .B(n739), .ZN(n742) );
  NOR2_X1 U793 ( .A1(n742), .A2(n741), .ZN(n750) );
  XNOR2_X1 U794 ( .A(n743), .B(KEYINPUT126), .ZN(n748) );
  XOR2_X1 U795 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n745) );
  NAND2_X1 U796 ( .A1(G224), .A2(G953), .ZN(n744) );
  XNOR2_X1 U797 ( .A(n745), .B(n744), .ZN(n746) );
  NAND2_X1 U798 ( .A1(n746), .A2(G898), .ZN(n747) );
  NAND2_X1 U799 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U800 ( .A(n750), .B(n749), .ZN(G69) );
  XOR2_X1 U801 ( .A(KEYINPUT127), .B(n751), .Z(n754) );
  XNOR2_X1 U802 ( .A(G134), .B(n752), .ZN(n753) );
  XNOR2_X1 U803 ( .A(n754), .B(n753), .ZN(n756) );
  XNOR2_X1 U804 ( .A(n755), .B(n756), .ZN(n761) );
  INV_X1 U805 ( .A(n761), .ZN(n758) );
  XNOR2_X1 U806 ( .A(n758), .B(n757), .ZN(n760) );
  NAND2_X1 U807 ( .A1(n760), .A2(n759), .ZN(n765) );
  XNOR2_X1 U808 ( .A(G227), .B(n761), .ZN(n762) );
  NAND2_X1 U809 ( .A1(n762), .A2(G900), .ZN(n763) );
  NAND2_X1 U810 ( .A1(n763), .A2(G953), .ZN(n764) );
  NAND2_X1 U811 ( .A1(n765), .A2(n764), .ZN(G72) );
  XOR2_X1 U812 ( .A(G131), .B(n766), .Z(G33) );
  XNOR2_X1 U813 ( .A(G134), .B(n767), .ZN(G36) );
  XNOR2_X1 U814 ( .A(n768), .B(G122), .ZN(G24) );
  XOR2_X1 U815 ( .A(G140), .B(n769), .Z(G42) );
  XNOR2_X1 U816 ( .A(n770), .B(G119), .ZN(G21) );
  XOR2_X1 U817 ( .A(G137), .B(n771), .Z(G39) );
endmodule

