//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0002(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0003(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n204));
  NAND2_X1  g0004(.A1(G107), .A2(G264), .ZN(new_n205));
  NAND2_X1  g0005(.A1(G68), .A2(G238), .ZN(new_n206));
  NAND3_X1  g0006(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  AOI21_X1  g0007(.A(new_n207), .B1(G50), .B2(G226), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT67), .ZN(new_n210));
  XNOR2_X1  g0010(.A(KEYINPUT65), .B(G77), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  XOR2_X1   g0012(.A(KEYINPUT66), .B(G244), .Z(new_n213));
  OAI211_X1 g0013(.A(new_n208), .B(new_n210), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G20), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n215), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT0), .Z(new_n220));
  NOR2_X1   g0020(.A1(G58), .A2(G68), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NOR3_X1   g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NOR3_X1   g0026(.A1(new_n217), .A2(new_n220), .A3(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G250), .B(G257), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G264), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n230), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G68), .B(G77), .Z(new_n236));
  XOR2_X1   g0036(.A(G50), .B(G58), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G351));
  XNOR2_X1  g0042(.A(KEYINPUT3), .B(G33), .ZN(new_n243));
  INV_X1    g0043(.A(G1698), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G222), .ZN(new_n245));
  NAND2_X1  g0045(.A1(G223), .A2(G1698), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n243), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G41), .ZN(new_n249));
  OAI211_X1 g0049(.A(G1), .B(G13), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  OAI211_X1 g0051(.A(new_n247), .B(new_n251), .C1(new_n211), .C2(new_n243), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  OAI211_X1 g0053(.A(new_n253), .B(G274), .C1(G41), .C2(G45), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G226), .ZN(new_n258));
  AND3_X1   g0058(.A1(new_n252), .A2(new_n254), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G179), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n225), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n263), .B1(new_n253), .B2(G20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G50), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n253), .A2(G13), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G20), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G50), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NOR3_X1   g0070(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n224), .A2(new_n248), .ZN(new_n272));
  INV_X1    g0072(.A(G150), .ZN(new_n273));
  OAI22_X1  g0073(.A1(new_n271), .A2(new_n224), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(KEYINPUT68), .B1(new_n248), .B2(G20), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT68), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(new_n224), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n274), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n263), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n265), .B(new_n270), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n252), .A2(new_n258), .A3(new_n254), .ZN(new_n284));
  INV_X1    g0084(.A(G169), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n261), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n254), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n243), .A2(G232), .A3(new_n244), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT69), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT3), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G107), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n243), .A2(G238), .A3(G1698), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n243), .A2(KEYINPUT69), .A3(G232), .A4(new_n244), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n292), .A2(new_n297), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n289), .B1(new_n300), .B2(new_n251), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n256), .A2(new_n213), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(new_n260), .A3(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n268), .A2(new_n211), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT70), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n212), .A2(new_n224), .B1(new_n279), .B2(new_n272), .ZN(new_n307));
  XNOR2_X1  g0107(.A(KEYINPUT15), .B(G87), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n275), .B2(new_n277), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n263), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n264), .A2(G77), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n306), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI211_X1 g0112(.A(new_n302), .B(new_n289), .C1(new_n300), .C2(new_n251), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n304), .B(new_n312), .C1(new_n313), .C2(G169), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n280), .A2(new_n278), .ZN(new_n316));
  INV_X1    g0116(.A(G50), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n221), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(G20), .A2(G33), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n318), .A2(G20), .B1(G150), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n282), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n282), .B1(G1), .B2(new_n224), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(new_n317), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n321), .A2(new_n323), .A3(new_n269), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n324), .A2(KEYINPUT9), .B1(new_n259), .B2(G190), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n284), .A2(G200), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT9), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n283), .A2(KEYINPUT72), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT72), .B1(new_n283), .B2(new_n327), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n325), .B(new_n326), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT10), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n283), .A2(new_n327), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT72), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n328), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT10), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n336), .A2(new_n337), .A3(new_n326), .A4(new_n325), .ZN(new_n338));
  AOI211_X1 g0138(.A(new_n288), .B(new_n315), .C1(new_n332), .C2(new_n338), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n306), .A2(new_n310), .A3(new_n311), .ZN(new_n340));
  INV_X1    g0140(.A(G200), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n313), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT71), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n313), .A2(G190), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT71), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n340), .B(new_n345), .C1(new_n313), .C2(new_n341), .ZN(new_n346));
  AND3_X1   g0146(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  OR2_X1    g0147(.A1(G223), .A2(G1698), .ZN(new_n348));
  INV_X1    g0148(.A(G226), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G1698), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n293), .A2(new_n348), .A3(new_n295), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G33), .A2(G87), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n251), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n257), .A2(G232), .ZN(new_n355));
  INV_X1    g0155(.A(G190), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .A4(new_n254), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT79), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n354), .A2(new_n355), .A3(new_n254), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n341), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n289), .B1(new_n353), .B2(new_n251), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT79), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n361), .A2(new_n362), .A3(new_n356), .A4(new_n355), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n358), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G58), .ZN(new_n365));
  INV_X1    g0165(.A(G68), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(G20), .B1(new_n367), .B2(new_n221), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n319), .A2(G159), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT7), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n243), .B2(G20), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n296), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n370), .B1(new_n374), .B2(G68), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n282), .B1(new_n375), .B2(KEYINPUT16), .ZN(new_n376));
  XOR2_X1   g0176(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n248), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n295), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT77), .B1(new_n248), .B2(KEYINPUT3), .ZN(new_n381));
  OAI211_X1 g0181(.A(KEYINPUT7), .B(new_n224), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n366), .B1(new_n382), .B2(new_n372), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n378), .B1(new_n383), .B2(new_n370), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n376), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n280), .A2(new_n268), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(new_n280), .B2(new_n264), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n364), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT17), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n387), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(new_n376), .B2(new_n384), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n359), .A2(new_n260), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n285), .B1(new_n361), .B2(new_n355), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g0195(.A(KEYINPUT78), .B(KEYINPUT18), .C1(new_n392), .C2(new_n395), .ZN(new_n396));
  NOR3_X1   g0196(.A1(new_n243), .A2(new_n371), .A3(G20), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT7), .B1(new_n296), .B2(new_n224), .ZN(new_n398));
  OAI21_X1  g0198(.A(G68), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n370), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT16), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n263), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n382), .A2(new_n372), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G68), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n377), .B1(new_n405), .B2(new_n400), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n387), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  OR2_X1    g0207(.A1(new_n393), .A2(new_n394), .ZN(new_n408));
  XOR2_X1   g0208(.A(KEYINPUT78), .B(KEYINPUT18), .Z(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n392), .A2(KEYINPUT17), .A3(new_n364), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n390), .A2(new_n396), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n347), .A2(new_n412), .ZN(new_n413));
  AND3_X1   g0213(.A1(new_n250), .A2(G238), .A3(new_n255), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n293), .A2(new_n295), .A3(G232), .A4(G1698), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n293), .A2(new_n295), .A3(G226), .A4(new_n244), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G97), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n414), .B1(new_n418), .B2(new_n251), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT74), .B(KEYINPUT13), .ZN(new_n420));
  XOR2_X1   g0220(.A(new_n254), .B(KEYINPUT73), .Z(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n419), .A2(new_n421), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT13), .ZN(new_n424));
  OAI211_X1 g0224(.A(G190), .B(new_n422), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n418), .A2(new_n251), .ZN(new_n426));
  INV_X1    g0226(.A(new_n414), .ZN(new_n427));
  AND4_X1   g0227(.A1(new_n420), .A2(new_n426), .A3(new_n427), .A4(new_n421), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n420), .B1(new_n419), .B2(new_n421), .ZN(new_n429));
  OAI21_X1  g0229(.A(G200), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n224), .A2(G68), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n267), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n432), .B(KEYINPUT12), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n366), .B2(new_n322), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n431), .B1(new_n278), .B2(G77), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n319), .A2(G50), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT11), .B1(new_n438), .B2(new_n282), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT11), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n437), .A2(new_n440), .A3(new_n263), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n434), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n425), .A2(new_n430), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(G169), .B1(new_n428), .B2(new_n429), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT14), .ZN(new_n445));
  OAI211_X1 g0245(.A(G179), .B(new_n422), .C1(new_n423), .C2(new_n424), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT14), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n447), .B(G169), .C1(new_n428), .C2(new_n429), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n445), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n442), .ZN(new_n450));
  AOI211_X1 g0250(.A(KEYINPUT75), .B(new_n443), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT75), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n449), .A2(new_n450), .ZN(new_n453));
  INV_X1    g0253(.A(new_n443), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n339), .B(new_n413), .C1(new_n451), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT80), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n453), .A2(new_n454), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT75), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n453), .A2(new_n452), .A3(new_n454), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT80), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n461), .A2(new_n462), .A3(new_n413), .A4(new_n339), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n224), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT86), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OR3_X1    g0268(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n465), .A2(KEYINPUT86), .A3(new_n224), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n243), .A2(new_n224), .A3(G68), .ZN(new_n472));
  INV_X1    g0272(.A(G97), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n473), .B1(new_n275), .B2(new_n277), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n471), .B(new_n472), .C1(KEYINPUT19), .C2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n266), .A2(new_n224), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n475), .A2(new_n263), .B1(new_n308), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n268), .B(new_n282), .C1(G1), .C2(new_n248), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G87), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n253), .A2(G45), .ZN(new_n481));
  OR2_X1    g0281(.A1(new_n481), .A2(G274), .ZN(new_n482));
  INV_X1    g0282(.A(G250), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n250), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n293), .A2(new_n295), .A3(G238), .A4(new_n244), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT85), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT85), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n243), .A2(new_n489), .A3(G238), .A4(new_n244), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n243), .A2(G244), .A3(G1698), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G33), .A2(G116), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n488), .A2(new_n490), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n486), .B1(new_n493), .B2(new_n251), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n477), .B(new_n480), .C1(new_n341), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(G190), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n472), .B1(new_n474), .B2(KEYINPUT19), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n263), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OR2_X1    g0300(.A1(new_n478), .A2(new_n308), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n476), .A2(new_n308), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n493), .A2(new_n251), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(new_n260), .A3(new_n485), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n494), .A2(G169), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n495), .A2(new_n497), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT82), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(new_n481), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G41), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n515), .A2(KEYINPUT82), .A3(new_n253), .A4(G45), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n512), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n517), .A2(G270), .A3(new_n250), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n512), .A2(new_n516), .A3(G274), .A4(new_n513), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(new_n251), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT87), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n244), .A2(G257), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G264), .A2(G1698), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n243), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n524), .B(new_n251), .C1(G303), .C2(new_n243), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n517), .A2(G270), .A3(new_n250), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT87), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n526), .B(new_n527), .C1(new_n251), .C2(new_n519), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n521), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G283), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n530), .B(new_n224), .C1(G33), .C2(new_n473), .ZN(new_n531));
  INV_X1    g0331(.A(G116), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G20), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n531), .A2(KEYINPUT20), .A3(new_n263), .A4(new_n533), .ZN(new_n534));
  OR2_X1    g0334(.A1(new_n534), .A2(KEYINPUT88), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(KEYINPUT88), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n531), .A2(new_n263), .A3(new_n533), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n535), .B(new_n536), .C1(KEYINPUT20), .C2(new_n537), .ZN(new_n538));
  OR2_X1    g0338(.A1(new_n266), .A2(new_n533), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n479), .A2(G116), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n529), .A2(G169), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT21), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n529), .A2(KEYINPUT21), .A3(G169), .A4(new_n541), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n521), .A2(new_n528), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n546), .A2(G179), .A3(new_n541), .A4(new_n525), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT89), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n529), .A2(G200), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n541), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n529), .B2(new_n356), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n549), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n546), .A2(G190), .A3(new_n525), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n555), .A2(KEYINPUT89), .A3(new_n552), .A4(new_n550), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n548), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT23), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n224), .B2(G107), .ZN(new_n559));
  INV_X1    g0359(.A(G107), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(KEYINPUT23), .A3(G20), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n224), .A2(G33), .A3(G116), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n293), .A2(new_n295), .A3(new_n224), .A4(G87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(KEYINPUT90), .A2(KEYINPUT22), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n562), .B(new_n563), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  OR2_X1    g0367(.A1(KEYINPUT90), .A2(KEYINPUT22), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n564), .A2(new_n568), .A3(new_n565), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(KEYINPUT24), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT24), .ZN(new_n571));
  INV_X1    g0371(.A(new_n569), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n571), .B1(new_n572), .B2(new_n566), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n570), .A2(new_n263), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n479), .A2(G107), .ZN(new_n575));
  NOR3_X1   g0375(.A1(new_n266), .A2(new_n224), .A3(G107), .ZN(new_n576));
  XNOR2_X1  g0376(.A(new_n576), .B(KEYINPUT25), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n517), .A2(G264), .A3(new_n250), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n293), .A2(new_n295), .A3(G250), .A4(new_n244), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT91), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n243), .A2(KEYINPUT91), .A3(G250), .A4(new_n244), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g0385(.A(KEYINPUT92), .B(G294), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G257), .A2(G1698), .ZN(new_n588));
  OAI22_X1  g0388(.A1(new_n587), .A2(new_n248), .B1(new_n296), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n251), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(KEYINPUT93), .B1(new_n519), .B2(new_n251), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n580), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(KEYINPUT93), .B(new_n251), .C1(new_n585), .C2(new_n589), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n592), .A2(new_n356), .A3(new_n593), .ZN(new_n594));
  OR2_X1    g0394(.A1(new_n519), .A2(new_n251), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n517), .A2(G264), .A3(new_n250), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n590), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n597), .A2(new_n341), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n579), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n285), .B1(new_n592), .B2(new_n593), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n597), .A2(new_n260), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n578), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n243), .A2(KEYINPUT4), .A3(G244), .A4(new_n244), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n293), .A2(new_n295), .A3(G244), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT4), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n604), .A2(new_n607), .A3(new_n530), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n243), .A2(G250), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n244), .B1(new_n609), .B2(KEYINPUT4), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n251), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n517), .A2(G257), .A3(new_n250), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n611), .A2(new_n260), .A3(new_n595), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT83), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n611), .A2(new_n595), .A3(new_n612), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n285), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n517), .A2(G257), .A3(new_n250), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n617), .A2(new_n520), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT83), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n618), .A2(new_n619), .A3(new_n260), .A4(new_n611), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n560), .B1(new_n382), .B2(new_n372), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT6), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n622), .A2(new_n473), .A3(G107), .ZN(new_n623));
  XNOR2_X1  g0423(.A(G97), .B(G107), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n623), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(G77), .ZN(new_n626));
  OAI22_X1  g0426(.A1(new_n625), .A2(new_n224), .B1(new_n626), .B2(new_n272), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n263), .B1(new_n621), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n268), .A2(G97), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n479), .B2(G97), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n614), .A2(new_n616), .A3(new_n620), .A4(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT81), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n628), .A2(KEYINPUT81), .A3(new_n630), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n615), .A2(new_n341), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n618), .A2(new_n356), .A3(new_n611), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n635), .A2(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT84), .B1(new_n633), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  INV_X1    g0441(.A(new_n636), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT81), .B1(new_n628), .B2(new_n630), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT84), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n645), .A3(new_n632), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n603), .B1(new_n640), .B2(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n464), .A2(new_n509), .A3(new_n557), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n648), .B(KEYINPUT94), .ZN(G372));
  NAND2_X1  g0449(.A1(new_n332), .A2(new_n338), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n407), .A2(new_n408), .A3(KEYINPUT96), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT96), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n392), .B2(new_n395), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n651), .A2(new_n653), .A3(KEYINPUT18), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT18), .B1(new_n651), .B2(new_n653), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n390), .A2(new_n411), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n454), .A2(new_n315), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n453), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n650), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n662), .A2(new_n287), .ZN(new_n663));
  INV_X1    g0463(.A(new_n464), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n614), .A2(new_n616), .A3(new_n620), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n642), .A2(new_n643), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  INV_X1    g0467(.A(new_n494), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(G200), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n669), .A2(new_n496), .A3(new_n480), .A4(new_n477), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n665), .A2(new_n666), .A3(new_n667), .A4(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT26), .B1(new_n508), .B2(new_n632), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n506), .A2(new_n507), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n671), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT95), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n671), .A2(new_n672), .A3(KEYINPUT95), .A4(new_n674), .ZN(new_n678));
  AND4_X1   g0478(.A1(new_n544), .A2(new_n602), .A3(new_n545), .A4(new_n547), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n599), .A2(new_n644), .A3(new_n632), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n677), .A2(new_n678), .B1(new_n681), .B2(new_n509), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n663), .B1(new_n664), .B2(new_n682), .ZN(G369));
  OR3_X1    g0483(.A1(new_n266), .A2(KEYINPUT27), .A3(G20), .ZN(new_n684));
  OAI21_X1  g0484(.A(KEYINPUT27), .B1(new_n266), .B2(G20), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(G213), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(G343), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n552), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n548), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n554), .A2(new_n556), .ZN(new_n692));
  INV_X1    g0492(.A(new_n548), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n691), .B1(new_n694), .B2(new_n690), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G330), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n599), .B(new_n602), .C1(new_n579), .C2(new_n689), .ZN(new_n698));
  INV_X1    g0498(.A(new_n602), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n688), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT97), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n698), .A2(new_n700), .A3(KEYINPUT97), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n697), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n699), .A2(new_n689), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n693), .A2(new_n688), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n708), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n706), .A2(new_n710), .ZN(G399));
  INV_X1    g0511(.A(new_n218), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G41), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n469), .A2(G116), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(G1), .A3(new_n715), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n716), .A2(KEYINPUT98), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(KEYINPUT98), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n717), .B(new_n718), .C1(new_n223), .C2(new_n714), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n682), .B2(new_n688), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n509), .A2(new_n667), .A3(new_n633), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n665), .A2(new_n670), .A3(new_n666), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n673), .B1(new_n724), .B2(KEYINPUT26), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n633), .A2(new_n639), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n726), .B(new_n599), .C1(new_n548), .C2(new_n699), .ZN(new_n727));
  INV_X1    g0527(.A(new_n670), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n723), .B(new_n725), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(KEYINPUT29), .A3(new_n689), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n722), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n647), .A2(new_n557), .A3(new_n509), .A4(new_n689), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n521), .A2(G179), .A3(new_n525), .A4(new_n528), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n590), .A2(new_n596), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT100), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(KEYINPUT100), .A2(KEYINPUT30), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n618), .A2(new_n494), .A3(new_n611), .A4(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n735), .A2(new_n738), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n738), .B1(new_n735), .B2(new_n742), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n494), .A2(KEYINPUT99), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n494), .A2(KEYINPUT99), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n529), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n615), .A2(new_n597), .A3(new_n260), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI211_X1 g0550(.A(KEYINPUT31), .B(new_n688), .C1(new_n745), .C2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT31), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n743), .A2(new_n744), .A3(new_n750), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n752), .B1(new_n753), .B2(new_n689), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n732), .A2(new_n751), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G330), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n731), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n720), .B1(new_n758), .B2(G1), .ZN(G364));
  INV_X1    g0559(.A(G13), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G20), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n253), .B1(new_n761), .B2(G45), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n713), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n697), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(G330), .B2(new_n695), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G13), .A2(G33), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n224), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT101), .Z(new_n769));
  AOI21_X1  g0569(.A(new_n225), .B1(G20), .B2(new_n285), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n238), .A2(G45), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n712), .A2(new_n243), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G45), .ZN(new_n776));
  INV_X1    g0576(.A(new_n223), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n773), .A2(new_n778), .B1(new_n532), .B2(new_n712), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n243), .A2(G355), .A3(new_n218), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n772), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n341), .A2(G179), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n224), .A2(G190), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G283), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n296), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n224), .A2(new_n356), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n260), .A2(G200), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT102), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n789), .B1(new_n787), .B2(new_n788), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n260), .A2(new_n341), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n787), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT104), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G322), .A2(new_n793), .B1(new_n796), .B2(G326), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G179), .A2(G200), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n224), .B1(new_n798), .B2(G190), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n794), .A2(new_n783), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT33), .B(G317), .Z(new_n801));
  OAI221_X1 g0601(.A(new_n797), .B1(new_n587), .B2(new_n799), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n783), .A2(new_n798), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n786), .B(new_n802), .C1(G329), .C2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G303), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n787), .A2(new_n782), .ZN(new_n807));
  INV_X1    g0607(.A(G311), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n783), .A2(new_n788), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n805), .B1(new_n806), .B2(new_n807), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n795), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n793), .A2(G58), .B1(G50), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n212), .B2(new_n809), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT103), .Z(new_n814));
  INV_X1    g0614(.A(new_n800), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n814), .B1(G68), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n799), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G97), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n804), .A2(G159), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT32), .ZN(new_n820));
  INV_X1    g0620(.A(new_n784), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n820), .B1(G107), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n807), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(G87), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n816), .A2(new_n818), .A3(new_n822), .A4(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n810), .B1(new_n825), .B2(new_n296), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n781), .B1(new_n826), .B2(new_n770), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n827), .B(new_n764), .C1(new_n695), .C2(new_n769), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n766), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(G396));
  NAND3_X1  g0630(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n312), .A2(new_n688), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n315), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n314), .A2(new_n688), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n677), .A2(new_n678), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n681), .A2(new_n509), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n838), .B1(new_n841), .B2(new_n689), .ZN(new_n842));
  NOR3_X1   g0642(.A1(new_n682), .A2(new_n688), .A3(new_n837), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(new_n756), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n713), .B2(new_n763), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n807), .A2(new_n317), .B1(new_n784), .B2(new_n366), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT108), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G137), .A2(new_n811), .B1(new_n815), .B2(G150), .ZN(new_n849));
  INV_X1    g0649(.A(G159), .ZN(new_n850));
  INV_X1    g0650(.A(new_n793), .ZN(new_n851));
  XOR2_X1   g0651(.A(KEYINPUT107), .B(G143), .Z(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n849), .B1(new_n850), .B2(new_n809), .C1(new_n851), .C2(new_n853), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT34), .ZN(new_n855));
  INV_X1    g0655(.A(G132), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n855), .B(new_n243), .C1(new_n856), .C2(new_n803), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n848), .B(new_n857), .C1(G58), .C2(new_n817), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n807), .A2(new_n560), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n793), .A2(G294), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n296), .B1(new_n795), .B2(new_n806), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n818), .B1(new_n808), .B2(new_n803), .ZN(new_n862));
  NOR3_X1   g0662(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n821), .A2(G87), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n863), .B(new_n864), .C1(new_n532), .C2(new_n809), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n859), .B(new_n865), .C1(G283), .C2(new_n815), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n770), .B1(new_n858), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n770), .A2(new_n767), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT105), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n764), .B1(new_n869), .B2(G77), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT106), .ZN(new_n871));
  INV_X1    g0671(.A(new_n767), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n867), .B(new_n871), .C1(new_n872), .C2(new_n838), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n846), .A2(new_n873), .ZN(G384));
  NAND3_X1  g0674(.A1(new_n841), .A2(new_n689), .A3(new_n838), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n836), .ZN(new_n876));
  INV_X1    g0676(.A(new_n686), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n378), .B1(new_n401), .B2(KEYINPUT109), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT109), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n375), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n376), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n387), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n412), .A2(new_n877), .A3(new_n882), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n881), .A2(new_n387), .B1(new_n395), .B2(new_n686), .ZN(new_n884));
  INV_X1    g0684(.A(new_n388), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT37), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n407), .A2(new_n408), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n407), .A2(new_n877), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT37), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n887), .A2(new_n888), .A3(new_n889), .A4(new_n388), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n883), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n883), .A2(new_n891), .A3(KEYINPUT38), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n450), .A2(new_n688), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n453), .A2(new_n454), .A3(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n450), .B(new_n688), .C1(new_n449), .C2(new_n443), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n876), .A2(new_n896), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n658), .A2(new_n686), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n453), .A2(new_n688), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n894), .A2(KEYINPUT39), .A3(new_n895), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n883), .A2(KEYINPUT38), .A3(new_n891), .ZN(new_n905));
  INV_X1    g0705(.A(new_n659), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n651), .A2(new_n653), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT18), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n906), .A2(new_n909), .A3(new_n654), .ZN(new_n910));
  INV_X1    g0710(.A(new_n888), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n888), .A2(new_n388), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT37), .B1(new_n907), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n890), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n905), .B1(new_n916), .B2(new_n893), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n903), .B(new_n904), .C1(new_n917), .C2(KEYINPUT39), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n901), .A2(new_n902), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n464), .A2(new_n722), .A3(new_n730), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n663), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n919), .B(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT40), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n888), .B1(new_n657), .B2(new_n906), .ZN(new_n924));
  INV_X1    g0724(.A(new_n915), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n893), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n923), .B1(new_n926), .B2(new_n895), .ZN(new_n927));
  INV_X1    g0727(.A(new_n900), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n837), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n755), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n755), .A2(new_n896), .A3(new_n929), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n927), .A2(new_n930), .B1(new_n931), .B2(new_n923), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n464), .A2(new_n755), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n932), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(G330), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n922), .B(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n253), .B2(new_n761), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT35), .ZN(new_n938));
  AOI211_X1 g0738(.A(new_n224), .B(new_n225), .C1(new_n625), .C2(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n939), .B(G116), .C1(new_n938), .C2(new_n625), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT36), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n223), .A2(new_n367), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n942), .A2(new_n212), .B1(G50), .B2(new_n366), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(G1), .A3(new_n760), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n937), .A2(new_n941), .A3(new_n944), .ZN(G367));
  NAND2_X1  g0745(.A1(new_n705), .A2(new_n709), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n666), .A2(new_n688), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n726), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n665), .A2(new_n666), .A3(new_n688), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT42), .B1(new_n946), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n708), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n633), .A2(new_n689), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT42), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n705), .A2(new_n955), .A3(new_n709), .A4(new_n950), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n952), .A2(new_n953), .A3(new_n954), .A4(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n689), .B1(new_n477), .B2(new_n480), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n673), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n508), .B2(new_n958), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n957), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n706), .A2(new_n951), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n957), .B(new_n961), .C1(new_n706), .C2(new_n951), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n713), .B(KEYINPUT41), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n706), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n710), .A2(new_n950), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT45), .ZN(new_n973));
  OR3_X1    g0773(.A1(new_n710), .A2(KEYINPUT44), .A3(new_n950), .ZN(new_n974));
  OAI21_X1  g0774(.A(KEYINPUT44), .B1(new_n710), .B2(new_n950), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n971), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT45), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n972), .B(new_n978), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n979), .A2(new_n706), .A3(new_n975), .A4(new_n974), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n705), .A2(new_n709), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n946), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT110), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n696), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n696), .A2(new_n983), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n982), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n981), .A2(new_n984), .A3(new_n946), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n989), .A2(new_n757), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n977), .A2(new_n980), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n970), .B1(new_n991), .B2(new_n758), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n968), .B1(new_n992), .B2(new_n763), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n823), .A2(KEYINPUT46), .A3(G116), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT46), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n807), .B2(new_n532), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n994), .B(new_n996), .C1(new_n587), .C2(new_n800), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(KEYINPUT111), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n785), .B2(new_n809), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n997), .A2(KEYINPUT111), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n796), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n296), .B1(new_n1001), .B2(new_n808), .ZN(new_n1002));
  INV_X1    g0802(.A(G317), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n784), .A2(new_n473), .B1(new_n803), .B2(new_n1003), .ZN(new_n1004));
  NOR4_X1   g0804(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n560), .B2(new_n799), .C1(new_n806), .C2(new_n851), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n793), .A2(G150), .B1(G68), .B2(new_n817), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT112), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n809), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(G50), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n823), .A2(G58), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1009), .A2(new_n243), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n796), .B2(new_n852), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n1007), .A2(new_n1008), .B1(G159), .B2(new_n815), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1014), .B(new_n1015), .C1(new_n212), .C2(new_n784), .ZN(new_n1016));
  INV_X1    g0816(.A(G137), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n803), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1006), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT47), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n770), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n960), .A2(new_n769), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n772), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n218), .B2(new_n308), .C1(new_n230), .C2(new_n775), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1021), .A2(new_n764), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n993), .A2(new_n1025), .ZN(G387));
  OAI21_X1  g0826(.A(new_n774), .B1(new_n234), .B2(new_n776), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n243), .A2(new_n218), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1027), .B1(new_n715), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n279), .A2(G50), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT50), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(G68), .A2(G77), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1031), .A2(new_n776), .A3(new_n1032), .A4(new_n715), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1029), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n712), .A2(new_n560), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n772), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n804), .A2(G326), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n823), .A2(new_n586), .B1(new_n817), .B2(G283), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n793), .A2(G317), .B1(G311), .B2(new_n815), .ZN(new_n1039));
  INV_X1    g0839(.A(G322), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1039), .B1(new_n806), .B2(new_n809), .C1(new_n1040), .C2(new_n1001), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT48), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1038), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT114), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g0846(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n1047));
  AOI211_X1 g0847(.A(new_n243), .B(new_n1037), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n532), .B2(new_n784), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n799), .A2(new_n308), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n800), .A2(new_n279), .B1(new_n803), .B2(new_n273), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(G97), .C2(new_n821), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n243), .B1(new_n809), .B2(new_n366), .C1(new_n850), .C2(new_n795), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G50), .B2(new_n793), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n212), .A2(new_n807), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1052), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT113), .Z(new_n1058));
  NAND2_X1  g0858(.A1(new_n1049), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1036), .B1(new_n1059), .B2(new_n770), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1060), .B(new_n764), .C1(new_n705), .C2(new_n769), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n987), .A2(new_n763), .A3(new_n988), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n714), .B1(new_n989), .B2(new_n757), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n990), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1063), .A2(new_n1066), .ZN(G393));
  AOI22_X1  g0867(.A1(new_n793), .A2(G159), .B1(G150), .B2(new_n811), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT51), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n799), .A2(new_n626), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n864), .B1(new_n366), .B2(new_n807), .C1(new_n279), .C2(new_n809), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n1069), .A2(new_n296), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n317), .B2(new_n800), .C1(new_n803), .C2(new_n853), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT116), .Z(new_n1074));
  OAI22_X1  g0874(.A1(new_n851), .A2(new_n808), .B1(new_n1003), .B2(new_n795), .ZN(new_n1075));
  XOR2_X1   g0875(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n1076));
  OR2_X1    g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n800), .A2(new_n806), .B1(new_n803), .B2(new_n1040), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G283), .B2(new_n823), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G294), .B2(new_n1010), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n817), .A2(G116), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1082), .A2(new_n296), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G107), .B2(new_n821), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n770), .B1(new_n1074), .B2(new_n1085), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n950), .A2(new_n769), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1023), .B1(new_n473), .B2(new_n218), .C1(new_n241), .C2(new_n775), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n764), .A4(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n977), .A2(new_n980), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1089), .B1(new_n1090), .B2(new_n762), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n714), .B1(new_n1090), .B2(new_n1065), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1091), .B1(new_n1092), .B2(new_n991), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(G390));
  AOI21_X1  g0894(.A(KEYINPUT38), .B1(new_n883), .B2(new_n891), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT39), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n905), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n910), .A2(new_n911), .B1(new_n890), .B2(new_n914), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n895), .B1(new_n1098), .B2(KEYINPUT38), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1097), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1100), .A2(new_n872), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n869), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n279), .ZN(new_n1103));
  XOR2_X1   g0903(.A(KEYINPUT54), .B(G143), .Z(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1105), .A2(new_n809), .ZN(new_n1106));
  INV_X1    g0906(.A(G125), .ZN(new_n1107));
  INV_X1    g0907(.A(G128), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n243), .B1(new_n803), .B2(new_n1107), .C1(new_n795), .C2(new_n1108), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1106), .B(new_n1109), .C1(G137), .C2(new_n815), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n793), .A2(G132), .B1(G50), .B2(new_n821), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n817), .A2(G159), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n807), .A2(new_n273), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT53), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .A4(new_n1114), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n296), .B1(new_n784), .B2(new_n366), .C1(new_n560), .C2(new_n800), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1070), .B(new_n1116), .C1(G116), .C2(new_n793), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G87), .A2(new_n823), .B1(new_n804), .B2(G294), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1117), .B(new_n1118), .C1(new_n473), .C2(new_n809), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n795), .A2(new_n785), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1115), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n770), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1101), .A2(new_n764), .A3(new_n1103), .A4(new_n1122), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n755), .A2(G330), .A3(new_n838), .A4(new_n900), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n900), .B1(new_n843), .B2(new_n835), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n903), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1100), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n729), .A2(new_n689), .A3(new_n834), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n836), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n903), .B(new_n917), .C1(new_n1130), .C2(new_n900), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1125), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1130), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1099), .B(new_n1127), .C1(new_n1133), .C2(new_n928), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n903), .B1(new_n876), .B2(new_n900), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1134), .B(new_n1124), .C1(new_n1135), .C2(new_n1100), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1123), .B1(new_n1137), .B2(new_n762), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n650), .A2(new_n287), .A3(new_n314), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n459), .B2(new_n460), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n462), .B1(new_n1140), .B2(new_n413), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n456), .A2(KEYINPUT80), .ZN(new_n1142));
  OAI211_X1 g0942(.A(G330), .B(new_n755), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n920), .A2(new_n663), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT118), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n920), .A2(new_n1143), .A3(KEYINPUT118), .A4(new_n663), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n755), .A2(G330), .A3(new_n838), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n928), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n1124), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n876), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n1130), .B2(new_n1151), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1148), .A2(new_n1132), .A3(new_n1136), .A4(new_n1153), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1154), .A2(new_n713), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1150), .A2(new_n1133), .A3(new_n1124), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1150), .A2(new_n1124), .B1(new_n836), .B2(new_n875), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n1137), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1138), .B1(new_n1155), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(G378));
  OAI21_X1  g0964(.A(new_n1148), .B1(new_n1137), .B2(new_n1159), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n650), .A2(new_n287), .ZN(new_n1166));
  XOR2_X1   g0966(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1167));
  XNOR2_X1  g0967(.A(new_n1166), .B(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n324), .A2(new_n686), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1168), .B(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n932), .B2(G330), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n931), .A2(new_n923), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1099), .A2(new_n755), .A3(KEYINPUT40), .A4(new_n929), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1173), .A2(G330), .A3(new_n1174), .A4(new_n1171), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n919), .B1(new_n1172), .B2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1173), .A2(G330), .A3(new_n1174), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1171), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n901), .A2(new_n902), .A3(new_n918), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n1181), .A3(new_n1175), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1177), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1165), .A2(KEYINPUT57), .A3(new_n1183), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1180), .A2(new_n1181), .A3(new_n1175), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1181), .B1(new_n1180), .B2(new_n1175), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT120), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT120), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1177), .A2(new_n1188), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1187), .A2(new_n1189), .B1(new_n1154), .B2(new_n1148), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n713), .B(new_n1184), .C1(new_n1190), .C2(KEYINPUT57), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(KEYINPUT3), .A2(G33), .ZN(new_n1192));
  AOI21_X1  g0992(.A(G50), .B1(new_n1192), .B2(new_n249), .ZN(new_n1193));
  AOI21_X1  g0993(.A(G41), .B1(new_n804), .B2(G124), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n809), .A2(new_n1017), .B1(new_n799), .B2(new_n273), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1105), .A2(new_n807), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(new_n793), .C2(G128), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1197), .B1(new_n1107), .B2(new_n795), .C1(new_n856), .C2(new_n800), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n248), .B(new_n1194), .C1(new_n1198), .C2(KEYINPUT59), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G159), .B2(new_n821), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1193), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1056), .B(new_n249), .C1(new_n366), .C2(new_n799), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n243), .B1(new_n821), .B2(G58), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n785), .B2(new_n803), .C1(new_n308), .C2(new_n809), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(G116), .C2(new_n811), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n473), .B2(new_n800), .C1(new_n560), .C2(new_n851), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT58), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n771), .B1(new_n1202), .B2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n764), .B1(new_n869), .B2(G50), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT119), .Z(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1209), .B(new_n1212), .C1(new_n1171), .C2(new_n767), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1213), .B1(new_n1214), .B2(new_n763), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1191), .A2(new_n1215), .ZN(G375));
  NAND2_X1  g1016(.A1(new_n928), .A2(new_n767), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n809), .A2(new_n273), .B1(new_n799), .B2(new_n317), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT122), .Z(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G132), .B2(new_n811), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n784), .A2(new_n365), .B1(new_n803), .B2(new_n1108), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n296), .B(new_n1221), .C1(new_n815), .C2(new_n1104), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1220), .B(new_n1222), .C1(new_n1017), .C2(new_n851), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G159), .B2(new_n823), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1050), .B1(G77), .B2(new_n821), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n806), .B2(new_n803), .C1(new_n851), .C2(new_n785), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n807), .A2(new_n473), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n811), .A2(G294), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n296), .B1(new_n809), .B2(new_n560), .C1(new_n532), .C2(new_n800), .ZN(new_n1229));
  NOR4_X1   g1029(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n770), .B1(new_n1224), .B2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1217), .A2(new_n764), .A3(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n366), .B2(new_n1102), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1153), .B2(new_n763), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT121), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1156), .A2(new_n1235), .A3(new_n1159), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1235), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1161), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1234), .B1(new_n1238), .B2(new_n970), .ZN(G381));
  INV_X1    g1039(.A(new_n1213), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1188), .B1(new_n1177), .B2(new_n1182), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1186), .A2(KEYINPUT120), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1240), .B1(new_n1243), .B2(new_n762), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1165), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT57), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n714), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1244), .B1(new_n1247), .B2(new_n1184), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1163), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n993), .A2(new_n1093), .A3(new_n1025), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1249), .A2(G381), .A3(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(G384), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(G393), .A2(G396), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .ZN(G407));
  OAI211_X1 g1054(.A(G407), .B(G213), .C1(G343), .C2(new_n1249), .ZN(G409));
  AOI21_X1  g1055(.A(new_n829), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1250), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1093), .B1(new_n993), .B2(new_n1025), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1257), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(G387), .A2(G390), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1257), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(new_n1262), .A3(new_n1250), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1260), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(G375), .A2(G378), .ZN(new_n1265));
  OAI21_X1  g1065(.A(KEYINPUT60), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1156), .A2(new_n1159), .A3(KEYINPUT60), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1267), .A2(new_n713), .A3(new_n1268), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1269), .A2(G384), .A3(new_n1234), .ZN(new_n1270));
  AOI21_X1  g1070(.A(G384), .B1(new_n1269), .B2(new_n1234), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n687), .A2(G213), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1190), .A2(new_n969), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1183), .A2(new_n763), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1163), .A2(new_n1274), .A3(new_n1240), .A4(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1265), .A2(new_n1272), .A3(new_n1273), .A4(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT61), .B1(new_n1277), .B2(KEYINPUT62), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1273), .B(new_n1276), .C1(new_n1248), .C2(new_n1163), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1273), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(G2897), .ZN(new_n1281));
  XOR2_X1   g1081(.A(new_n1281), .B(KEYINPUT125), .Z(new_n1282));
  NAND2_X1  g1082(.A1(new_n1280), .A2(KEYINPUT124), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1282), .B1(new_n1272), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1269), .A2(new_n1234), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1252), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1269), .A2(G384), .A3(new_n1234), .ZN(new_n1287));
  AND4_X1   g1087(.A1(new_n1286), .A2(new_n1287), .A3(new_n1283), .A4(new_n1282), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1279), .B1(new_n1284), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1278), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT123), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1291), .B1(new_n1279), .B2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1280), .B1(G375), .B2(G378), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1294), .A2(KEYINPUT123), .A3(new_n1272), .A4(new_n1276), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT62), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1264), .B1(new_n1290), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT126), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1298), .B1(new_n1284), .B2(new_n1288), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1272), .A2(new_n1283), .A3(new_n1282), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1286), .A2(new_n1287), .A3(new_n1283), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1282), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1300), .A2(new_n1303), .A3(KEYINPUT126), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1299), .A2(new_n1279), .A3(new_n1304), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1294), .A2(KEYINPUT63), .A3(new_n1272), .A4(new_n1276), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1264), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT61), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT63), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1293), .A2(new_n1310), .A3(new_n1295), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1305), .A2(new_n1309), .A3(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1297), .A2(new_n1312), .ZN(G405));
  NAND2_X1  g1113(.A1(new_n1265), .A2(new_n1249), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1260), .A2(new_n1263), .A3(KEYINPUT127), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(KEYINPUT127), .B1(new_n1260), .B2(new_n1263), .ZN(new_n1317));
  NOR3_X1   g1117(.A1(new_n1316), .A2(new_n1272), .A3(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT127), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1263), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1262), .B1(new_n1261), .B2(new_n1250), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1319), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1292), .B1(new_n1322), .B2(new_n1315), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1314), .B1(new_n1318), .B2(new_n1323), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1272), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1322), .A2(new_n1292), .A3(new_n1315), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1325), .A2(new_n1249), .A3(new_n1326), .A4(new_n1265), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1324), .A2(new_n1327), .ZN(G402));
endmodule


