//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n552,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  XOR2_X1   g028(.A(G325), .B(KEYINPUT64), .Z(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT65), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G125), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(KEYINPUT66), .A2(G113), .A3(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(G2105), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT67), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n473));
  OAI211_X1 g048(.A(new_n473), .B(G2105), .C1(new_n465), .C2(new_n470), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n476), .A2(KEYINPUT69), .A3(KEYINPUT3), .A4(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(new_n461), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n462), .A2(KEYINPUT68), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n477), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n481), .A2(G137), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n476), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(G2105), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G101), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n475), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G160));
  NAND2_X1  g064(.A1(new_n481), .A2(new_n482), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G136), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n481), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G124), .ZN(new_n495));
  OR2_X1    g070(.A1(G100), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G112), .C2(new_n482), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n492), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G162));
  NAND3_X1  g074(.A1(new_n481), .A2(G126), .A3(G2105), .ZN(new_n500));
  OR2_X1    g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n501), .B(G2104), .C1(G114), .C2(new_n482), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n482), .A2(G138), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n503), .B1(new_n481), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n503), .A2(new_n482), .A3(G138), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n506), .B1(new_n464), .B2(new_n463), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n500), .B(new_n502), .C1(new_n505), .C2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n517), .A2(new_n523), .ZN(G166));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(G51), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n521), .B2(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(KEYINPUT5), .A2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT5), .A2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n518), .A2(G89), .ZN(new_n532));
  NAND2_X1  g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n528), .A2(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  AOI22_X1  g111(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n516), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n519), .A2(new_n539), .B1(new_n521), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n538), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  AOI22_X1  g118(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n516), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n519), .A2(new_n546), .B1(new_n521), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT70), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  OR2_X1    g131(.A1(KEYINPUT6), .A2(G651), .ZN(new_n557));
  NAND2_X1  g132(.A1(KEYINPUT6), .A2(G651), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n511), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n556), .B1(new_n559), .B2(G53), .ZN(new_n560));
  AND2_X1   g135(.A1(KEYINPUT6), .A2(G651), .ZN(new_n561));
  NOR2_X1   g136(.A1(KEYINPUT6), .A2(G651), .ZN(new_n562));
  OAI211_X1 g137(.A(G53), .B(G543), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT71), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT72), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n567), .B1(new_n529), .B2(new_n530), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n512), .A2(KEYINPUT72), .A3(new_n513), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n514), .A2(new_n518), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G91), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n559), .A2(new_n556), .A3(G53), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT71), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n565), .A2(new_n573), .A3(new_n575), .A4(new_n579), .ZN(G299));
  INV_X1    g155(.A(G166), .ZN(G303));
  NAND2_X1  g156(.A1(new_n574), .A2(G87), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n559), .A2(G49), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G288));
  NAND2_X1  g161(.A1(new_n514), .A2(G61), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT73), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n587), .A2(new_n588), .B1(G73), .B2(G543), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n514), .A2(KEYINPUT73), .A3(G61), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n516), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(G86), .ZN(new_n592));
  INV_X1    g167(.A(G48), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n519), .A2(new_n592), .B1(new_n521), .B2(new_n593), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n591), .A2(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n516), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  INV_X1    g173(.A(G47), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n519), .A2(new_n598), .B1(new_n521), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n568), .A2(new_n569), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G66), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n516), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n559), .A2(G54), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n574), .A2(KEYINPUT10), .A3(G92), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n519), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n608), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n603), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n603), .B1(new_n616), .B2(G868), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  INV_X1    g194(.A(G299), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G297));
  OAI21_X1  g196(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n616), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n629), .B(G2104), .C1(G111), .C2(new_n482), .ZN(new_n630));
  INV_X1    g205(.A(G135), .ZN(new_n631));
  INV_X1    g206(.A(G123), .ZN(new_n632));
  OAI221_X1 g207(.A(new_n630), .B1(new_n490), .B2(new_n631), .C1(new_n632), .C2(new_n493), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT74), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(G2096), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n463), .A2(new_n464), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n485), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT12), .Z(new_n638));
  XOR2_X1   g213(.A(KEYINPUT13), .B(G2100), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n635), .A2(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2430), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT76), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT14), .ZN(new_n649));
  AND2_X1   g224(.A1(new_n649), .A2(KEYINPUT77), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(KEYINPUT77), .ZN(new_n651));
  OAI22_X1  g226(.A1(new_n650), .A2(new_n651), .B1(new_n644), .B2(new_n647), .ZN(new_n652));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(new_n655), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n642), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n656), .A2(new_n642), .A3(new_n657), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(G14), .ZN(new_n664));
  INV_X1    g239(.A(new_n662), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n660), .B1(new_n665), .B2(new_n658), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(KEYINPUT78), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n659), .A2(new_n662), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT78), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(new_n669), .A3(new_n660), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n664), .B1(new_n667), .B2(new_n670), .ZN(G401));
  XOR2_X1   g246(.A(KEYINPUT79), .B(KEYINPUT18), .Z(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT17), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT80), .Z(new_n679));
  XOR2_X1   g254(.A(G2072), .B(G2078), .Z(new_n680));
  INV_X1    g255(.A(new_n672), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n680), .B1(new_n675), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G2096), .B(G2100), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  OR2_X1    g261(.A1(new_n686), .A2(KEYINPUT19), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(KEYINPUT19), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1956), .B(G2474), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1961), .B(G1966), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT20), .Z(new_n694));
  NAND2_X1  g269(.A1(new_n690), .A2(new_n691), .ZN(new_n695));
  INV_X1    g270(.A(new_n692), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n689), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n687), .A2(KEYINPUT81), .A3(new_n688), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(G1991), .B(G1996), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT82), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT83), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n702), .B(new_n707), .Z(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(G229));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NOR2_X1   g285(.A1(G171), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G5), .B2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(G1961), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT96), .ZN(new_n715));
  INV_X1    g290(.A(G2084), .ZN(new_n716));
  NAND2_X1  g291(.A1(G160), .A2(G29), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  AND2_X1   g293(.A1(KEYINPUT24), .A2(G34), .ZN(new_n719));
  NOR2_X1   g294(.A1(KEYINPUT24), .A2(G34), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT93), .Z(new_n722));
  NAND2_X1  g297(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n715), .B1(new_n716), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n710), .A2(G21), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G168), .B2(new_n710), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n712), .A2(new_n713), .B1(G1966), .B2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G28), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(KEYINPUT30), .ZN(new_n729));
  AOI21_X1  g304(.A(G29), .B1(new_n728), .B2(KEYINPUT30), .ZN(new_n730));
  OR2_X1    g305(.A1(KEYINPUT31), .A2(G11), .ZN(new_n731));
  NAND2_X1  g306(.A1(KEYINPUT31), .A2(G11), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n729), .A2(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n727), .B(new_n733), .C1(G1966), .C2(new_n726), .ZN(new_n734));
  INV_X1    g309(.A(new_n723), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n734), .B1(G2084), .B2(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT89), .B(G1348), .Z(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G4), .A2(G16), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT88), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n615), .B2(new_n710), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT90), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n724), .B(new_n736), .C1(new_n738), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n491), .A2(G140), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n494), .A2(G128), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n482), .A2(G116), .ZN(new_n746));
  OAI21_X1  g321(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n744), .B(new_n745), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G29), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n718), .A2(G26), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT92), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT28), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G2067), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n710), .A2(G19), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT91), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n549), .B2(new_n710), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(G1341), .Z(new_n758));
  AND2_X1   g333(.A1(new_n718), .A2(G33), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n482), .A2(G103), .A3(G2104), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT25), .Z(new_n761));
  AOI22_X1  g336(.A1(new_n636), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n762));
  INV_X1    g337(.A(G139), .ZN(new_n763));
  OAI221_X1 g338(.A(new_n761), .B1(new_n762), .B2(new_n482), .C1(new_n763), .C2(new_n490), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n759), .B1(new_n764), .B2(G29), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n766), .A2(G2072), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(G2072), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n758), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n634), .A2(new_n718), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT95), .Z(new_n771));
  NOR4_X1   g346(.A1(new_n743), .A2(new_n754), .A3(new_n769), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n710), .A2(G20), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT23), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n620), .B2(new_n710), .ZN(new_n775));
  INV_X1    g350(.A(G1956), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n718), .A2(G35), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT98), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G162), .B2(new_n718), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT29), .Z(new_n781));
  INV_X1    g356(.A(G2090), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n777), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT99), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n718), .A2(G32), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n491), .A2(G141), .B1(G105), .B2(new_n485), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n494), .A2(G129), .ZN(new_n787));
  NAND3_X1  g362(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT94), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT26), .ZN(new_n790));
  AND3_X1   g365(.A1(new_n786), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n785), .B1(new_n791), .B2(new_n718), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT27), .Z(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(G1996), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n782), .B2(new_n781), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n793), .A2(G1996), .B1(new_n742), .B2(new_n738), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n718), .A2(G27), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G164), .B2(new_n718), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT97), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G2078), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n772), .A2(new_n784), .A3(new_n797), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n710), .A2(G23), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n585), .B2(new_n710), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT33), .B(G1976), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n591), .A2(new_n594), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(G16), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G6), .B2(G16), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT32), .B(G1981), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n806), .A2(KEYINPUT84), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(KEYINPUT84), .B2(new_n806), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n710), .A2(G22), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT85), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G166), .B2(new_n710), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(G1971), .Z(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n809), .B2(new_n811), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT34), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT86), .Z(new_n822));
  OR2_X1    g397(.A1(G25), .A2(G29), .ZN(new_n823));
  OR2_X1    g398(.A1(G95), .A2(G2105), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n824), .B(G2104), .C1(G107), .C2(new_n482), .ZN(new_n825));
  INV_X1    g400(.A(G131), .ZN(new_n826));
  INV_X1    g401(.A(G119), .ZN(new_n827));
  OAI221_X1 g402(.A(new_n825), .B1(new_n490), .B2(new_n826), .C1(new_n827), .C2(new_n493), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n823), .B1(new_n828), .B2(new_n718), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT35), .B(G1991), .Z(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n710), .A2(G24), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n601), .B2(new_n710), .ZN(new_n833));
  INV_X1    g408(.A(G1986), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n829), .A2(new_n830), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI211_X1 g412(.A(new_n831), .B(new_n837), .C1(new_n819), .C2(new_n820), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n822), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT87), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n839), .A2(new_n840), .A3(KEYINPUT36), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(KEYINPUT36), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n822), .A2(new_n842), .A3(new_n838), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n802), .B1(new_n841), .B2(new_n843), .ZN(G311));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n843), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n772), .A2(new_n797), .A3(new_n801), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n845), .A2(new_n784), .A3(new_n846), .ZN(G150));
  NOR2_X1   g422(.A1(new_n615), .A2(new_n623), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT101), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n848), .B(new_n850), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(new_n516), .ZN(new_n853));
  INV_X1    g428(.A(G93), .ZN(new_n854));
  INV_X1    g429(.A(G55), .ZN(new_n855));
  OAI22_X1  g430(.A1(new_n519), .A2(new_n854), .B1(new_n521), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n549), .A2(new_n857), .ZN(new_n858));
  OAI22_X1  g433(.A1(new_n545), .A2(new_n548), .B1(new_n853), .B2(new_n856), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n851), .B(new_n860), .Z(new_n861));
  OR2_X1    g436(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n862));
  INV_X1    g437(.A(G860), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n857), .A2(new_n863), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(G145));
  XNOR2_X1  g443(.A(new_n634), .B(new_n498), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n488), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n791), .B(new_n764), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n491), .A2(G142), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n494), .A2(G130), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n482), .A2(G118), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n872), .B(new_n873), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n638), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n871), .A2(new_n877), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n748), .B(new_n508), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n828), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n878), .A3(new_n879), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n870), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT102), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n870), .B1(new_n884), .B2(new_n885), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n888), .A2(G37), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT103), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(new_n892), .A3(new_n889), .ZN(new_n893));
  XNOR2_X1  g468(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n894), .B1(new_n891), .B2(new_n893), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(G395));
  XNOR2_X1  g472(.A(new_n807), .B(G290), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n585), .B(G166), .Z(new_n899));
  XNOR2_X1  g474(.A(new_n898), .B(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n900), .B(KEYINPUT42), .Z(new_n901));
  XNOR2_X1  g476(.A(new_n625), .B(new_n860), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n616), .A2(G299), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n615), .A2(new_n620), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n904), .B(KEYINPUT105), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n903), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n909), .B1(new_n616), .B2(G299), .ZN(new_n910));
  AOI22_X1  g485(.A1(new_n908), .A2(new_n909), .B1(new_n904), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n906), .B1(new_n911), .B2(new_n902), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT106), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n901), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n912), .A2(new_n913), .ZN(new_n915));
  XOR2_X1   g490(.A(new_n914), .B(new_n915), .Z(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(G868), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(G868), .B2(new_n857), .ZN(G295));
  OAI21_X1  g493(.A(new_n917), .B1(G868), .B2(new_n857), .ZN(G331));
  INV_X1    g494(.A(new_n900), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n860), .B(G301), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(G168), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n905), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT108), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(new_n925), .A3(new_n905), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n905), .A2(new_n909), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n907), .A2(new_n910), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n922), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n920), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n932));
  INV_X1    g507(.A(G37), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n923), .B1(new_n911), .B2(new_n922), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n934), .A2(new_n920), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n931), .A2(new_n932), .A3(new_n933), .A4(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(new_n937), .A3(new_n920), .ZN(new_n938));
  OAI221_X1 g513(.A(new_n923), .B1(KEYINPUT107), .B2(new_n900), .C1(new_n911), .C2(new_n922), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n933), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n936), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n932), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n931), .A2(new_n933), .A3(new_n935), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n943), .B1(new_n944), .B2(new_n932), .ZN(new_n945));
  MUX2_X1   g520(.A(new_n942), .B(new_n945), .S(KEYINPUT44), .Z(G397));
  NOR2_X1   g521(.A1(new_n748), .A2(G2067), .ZN(new_n947));
  INV_X1    g522(.A(G1384), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n481), .A2(new_n504), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n507), .B1(new_n949), .B2(KEYINPUT4), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n500), .A2(new_n502), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT109), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT45), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n475), .A2(G40), .A3(new_n487), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G1996), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT110), .Z(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n748), .B(G2067), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT111), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(new_n960), .B2(new_n791), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n963), .A2(new_n791), .B1(new_n959), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n830), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n828), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n947), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n959), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n828), .A2(new_n968), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n959), .B1(new_n972), .B2(new_n969), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n967), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(G290), .A2(G1986), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n959), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g551(.A(new_n976), .B(KEYINPUT48), .Z(new_n977));
  OAI22_X1  g552(.A1(new_n970), .A2(new_n971), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n971), .B1(new_n965), .B2(new_n791), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n979), .B1(new_n962), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT125), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n982), .B1(new_n963), .B2(KEYINPUT46), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n962), .A2(KEYINPUT125), .A3(new_n980), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n985), .A2(KEYINPUT47), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(KEYINPUT47), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n978), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT123), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n948), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(G2078), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n992), .A2(G40), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n487), .A2(new_n471), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n957), .A2(new_n990), .A3(new_n994), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n475), .A2(G40), .A3(new_n487), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n952), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n998), .A3(new_n990), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n991), .B1(new_n999), .B2(G2078), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n952), .A2(KEYINPUT50), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n508), .A2(new_n1002), .A3(new_n948), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n996), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n713), .ZN(new_n1005));
  AND4_X1   g580(.A1(G301), .A2(new_n995), .A3(new_n1000), .A4(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT122), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n996), .A2(new_n998), .A3(new_n990), .A4(new_n992), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1007), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1000), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1006), .B1(new_n1011), .B2(G171), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n989), .B1(new_n1012), .B2(KEYINPUT54), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1002), .B1(new_n508), .B2(new_n948), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(new_n958), .ZN(new_n1016));
  AOI21_X1  g591(.A(G1961), .B1(new_n1016), .B2(new_n1003), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1008), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT122), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(G301), .B1(new_n1021), .B2(new_n1000), .ZN(new_n1022));
  OAI211_X1 g597(.A(KEYINPUT123), .B(new_n1014), .C1(new_n1022), .C2(new_n1006), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1013), .A2(new_n1023), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n996), .A2(new_n998), .A3(new_n990), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT56), .B(G2072), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1025), .A2(new_n1026), .B1(new_n1004), .B2(new_n776), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n576), .A2(new_n577), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n573), .A2(new_n575), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT116), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1029), .A2(new_n1033), .A3(new_n1030), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT117), .B1(G299), .B2(new_n1030), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n573), .A2(new_n575), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n576), .A2(new_n578), .A3(new_n577), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n578), .B1(new_n576), .B2(new_n577), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1037), .A2(new_n1040), .A3(new_n1041), .A4(KEYINPUT57), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1036), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1035), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1027), .A2(new_n1044), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n958), .A2(G2067), .A3(new_n952), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n738), .B1(new_n1016), .B2(new_n1003), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1045), .B(new_n616), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1044), .A2(KEYINPUT118), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1004), .A2(new_n776), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n996), .A2(new_n998), .A3(new_n990), .A4(new_n1026), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1035), .A2(new_n1043), .A3(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1049), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1048), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n608), .A2(KEYINPUT121), .A3(new_n609), .A4(new_n614), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT60), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n615), .A2(new_n1059), .ZN(new_n1060));
  NOR4_X1   g635(.A1(new_n1047), .A2(new_n1046), .A3(new_n1058), .A4(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1046), .B1(new_n1004), .B2(new_n737), .ZN(new_n1062));
  OR2_X1    g637(.A1(new_n1062), .A2(KEYINPUT60), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1058), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1062), .A2(new_n1064), .B1(new_n1059), .B2(new_n615), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1061), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT61), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(new_n1027), .B2(new_n1044), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1055), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n999), .B2(G1996), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n958), .B1(new_n997), .B2(new_n952), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1072), .A2(KEYINPUT119), .A3(new_n960), .A4(new_n990), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT58), .B(G1341), .Z(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(new_n958), .B2(new_n952), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1071), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n549), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(KEYINPUT59), .A3(new_n549), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1066), .A2(new_n1069), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1036), .A2(new_n1042), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1052), .A2(KEYINPUT120), .A3(new_n1082), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1083), .A2(new_n1045), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n1027), .B2(new_n1044), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT61), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1056), .B1(new_n1081), .B2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(G301), .B(new_n1000), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n995), .A2(new_n1000), .A3(new_n1005), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1014), .B1(new_n1090), .B2(G171), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT49), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT114), .ZN(new_n1094));
  OAI21_X1  g669(.A(G1981), .B1(new_n591), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1095), .A2(new_n807), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n587), .A2(new_n588), .ZN(new_n1097));
  NAND2_X1  g672(.A1(G73), .A2(G543), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(new_n590), .A3(new_n1098), .ZN(new_n1099));
  AOI221_X4 g674(.A(new_n594), .B1(new_n1094), .B2(G1981), .C1(new_n1099), .C2(G651), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1093), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(G1981), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1099), .A2(G651), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n1103), .B2(KEYINPUT114), .ZN(new_n1104));
  NAND2_X1  g679(.A1(G305), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1100), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n1106), .A3(KEYINPUT49), .ZN(new_n1107));
  INV_X1    g682(.A(G8), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1108), .B1(new_n996), .B2(new_n953), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1101), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n585), .A2(G1976), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT52), .ZN(new_n1113));
  INV_X1    g688(.A(G1976), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT52), .B1(G288), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1109), .A2(new_n1111), .A3(new_n1115), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1110), .A2(new_n1113), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT113), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n1004), .B2(G2090), .ZN(new_n1119));
  XOR2_X1   g694(.A(KEYINPUT112), .B(G1971), .Z(new_n1120));
  NAND2_X1  g695(.A1(new_n999), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1016), .A2(KEYINPUT113), .A3(new_n782), .A4(new_n1003), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1119), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(G166), .A2(new_n1108), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(KEYINPUT55), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(G8), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1004), .A2(KEYINPUT115), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT115), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1016), .A2(new_n1128), .A3(new_n1003), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1127), .A2(new_n1129), .A3(new_n782), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1108), .B1(new_n1130), .B2(new_n1121), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1117), .B(new_n1126), .C1(new_n1125), .C2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(G1966), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n999), .A2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n996), .A2(new_n1001), .A3(new_n716), .A4(new_n1003), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1134), .A2(G168), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT51), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1136), .A2(new_n1137), .A3(G8), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(G286), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1140), .A2(G8), .A3(new_n1136), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1138), .B1(new_n1141), .B2(KEYINPUT51), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1092), .A2(new_n1132), .A3(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1024), .A2(new_n1088), .A3(new_n1143), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1123), .A2(G8), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1117), .A2(new_n1145), .A3(new_n1125), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1109), .ZN(new_n1147));
  NOR2_X1   g722(.A1(G288), .A2(G1976), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1110), .A2(new_n1148), .B1(new_n1102), .B2(new_n807), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1146), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n1145), .A2(new_n1125), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1139), .A2(G8), .A3(G168), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT63), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1151), .A2(new_n1126), .A3(new_n1117), .A4(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1153), .B1(new_n1132), .B2(new_n1152), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1150), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1144), .A2(KEYINPUT124), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT124), .B1(new_n1144), .B2(new_n1157), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1141), .A2(KEYINPUT51), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1138), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1022), .B1(new_n1162), .B2(KEYINPUT62), .ZN(new_n1163));
  AOI211_X1 g738(.A(new_n1132), .B(new_n1163), .C1(KEYINPUT62), .C2(new_n1162), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1158), .A2(new_n1159), .A3(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n601), .A2(new_n834), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n959), .B1(new_n975), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n967), .A2(new_n1167), .A3(new_n973), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n988), .B1(new_n1165), .B2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  AOI22_X1  g744(.A1(new_n891), .A2(new_n893), .B1(new_n941), .B2(new_n936), .ZN(new_n1171));
  NOR2_X1   g745(.A1(G227), .A2(new_n458), .ZN(new_n1172));
  INV_X1    g746(.A(new_n1172), .ZN(new_n1173));
  OAI21_X1  g747(.A(KEYINPUT126), .B1(G401), .B2(new_n1173), .ZN(new_n1174));
  AND2_X1   g748(.A1(new_n663), .A2(G14), .ZN(new_n1175));
  AOI21_X1  g749(.A(new_n669), .B1(new_n668), .B2(new_n660), .ZN(new_n1176));
  AOI211_X1 g750(.A(KEYINPUT78), .B(new_n661), .C1(new_n659), .C2(new_n662), .ZN(new_n1177));
  OAI21_X1  g751(.A(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n1179));
  NAND3_X1  g753(.A1(new_n1178), .A2(new_n1179), .A3(new_n1172), .ZN(new_n1180));
  NAND3_X1  g754(.A1(new_n1174), .A2(new_n1180), .A3(new_n708), .ZN(new_n1181));
  NAND2_X1  g755(.A1(new_n1181), .A2(KEYINPUT127), .ZN(new_n1182));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n1183));
  NAND4_X1  g757(.A1(new_n1174), .A2(new_n1180), .A3(new_n1183), .A4(new_n708), .ZN(new_n1184));
  AND3_X1   g758(.A1(new_n1171), .A2(new_n1182), .A3(new_n1184), .ZN(G308));
  NAND3_X1  g759(.A1(new_n1171), .A2(new_n1182), .A3(new_n1184), .ZN(G225));
endmodule


