//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT68), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT68), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n192), .A3(G116), .ZN(new_n193));
  OR3_X1    g007(.A1(new_n189), .A2(KEYINPUT69), .A3(G116), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT69), .B1(new_n189), .B2(G116), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT2), .B(G113), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT70), .ZN(new_n199));
  INV_X1    g013(.A(new_n197), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n200), .A2(new_n193), .A3(new_n194), .A4(new_n195), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n198), .A2(new_n199), .A3(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n196), .A2(KEYINPUT70), .A3(new_n197), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  INV_X1    g020(.A(G134), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT64), .A2(G137), .ZN(new_n208));
  NOR2_X1   g022(.A1(KEYINPUT64), .A2(G137), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G137), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G134), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n206), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n211), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT64), .A2(G137), .ZN(new_n216));
  AND2_X1   g030(.A1(KEYINPUT11), .A2(G134), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(KEYINPUT11), .B1(new_n211), .B2(G134), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(G131), .B1(new_n207), .B2(G137), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT65), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n218), .A2(new_n220), .A3(new_n224), .A4(new_n221), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n213), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G143), .ZN(new_n228));
  INV_X1    g042(.A(G143), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n232), .B(KEYINPUT1), .C1(new_n229), .C2(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G128), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n232), .B1(new_n228), .B2(KEYINPUT1), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n231), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(G143), .B(G146), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT1), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n238), .A3(G128), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n226), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n207), .A2(G137), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n218), .A2(new_n220), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n206), .B1(new_n243), .B2(KEYINPUT66), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n218), .A2(new_n220), .A3(new_n245), .A4(new_n242), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n244), .A2(new_n246), .B1(new_n223), .B2(new_n225), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT0), .ZN(new_n248));
  INV_X1    g062(.A(G128), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n237), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n231), .A2(KEYINPUT0), .A3(G128), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n249), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n241), .B1(new_n247), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT30), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n243), .A2(KEYINPUT66), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(G131), .A3(new_n246), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n223), .A2(new_n225), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n260), .B1(new_n259), .B2(new_n261), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n262), .A2(new_n263), .A3(new_n254), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n240), .B1(new_n226), .B2(new_n265), .ZN(new_n266));
  AOI211_X1 g080(.A(KEYINPUT72), .B(new_n213), .C1(new_n223), .C2(new_n225), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT30), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n205), .B(new_n257), .C1(new_n264), .C2(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT73), .B(G237), .ZN(new_n270));
  INV_X1    g084(.A(G953), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(G210), .A3(new_n271), .ZN(new_n272));
  OR2_X1    g086(.A1(new_n272), .A2(KEYINPUT27), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(KEYINPUT27), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT26), .B(G101), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n273), .A2(new_n274), .A3(new_n276), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n236), .A2(new_n239), .ZN(new_n281));
  INV_X1    g095(.A(new_n213), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n208), .A2(new_n209), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n219), .B1(new_n283), .B2(new_n217), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n224), .B1(new_n284), .B2(new_n221), .ZN(new_n285));
  INV_X1    g099(.A(new_n225), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n281), .B1(new_n287), .B2(KEYINPUT72), .ZN(new_n288));
  INV_X1    g102(.A(new_n267), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n205), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n259), .A2(new_n261), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT71), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n247), .A2(new_n260), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n293), .A3(new_n253), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n280), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n269), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT74), .B1(new_n296), .B2(KEYINPUT31), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(KEYINPUT31), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT31), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n269), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n297), .B1(new_n301), .B2(KEYINPUT74), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT28), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n204), .B1(new_n266), .B2(new_n267), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n303), .B1(new_n264), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT76), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n290), .A2(new_n294), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(KEYINPUT76), .A3(new_n303), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n226), .A2(new_n240), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n254), .B1(new_n259), .B2(new_n261), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n205), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n290), .A2(new_n294), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n255), .A2(KEYINPUT75), .A3(new_n205), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n303), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n280), .B1(new_n310), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n188), .B1(new_n302), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n266), .A2(new_n267), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n205), .B1(new_n264), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n303), .B1(new_n321), .B2(new_n308), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT29), .B1(new_n310), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n313), .A2(new_n314), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n308), .A2(new_n316), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT28), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT29), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n326), .A2(new_n327), .A3(new_n307), .A4(new_n309), .ZN(new_n328));
  INV_X1    g142(.A(new_n280), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n323), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n269), .A2(new_n308), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(new_n329), .ZN(new_n332));
  AOI21_X1  g146(.A(G902), .B1(new_n332), .B2(new_n327), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n319), .A2(KEYINPUT32), .B1(new_n334), .B2(G472), .ZN(new_n335));
  XOR2_X1   g149(.A(KEYINPUT77), .B(KEYINPUT32), .Z(new_n336));
  AND3_X1   g150(.A1(new_n269), .A2(new_n295), .A3(new_n299), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n299), .B1(new_n269), .B2(new_n295), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT74), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n298), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n318), .A3(new_n341), .ZN(new_n342));
  AOI211_X1 g156(.A(KEYINPUT78), .B(new_n336), .C1(new_n342), .C2(new_n187), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n187), .ZN(new_n345));
  INV_X1    g159(.A(new_n336), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n335), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G234), .ZN(new_n349));
  OAI21_X1  g163(.A(G217), .B1(new_n349), .B2(G902), .ZN(new_n350));
  INV_X1    g164(.A(G902), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(G125), .B(G140), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT16), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT16), .ZN(new_n356));
  INV_X1    g170(.A(G140), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n355), .A2(new_n356), .A3(new_n357), .A4(G125), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n357), .A3(G125), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT82), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n354), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n361), .A2(new_n227), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n353), .B(KEYINPUT84), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n227), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n249), .A2(KEYINPUT23), .A3(G119), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n365), .B(KEYINPUT80), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n190), .A2(new_n192), .A3(G128), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT23), .ZN(new_n368));
  OR2_X1    g182(.A1(new_n368), .A2(KEYINPUT81), .ZN(new_n369));
  AOI21_X1  g183(.A(G128), .B1(new_n190), .B2(new_n192), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(new_n368), .B2(KEYINPUT81), .ZN(new_n371));
  AOI211_X1 g185(.A(G110), .B(new_n366), .C1(new_n369), .C2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n367), .B1(new_n189), .B2(G128), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT24), .B(G110), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n362), .B(new_n364), .C1(new_n372), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n361), .A2(new_n227), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT83), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT83), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n361), .A2(new_n380), .A3(new_n227), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n381), .A3(new_n362), .ZN(new_n382));
  OR2_X1    g196(.A1(new_n373), .A2(new_n374), .ZN(new_n383));
  INV_X1    g197(.A(G110), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n366), .B1(new_n369), .B2(new_n371), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n382), .B(new_n383), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n377), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT22), .B(G137), .ZN(new_n388));
  INV_X1    g202(.A(G221), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n389), .A2(new_n349), .A3(G953), .ZN(new_n390));
  XOR2_X1   g204(.A(new_n388), .B(new_n390), .Z(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n391), .B1(new_n377), .B2(new_n386), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT86), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT86), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n397), .B1(new_n393), .B2(new_n394), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n352), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NOR3_X1   g213(.A1(new_n393), .A2(G902), .A3(new_n394), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT85), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(KEYINPUT25), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  NOR4_X1   g218(.A1(new_n393), .A2(new_n394), .A3(G902), .A4(new_n402), .ZN(new_n405));
  OR2_X1    g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n350), .B(KEYINPUT79), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n399), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n270), .A2(G214), .A3(new_n271), .ZN(new_n409));
  XOR2_X1   g223(.A(KEYINPUT95), .B(G143), .Z(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n229), .A2(KEYINPUT95), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n270), .A2(G214), .A3(new_n271), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(KEYINPUT18), .A2(G131), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n206), .B1(new_n411), .B2(new_n413), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT18), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n353), .B(KEYINPUT96), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G146), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n364), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n417), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n418), .A2(KEYINPUT17), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n424), .A2(new_n381), .A3(new_n362), .A4(new_n379), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n411), .A2(new_n206), .A3(new_n413), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n427), .A2(KEYINPUT17), .A3(new_n418), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n423), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(G113), .B(G122), .ZN(new_n430));
  INV_X1    g244(.A(G104), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n430), .B(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT97), .ZN(new_n434));
  AOI21_X1  g248(.A(G902), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n379), .A2(new_n362), .ZN(new_n436));
  INV_X1    g250(.A(new_n418), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT17), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(new_n426), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n436), .A2(new_n439), .A3(new_n381), .A4(new_n424), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n440), .A2(KEYINPUT97), .A3(new_n433), .A4(new_n423), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n435), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G475), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n415), .A2(new_n416), .B1(new_n364), .B2(new_n421), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n432), .B1(new_n444), .B2(new_n419), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n420), .A2(KEYINPUT19), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT19), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n363), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n448), .A3(new_n227), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n449), .B(new_n362), .C1(new_n418), .C2(new_n427), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n429), .A2(new_n432), .B1(new_n445), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT20), .ZN(new_n452));
  NOR2_X1   g266(.A1(G475), .A2(G902), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n452), .B1(new_n451), .B2(new_n453), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n443), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G478), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(KEYINPUT15), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(G116), .B(G122), .ZN(new_n460));
  INV_X1    g274(.A(G107), .ZN(new_n461));
  OR2_X1    g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n461), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n249), .A2(G143), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n229), .A2(G128), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n207), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n465), .A2(KEYINPUT13), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(new_n466), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n465), .A2(KEYINPUT13), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n207), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT98), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n473), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT98), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n462), .A2(new_n463), .B1(new_n207), .B2(new_n467), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G122), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G116), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n461), .B1(new_n481), .B2(KEYINPUT14), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(new_n460), .ZN(new_n483));
  OAI21_X1  g297(.A(G134), .B1(new_n465), .B2(new_n466), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n468), .A2(KEYINPUT99), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT99), .B1(new_n468), .B2(new_n484), .ZN(new_n487));
  OR2_X1    g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n479), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT9), .B(G234), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(G217), .A3(new_n271), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n492), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n479), .A2(new_n488), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n459), .B1(new_n496), .B2(new_n351), .ZN(new_n497));
  AOI211_X1 g311(.A(G902), .B(new_n458), .C1(new_n493), .C2(new_n495), .ZN(new_n498));
  OR2_X1    g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n456), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(G234), .A2(G237), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n501), .A2(G952), .A3(new_n271), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n501), .A2(G902), .A3(G953), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  XOR2_X1   g319(.A(KEYINPUT21), .B(G898), .Z(new_n506));
  OAI21_X1  g320(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n500), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(G469), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n461), .A2(KEYINPUT88), .A3(G104), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n431), .A2(G107), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT88), .B1(new_n461), .B2(G104), .ZN(new_n513));
  OAI21_X1  g327(.A(G101), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT3), .B1(new_n431), .B2(G107), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT3), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n461), .A3(G104), .ZN(new_n517));
  INV_X1    g331(.A(G101), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n515), .A2(new_n517), .A3(new_n518), .A4(new_n511), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n514), .A2(KEYINPUT10), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT90), .B1(new_n281), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n514), .A2(new_n519), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT90), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n522), .A2(new_n240), .A3(new_n523), .A4(KEYINPUT10), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n515), .A2(new_n517), .A3(new_n511), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G101), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(KEYINPUT4), .A3(new_n519), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT4), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n526), .A2(new_n529), .A3(G101), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n249), .B1(new_n228), .B2(KEYINPUT1), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n239), .B1(new_n532), .B2(new_n237), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n519), .A3(new_n514), .ZN(new_n534));
  XOR2_X1   g348(.A(KEYINPUT89), .B(KEYINPUT10), .Z(new_n535));
  AOI22_X1  g349(.A1(new_n531), .A2(new_n253), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n525), .B(new_n536), .C1(new_n263), .C2(new_n262), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n271), .A2(G227), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(KEYINPUT87), .ZN(new_n539));
  XNOR2_X1  g353(.A(G110), .B(G140), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n534), .B1(new_n522), .B2(new_n240), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n292), .A2(new_n293), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT12), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n247), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n545), .A2(new_n546), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n525), .A2(new_n536), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(new_n292), .A3(new_n293), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n542), .B1(new_n551), .B2(new_n537), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n509), .B(new_n351), .C1(new_n549), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(G469), .A2(G902), .ZN(new_n554));
  INV_X1    g368(.A(new_n537), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n541), .B1(new_n548), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n551), .A2(new_n542), .A3(new_n537), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n553), .B(new_n554), .C1(new_n558), .C2(new_n509), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n389), .B1(new_n491), .B2(new_n351), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(G214), .B1(G237), .B2(G902), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n193), .A2(new_n194), .A3(KEYINPUT5), .A4(new_n195), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n566), .B(G113), .C1(KEYINPUT5), .C2(new_n193), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n201), .A3(new_n522), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n528), .A2(new_n530), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n568), .B1(new_n204), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(G110), .B(G122), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n571), .B(new_n568), .C1(new_n204), .C2(new_n569), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(KEYINPUT6), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT6), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n570), .A2(new_n576), .A3(new_n572), .ZN(new_n577));
  INV_X1    g391(.A(G125), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n281), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n254), .A2(G125), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n271), .A2(G224), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n575), .A2(new_n577), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT91), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n575), .A2(new_n583), .A3(KEYINPUT91), .A4(new_n577), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT92), .B(KEYINPUT8), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n571), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n522), .A2(new_n201), .ZN(new_n591));
  OR2_X1    g405(.A1(new_n566), .A2(KEYINPUT93), .ZN(new_n592));
  OAI21_X1  g406(.A(G113), .B1(new_n193), .B2(KEYINPUT5), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(KEYINPUT93), .B2(new_n566), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n591), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n522), .B1(new_n567), .B2(new_n201), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n590), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT7), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n582), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n240), .A2(G125), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n599), .B1(new_n600), .B2(KEYINPUT94), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n601), .B1(new_n581), .B2(KEYINPUT94), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n579), .A2(new_n580), .A3(new_n599), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n597), .A2(new_n602), .A3(new_n574), .A4(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n351), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n588), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(G210), .B1(G237), .B2(G902), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n588), .A2(new_n608), .A3(new_n606), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n565), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n508), .A2(new_n563), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n348), .A2(new_n408), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G101), .ZN(G3));
  NAND2_X1  g429(.A1(new_n342), .A2(new_n351), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(G472), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n617), .A2(new_n408), .A3(new_n563), .A4(new_n345), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT100), .ZN(new_n620));
  INV_X1    g434(.A(new_n495), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n494), .B1(new_n479), .B2(new_n488), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n457), .B(new_n351), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(G478), .A2(G902), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n621), .A2(KEYINPUT33), .A3(new_n622), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n493), .B2(new_n495), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n625), .B1(new_n629), .B2(G478), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n456), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n612), .A2(new_n620), .A3(new_n507), .A4(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n608), .B1(new_n588), .B2(new_n606), .ZN(new_n634));
  AOI211_X1 g448(.A(new_n609), .B(new_n605), .C1(new_n586), .C2(new_n587), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n564), .B(new_n507), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(KEYINPUT100), .B1(new_n636), .B2(new_n631), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n619), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT34), .B(G104), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT101), .B(KEYINPUT102), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  INV_X1    g457(.A(new_n456), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n499), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n636), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n619), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n617), .A2(new_n345), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n407), .B1(new_n404), .B2(new_n405), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n392), .A2(KEYINPUT36), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n387), .B(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n654), .A2(new_n351), .A3(new_n350), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n650), .B1(new_n651), .B2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n617), .A2(KEYINPUT103), .A3(new_n345), .A4(new_n656), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n658), .A2(new_n613), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT104), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT37), .B(G110), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  OR2_X1    g477(.A1(new_n505), .A2(G900), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n503), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n644), .A2(new_n499), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  AND4_X1   g481(.A1(new_n612), .A2(new_n563), .A3(new_n667), .A4(new_n656), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n348), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  NOR2_X1   g484(.A1(new_n634), .A2(new_n635), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT38), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n456), .A2(new_n499), .A3(new_n564), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n672), .A2(new_n656), .A3(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(G472), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n280), .B1(new_n269), .B2(new_n308), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(G902), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n321), .A2(new_n280), .A3(new_n308), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n675), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n679), .B1(new_n319), .B2(KEYINPUT32), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n680), .B1(new_n347), .B2(new_n343), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n665), .B(KEYINPUT39), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n563), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n683), .A2(KEYINPUT40), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(KEYINPUT40), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n674), .A2(new_n681), .A3(new_n684), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G143), .ZN(G45));
  AND3_X1   g501(.A1(new_n563), .A2(new_n612), .A3(new_n656), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n630), .A2(new_n456), .A3(new_n665), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n630), .A2(new_n456), .A3(KEYINPUT105), .A4(new_n665), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n348), .A2(new_n688), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT106), .B(G146), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G48));
  OAI21_X1  g511(.A(new_n351), .B1(new_n549), .B2(new_n552), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(G469), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n699), .A2(new_n700), .A3(new_n553), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n698), .A2(KEYINPUT107), .A3(G469), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n560), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n348), .A2(new_n638), .A3(new_n408), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT41), .B(G113), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G15));
  NAND4_X1  g520(.A1(new_n348), .A2(new_n408), .A3(new_n646), .A4(new_n703), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G116), .ZN(G18));
  AND4_X1   g522(.A1(new_n612), .A2(new_n703), .A3(new_n508), .A4(new_n656), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n348), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  NOR2_X1   g525(.A1(new_n671), .A2(new_n673), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n712), .A2(new_n507), .A3(new_n703), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n675), .B1(new_n342), .B2(new_n351), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n396), .A2(new_n398), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n652), .B1(new_n352), .B2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n301), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n280), .B1(new_n310), .B2(new_n322), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n188), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n714), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n713), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  NOR3_X1   g536(.A1(new_n693), .A2(new_n714), .A3(new_n719), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n703), .A2(new_n612), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n723), .A2(new_n656), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G125), .ZN(G27));
  NAND2_X1  g541(.A1(new_n671), .A2(new_n564), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n693), .A2(new_n728), .A3(new_n562), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n348), .A2(new_n408), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT42), .B1(new_n730), .B2(KEYINPUT108), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n348), .A2(new_n729), .A3(new_n732), .A4(new_n408), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n319), .A2(KEYINPUT32), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n335), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n408), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n729), .A2(KEYINPUT42), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n734), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n716), .B1(new_n735), .B2(new_n335), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n740), .A2(KEYINPUT109), .A3(KEYINPUT42), .A4(new_n729), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n731), .A2(new_n733), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT110), .B(G131), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G33));
  NOR2_X1   g558(.A1(new_n728), .A2(new_n562), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n348), .A2(new_n408), .A3(new_n667), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G134), .ZN(G36));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n509), .B1(new_n558), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n749), .B1(new_n748), .B2(new_n558), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n554), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g567(.A(new_n753), .B(KEYINPUT111), .Z(new_n754));
  INV_X1    g568(.A(new_n553), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n755), .B1(new_n751), .B2(new_n752), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n560), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n682), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n644), .A2(new_n630), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT43), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n651), .A3(new_n656), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n728), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n763), .B1(new_n762), .B2(new_n761), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n758), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G137), .ZN(G39));
  OR4_X1    g580(.A1(new_n348), .A2(new_n408), .A3(new_n693), .A4(new_n728), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n757), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n757), .A2(new_n769), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n768), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G140), .ZN(G42));
  AND2_X1   g587(.A1(new_n669), .A2(new_n726), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n656), .B1(new_n503), .B2(new_n664), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n681), .A2(new_n563), .A3(new_n712), .A4(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n774), .A2(KEYINPUT52), .A3(new_n695), .A4(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT115), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n776), .A2(new_n695), .A3(new_n669), .A4(new_n726), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n730), .A2(KEYINPUT108), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT42), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n786), .A2(new_n787), .A3(new_n733), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n739), .A2(new_n741), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n500), .A2(new_n665), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n723), .B1(new_n348), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n745), .A2(new_n656), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n746), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n645), .A2(new_n631), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(new_n612), .A3(new_n507), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n618), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n660), .A2(new_n614), .A3(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n348), .A2(new_n709), .B1(new_n713), .B2(new_n720), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n704), .A3(new_n707), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n802), .A2(new_n704), .A3(new_n707), .A4(KEYINPUT113), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n790), .A2(new_n801), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n784), .A2(new_n785), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT78), .B1(new_n319), .B2(new_n336), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n345), .A2(new_n344), .A3(new_n346), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n791), .B1(new_n813), .B2(new_n335), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n656), .B(new_n745), .C1(new_n814), .C2(new_n723), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n716), .B1(new_n813), .B2(new_n335), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n798), .B1(new_n816), .B2(new_n613), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n815), .A2(new_n817), .A3(new_n660), .A4(new_n746), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n742), .A2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n805), .A2(new_n806), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(new_n820), .A3(KEYINPUT114), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n777), .A2(new_n781), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n810), .A2(new_n821), .B1(KEYINPUT53), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT54), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n803), .A2(new_n785), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n790), .A2(new_n801), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n784), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n830));
  INV_X1    g644(.A(new_n822), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n830), .B(new_n785), .C1(new_n807), .C2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n830), .B1(new_n823), .B2(new_n785), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n829), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n835), .A2(KEYINPUT54), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n825), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n770), .A2(new_n771), .ZN(new_n838));
  INV_X1    g652(.A(new_n701), .ZN(new_n839));
  INV_X1    g653(.A(new_n702), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n838), .B1(new_n561), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n760), .A2(new_n502), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n844), .A2(new_n720), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n842), .A2(new_n564), .A3(new_n671), .A4(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n703), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT118), .B1(new_n847), .B2(new_n564), .ZN(new_n848));
  OR3_X1    g662(.A1(new_n847), .A2(KEYINPUT118), .A3(new_n564), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n845), .A2(new_n672), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n850), .B(KEYINPUT50), .Z(new_n851));
  NOR2_X1   g665(.A1(new_n847), .A2(new_n728), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n844), .A2(new_n852), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n853), .A2(new_n714), .A3(new_n657), .A4(new_n719), .ZN(new_n854));
  INV_X1    g668(.A(new_n681), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n408), .A2(new_n855), .A3(new_n502), .A4(new_n852), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n630), .A2(new_n456), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n854), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n846), .A2(new_n851), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT51), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n859), .A2(new_n860), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n845), .A2(new_n725), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(G952), .A3(new_n271), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n853), .A2(new_n737), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT48), .ZN(new_n866));
  AOI211_X1 g680(.A(new_n864), .B(new_n866), .C1(new_n632), .C2(new_n856), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n861), .A2(new_n862), .A3(new_n867), .ZN(new_n868));
  OAI22_X1  g682(.A1(new_n837), .A2(new_n868), .B1(G952), .B2(G953), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n841), .B(KEYINPUT49), .Z(new_n870));
  NOR3_X1   g684(.A1(new_n716), .A2(new_n565), .A3(new_n560), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n672), .A2(new_n759), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n872), .A3(new_n855), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n869), .A2(new_n873), .ZN(G75));
  NOR2_X1   g688(.A1(new_n271), .A2(G952), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n827), .B1(new_n778), .B2(new_n783), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n785), .B1(new_n807), .B2(new_n831), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT117), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n877), .B1(new_n879), .B2(new_n832), .ZN(new_n880));
  INV_X1    g694(.A(G210), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n880), .A2(new_n881), .A3(new_n351), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n575), .A2(new_n577), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(new_n583), .ZN(new_n884));
  XOR2_X1   g698(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n885));
  XNOR2_X1  g699(.A(new_n884), .B(new_n885), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n886), .A2(KEYINPUT56), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n876), .B1(new_n882), .B2(new_n887), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n882), .A2(KEYINPUT120), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT56), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n882), .A2(KEYINPUT120), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n888), .B1(new_n892), .B2(new_n886), .ZN(G51));
  XNOR2_X1  g707(.A(new_n835), .B(KEYINPUT54), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n554), .B(KEYINPUT57), .Z(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n896), .B1(new_n552), .B2(new_n549), .ZN(new_n897));
  OR3_X1    g711(.A1(new_n880), .A2(new_n351), .A3(new_n750), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n875), .B1(new_n897), .B2(new_n898), .ZN(G54));
  NAND2_X1  g713(.A1(KEYINPUT58), .A2(G475), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT121), .Z(new_n901));
  NAND3_X1  g715(.A1(new_n835), .A2(G902), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n451), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n876), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n903), .B2(new_n902), .ZN(G60));
  INV_X1    g719(.A(new_n629), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n624), .B(KEYINPUT59), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n906), .B1(new_n837), .B2(new_n907), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n894), .A2(new_n906), .A3(new_n907), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n908), .A2(new_n909), .A3(new_n875), .ZN(G63));
  XNOR2_X1  g724(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n913));
  NAND2_X1  g727(.A1(G217), .A2(G902), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT60), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n880), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n915), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n835), .A2(KEYINPUT122), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n916), .A2(new_n918), .A3(new_n715), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n876), .ZN(new_n920));
  INV_X1    g734(.A(new_n654), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n916), .B2(new_n918), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n912), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n916), .A2(new_n918), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n654), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n925), .A2(new_n876), .A3(new_n919), .A4(new_n911), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n923), .A2(new_n926), .ZN(G66));
  AND3_X1   g741(.A1(new_n820), .A2(new_n660), .A3(new_n817), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n271), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n506), .A2(G224), .A3(G953), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(G898), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n883), .B1(new_n932), .B2(G953), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n931), .B(new_n933), .ZN(G69));
  OAI21_X1  g748(.A(new_n257), .B1(new_n264), .B2(new_n268), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n446), .A2(new_n448), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n935), .B(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n740), .A2(new_n712), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n772), .B1(new_n758), .B2(new_n938), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n774), .A2(new_n695), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n765), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n765), .A2(KEYINPUT125), .A3(new_n940), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n939), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n790), .A2(new_n746), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT126), .ZN(new_n947));
  AOI21_X1  g761(.A(G953), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n271), .A2(G900), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT127), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n948), .A2(KEYINPUT127), .A3(new_n949), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n937), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(G227), .A2(G900), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(G953), .ZN(new_n955));
  INV_X1    g769(.A(new_n937), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n728), .B1(new_n631), .B2(new_n645), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n816), .A2(new_n563), .A3(new_n682), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n765), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT124), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n940), .A2(new_n686), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT62), .Z(new_n962));
  AND3_X1   g776(.A1(new_n960), .A2(new_n772), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n956), .B1(new_n963), .B2(G953), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n953), .A2(new_n955), .A3(new_n964), .ZN(new_n965));
  OR3_X1    g779(.A1(new_n948), .A2(KEYINPUT127), .A3(new_n949), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n950), .ZN(new_n967));
  OAI211_X1 g781(.A(G953), .B(new_n954), .C1(new_n967), .C2(new_n956), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n965), .A2(new_n968), .ZN(G72));
  OR2_X1    g783(.A1(new_n332), .A2(new_n676), .ZN(new_n970));
  NAND2_X1  g784(.A1(G472), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT63), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n876), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n970), .A2(new_n972), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n824), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n963), .A2(new_n676), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n945), .A2(new_n332), .A3(new_n947), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI211_X1 g793(.A(new_n974), .B(new_n976), .C1(new_n979), .C2(new_n928), .ZN(G57));
endmodule


