//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT67), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(KEYINPUT67), .ZN(new_n191));
  OAI21_X1  g005(.A(G119), .B1(new_n189), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n193), .B1(new_n190), .B2(G119), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT66), .A3(G116), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n192), .A2(KEYINPUT5), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT5), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(new_n195), .A3(G116), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n198), .A2(G113), .A3(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT2), .B(G113), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n192), .A2(new_n203), .A3(new_n197), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT3), .B1(new_n206), .B2(G107), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G104), .ZN(new_n210));
  INV_X1    g024(.A(G101), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n206), .A2(G107), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n207), .A2(new_n210), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n209), .A2(G104), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n206), .A2(G107), .ZN(new_n215));
  OAI21_X1  g029(.A(G101), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n205), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT74), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n213), .A2(new_n216), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n201), .A2(new_n204), .A3(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n218), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  XOR2_X1   g036(.A(G110), .B(G122), .Z(new_n223));
  XOR2_X1   g037(.A(new_n223), .B(KEYINPUT8), .Z(new_n224));
  NAND3_X1  g038(.A1(new_n205), .A2(KEYINPUT74), .A3(new_n217), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n207), .A2(new_n210), .A3(new_n212), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G101), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT4), .A3(new_n213), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n230), .A3(G101), .ZN(new_n231));
  INV_X1    g045(.A(new_n204), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n203), .B1(new_n192), .B2(new_n197), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n229), .B(new_n231), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n223), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n221), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G143), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G146), .ZN(new_n238));
  INV_X1    g052(.A(G146), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G143), .ZN(new_n240));
  NAND2_X1  g054(.A1(KEYINPUT0), .A2(G128), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n238), .A2(new_n240), .ZN(new_n243));
  XOR2_X1   g057(.A(KEYINPUT0), .B(G128), .Z(new_n244));
  OAI21_X1  g058(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G125), .ZN(new_n246));
  INV_X1    g060(.A(G128), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(KEYINPUT1), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(new_n238), .A3(new_n240), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(new_n239), .A3(G143), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n237), .B(G146), .C1(new_n247), .C2(KEYINPUT1), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G125), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G224), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G953), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n246), .B(new_n254), .C1(KEYINPUT75), .C2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n256), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT7), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n257), .B(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n226), .A2(new_n236), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n234), .A2(new_n221), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n262), .A2(new_n223), .B1(new_n263), .B2(KEYINPUT6), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(KEYINPUT6), .ZN(new_n265));
  AOI211_X1 g079(.A(new_n235), .B(new_n265), .C1(new_n234), .C2(new_n221), .ZN(new_n266));
  INV_X1    g080(.A(new_n236), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n246), .A2(new_n254), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n269), .B(new_n258), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n187), .B(new_n261), .C1(new_n268), .C2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(G210), .B1(G237), .B2(G902), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n262), .A2(new_n223), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n265), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT6), .A4(new_n223), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(new_n236), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(G902), .B1(new_n279), .B2(new_n270), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(new_n273), .A3(new_n261), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n275), .A2(KEYINPUT76), .A3(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(G214), .B1(G237), .B2(G902), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT76), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n280), .A2(new_n284), .A3(new_n273), .A4(new_n261), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G953), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G952), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n288), .B1(G234), .B2(G237), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT21), .B(G898), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n290), .B(KEYINPUT84), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  AOI211_X1 g106(.A(new_n187), .B(new_n287), .C1(G234), .C2(G237), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n289), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G237), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n287), .A3(G214), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT77), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n297), .A3(G143), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(G143), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n237), .A2(KEYINPUT77), .ZN(new_n300));
  NOR2_X1   g114(.A1(G237), .A2(G953), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n299), .A2(new_n300), .A3(G214), .A4(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G131), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT17), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n298), .A2(new_n302), .A3(G131), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT16), .ZN(new_n309));
  INV_X1    g123(.A(G140), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G125), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n253), .A2(G140), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT70), .ZN(new_n313));
  OR3_X1    g127(.A1(new_n310), .A2(KEYINPUT70), .A3(G125), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n309), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n311), .A2(KEYINPUT16), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n239), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n313), .A2(new_n314), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT16), .ZN(new_n319));
  INV_X1    g133(.A(new_n316), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(G146), .A3(new_n320), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n298), .A2(new_n302), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(KEYINPUT17), .A3(G131), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n308), .A2(new_n317), .A3(new_n321), .A4(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(G113), .B(G122), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(new_n206), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n322), .A2(KEYINPUT18), .A3(G131), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT18), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n303), .A2(new_n328), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n311), .A2(new_n312), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n239), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n318), .B2(new_n239), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n327), .A2(new_n329), .A3(new_n332), .A4(new_n305), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n324), .A2(new_n326), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT79), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n326), .B1(new_n324), .B2(new_n333), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n324), .A2(new_n333), .ZN(new_n339));
  INV_X1    g153(.A(new_n326), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(KEYINPUT79), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n187), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT80), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(G902), .B1(new_n337), .B2(KEYINPUT79), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n344), .B(new_n345), .C1(new_n337), .C2(new_n336), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(G475), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G478), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(KEYINPUT15), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  XOR2_X1   g164(.A(KEYINPUT9), .B(G234), .Z(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G217), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n352), .A2(new_n353), .A3(G953), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(G122), .B1(new_n189), .B2(new_n191), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n190), .A2(G122), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n209), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT81), .B1(new_n247), .B2(G143), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n237), .A3(G128), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G134), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT64), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT64), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G134), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n237), .A2(G128), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n363), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n368), .B1(new_n363), .B2(new_n370), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n359), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT14), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT67), .B(G116), .ZN(new_n375));
  INV_X1    g189(.A(G122), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n374), .B(new_n358), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n190), .A2(KEYINPUT67), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n188), .A2(G116), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT14), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n377), .A2(new_n381), .A3(G107), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT83), .B1(new_n373), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n372), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n363), .A2(new_n368), .A3(new_n370), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n377), .A2(new_n381), .A3(G107), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT83), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .A4(new_n359), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n383), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT13), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n361), .B1(G128), .B2(new_n237), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n247), .A2(KEYINPUT81), .A3(G143), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n360), .A2(new_n362), .A3(KEYINPUT13), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n370), .A3(new_n395), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n396), .A2(KEYINPUT82), .A3(G134), .ZN(new_n397));
  AOI21_X1  g211(.A(KEYINPUT82), .B1(new_n396), .B2(G134), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n209), .B1(new_n356), .B2(new_n358), .ZN(new_n399));
  NOR3_X1   g213(.A1(new_n380), .A2(G107), .A3(new_n357), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n385), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n397), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n355), .B1(new_n390), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT82), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n360), .A2(new_n362), .A3(KEYINPUT13), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT13), .B1(new_n360), .B2(new_n362), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n405), .A2(new_n406), .A3(new_n369), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n404), .B1(new_n407), .B2(new_n364), .ZN(new_n408));
  OAI21_X1  g222(.A(G107), .B1(new_n380), .B2(new_n357), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n371), .B1(new_n409), .B2(new_n359), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n396), .A2(KEYINPUT82), .A3(G134), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n412), .A2(new_n354), .A3(new_n383), .A4(new_n389), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n403), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n350), .B1(new_n414), .B2(new_n187), .ZN(new_n415));
  AOI211_X1 g229(.A(G902), .B(new_n349), .C1(new_n403), .C2(new_n413), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G475), .ZN(new_n418));
  INV_X1    g232(.A(new_n334), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT78), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT19), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT19), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n330), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n420), .B1(new_n424), .B2(G146), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n305), .A2(new_n307), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n421), .A2(new_n423), .A3(KEYINPUT78), .A4(new_n239), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n425), .A2(new_n426), .A3(new_n321), .A4(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n326), .B1(new_n428), .B2(new_n333), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n418), .B(new_n187), .C1(new_n419), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT20), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n428), .A2(new_n333), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n334), .B1(new_n432), .B2(new_n326), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n433), .A2(new_n434), .A3(new_n418), .A4(new_n187), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n347), .A2(new_n417), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n287), .A2(G221), .A3(G234), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(KEYINPUT22), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(G137), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n195), .A2(G128), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n247), .A2(G119), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  XOR2_X1   g258(.A(KEYINPUT24), .B(G110), .Z(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT23), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n443), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n247), .A2(KEYINPUT23), .A3(G119), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n442), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G110), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  AOI211_X1 g267(.A(new_n447), .B(new_n453), .C1(new_n321), .C2(new_n317), .ZN(new_n454));
  OAI22_X1  g268(.A1(new_n451), .A2(G110), .B1(new_n444), .B2(new_n445), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n321), .A2(new_n331), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n441), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n321), .A2(new_n317), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(new_n452), .A3(new_n446), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n456), .A3(new_n440), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(new_n187), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n353), .B1(G234), .B2(new_n187), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT25), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n458), .A2(new_n461), .A3(KEYINPUT25), .A4(new_n187), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n464), .B1(new_n468), .B2(new_n463), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NOR4_X1   g284(.A1(new_n286), .A2(new_n294), .A3(new_n437), .A4(new_n470), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n217), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n252), .A2(new_n213), .A3(new_n216), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT12), .ZN(new_n476));
  INV_X1    g290(.A(G137), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT11), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n368), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(KEYINPUT11), .A3(G134), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT11), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G137), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n479), .A2(new_n484), .A3(new_n304), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n365), .A2(new_n367), .B1(KEYINPUT11), .B2(new_n477), .ZN(new_n486));
  OAI21_X1  g300(.A(G131), .B1(new_n486), .B2(new_n483), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n475), .A2(new_n476), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n476), .B1(new_n475), .B2(new_n488), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT72), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n229), .A2(new_n245), .A3(new_n231), .ZN(new_n493));
  INV_X1    g307(.A(new_n488), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT10), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n495), .B1(new_n220), .B2(new_n252), .ZN(new_n496));
  AND4_X1   g310(.A1(new_n495), .A2(new_n252), .A3(new_n213), .A4(new_n216), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n493), .B(new_n494), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(G110), .B(G140), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(KEYINPUT71), .ZN(new_n500));
  INV_X1    g314(.A(G227), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(G953), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n500), .B(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n491), .A2(new_n492), .A3(new_n498), .A4(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n217), .B(new_n252), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT12), .B1(new_n505), .B2(new_n494), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n475), .A2(new_n476), .A3(new_n488), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n506), .A2(new_n498), .A3(new_n503), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT72), .ZN(new_n509));
  INV_X1    g323(.A(new_n503), .ZN(new_n510));
  INV_X1    g324(.A(new_n498), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n474), .A2(KEYINPUT10), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n220), .A2(new_n495), .A3(new_n252), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n494), .B1(new_n514), .B2(new_n493), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n510), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n504), .A2(new_n509), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G469), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n518), .A3(new_n187), .ZN(new_n519));
  NAND2_X1  g333(.A1(G469), .A2(G902), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n511), .A2(new_n515), .A3(new_n510), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n506), .A2(new_n498), .A3(new_n507), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n510), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(G469), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n519), .A2(new_n520), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(G221), .B1(new_n352), .B2(G902), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G472), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n304), .B1(new_n479), .B2(new_n484), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n486), .A2(G131), .A3(new_n483), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n245), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT65), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(G134), .A2(G137), .ZN(new_n535));
  INV_X1    g349(.A(new_n368), .ZN(new_n536));
  OAI211_X1 g350(.A(G131), .B(new_n535), .C1(new_n536), .C2(G137), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(new_n485), .A3(new_n252), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n488), .A2(KEYINPUT65), .A3(new_n245), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n534), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n232), .A2(new_n233), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n532), .A2(KEYINPUT30), .A3(new_n538), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n542), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT31), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n543), .A2(new_n532), .A3(new_n538), .ZN(new_n549));
  XOR2_X1   g363(.A(KEYINPUT26), .B(G101), .Z(new_n550));
  NAND2_X1  g364(.A1(new_n301), .A2(G210), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n547), .A2(new_n548), .A3(new_n549), .A4(new_n555), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n532), .A2(new_n538), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT28), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n558), .A3(new_n543), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n549), .A2(KEYINPUT28), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n540), .A2(new_n544), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n554), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n556), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n549), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n545), .B1(new_n540), .B2(new_n541), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n566), .B1(new_n567), .B2(new_n544), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n548), .B1(new_n568), .B2(new_n555), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n529), .B(new_n187), .C1(new_n565), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT32), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n547), .A2(new_n549), .A3(new_n555), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT31), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(new_n556), .A3(new_n564), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT32), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n574), .A2(new_n575), .A3(new_n529), .A4(new_n187), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT29), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n563), .B2(new_n554), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n555), .B1(new_n547), .B2(new_n549), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT69), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n559), .A2(new_n560), .B1(new_n540), .B2(new_n544), .ZN(new_n582));
  AOI21_X1  g396(.A(KEYINPUT29), .B1(new_n582), .B2(new_n555), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT69), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n583), .B(new_n584), .C1(new_n568), .C2(new_n555), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n557), .A2(new_n543), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n561), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(new_n554), .ZN(new_n589));
  AOI21_X1  g403(.A(G902), .B1(new_n589), .B2(KEYINPUT29), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n581), .A2(new_n585), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G472), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n528), .B1(new_n577), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n471), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  OAI21_X1  g409(.A(new_n187), .B1(new_n565), .B2(new_n569), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G472), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n597), .A2(new_n570), .A3(new_n527), .A4(new_n526), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(new_n470), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT85), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT87), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n601), .B1(new_n413), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n414), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n403), .B(new_n413), .C1(new_n602), .C2(new_n601), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(G478), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n414), .A2(new_n348), .A3(new_n187), .ZN(new_n607));
  NAND2_X1  g421(.A1(G478), .A2(G902), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n347), .A2(new_n436), .ZN(new_n610));
  INV_X1    g424(.A(new_n294), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n283), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n272), .A2(new_n274), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n614), .B1(new_n615), .B2(KEYINPUT86), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT86), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n275), .A2(new_n617), .A3(new_n281), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n600), .A2(new_n613), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT34), .B(G104), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  INV_X1    g437(.A(new_n417), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n624), .A2(new_n611), .A3(new_n347), .A4(new_n436), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n600), .A2(new_n620), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT88), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT35), .B(G107), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  AND2_X1   g444(.A1(new_n347), .A2(new_n436), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n468), .A2(new_n463), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n460), .A2(new_n456), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n441), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n463), .A2(G902), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n631), .A2(new_n611), .A3(new_n417), .A4(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n598), .A2(new_n639), .A3(new_n286), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT37), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G110), .ZN(G12));
  INV_X1    g456(.A(G900), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n289), .B1(new_n293), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n631), .A2(new_n624), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n616), .A2(new_n618), .A3(new_n638), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n593), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G128), .ZN(G30));
  INV_X1    g465(.A(KEYINPUT91), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n644), .B(KEYINPUT39), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n526), .A2(new_n527), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(new_n655), .B(KEYINPUT90), .Z(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT40), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n655), .B(KEYINPUT90), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT40), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n638), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n283), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n568), .A2(new_n554), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n555), .A2(new_n566), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n187), .B1(new_n665), .B2(new_n586), .ZN(new_n666));
  OAI21_X1  g480(.A(G472), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n577), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(KEYINPUT89), .Z(new_n669));
  AOI21_X1  g483(.A(new_n417), .B1(new_n347), .B2(new_n436), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n282), .A2(new_n285), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT38), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n669), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n652), .B1(new_n662), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n668), .B(KEYINPUT89), .ZN(new_n676));
  INV_X1    g490(.A(new_n670), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n676), .A2(new_n672), .A3(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n678), .A2(KEYINPUT91), .A3(new_n283), .A4(new_n661), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G143), .ZN(G45));
  INV_X1    g495(.A(KEYINPUT92), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n609), .A2(new_n610), .A3(new_n682), .A4(new_n645), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n609), .A2(new_n610), .A3(new_n645), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT92), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n593), .A2(new_n649), .A3(new_n683), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  AOI22_X1  g501(.A1(new_n571), .A2(new_n576), .B1(G472), .B2(new_n591), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n470), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n517), .A2(new_n187), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(G469), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n527), .A3(new_n519), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n619), .A2(new_n612), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT41), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G113), .ZN(G15));
  NOR2_X1   g510(.A1(new_n619), .A2(new_n692), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n577), .A2(new_n592), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n697), .A2(new_n698), .A3(new_n469), .A4(new_n626), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  INV_X1    g514(.A(new_n639), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n697), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G119), .ZN(G21));
  NAND2_X1  g517(.A1(new_n588), .A2(new_n554), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n573), .A2(new_n556), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n529), .A3(new_n187), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n597), .A2(new_n706), .A3(new_n469), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT93), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n597), .A2(new_n706), .A3(KEYINPUT93), .A4(new_n469), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n616), .A2(new_n618), .A3(new_n670), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n692), .A2(new_n294), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n711), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT94), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n712), .B1(new_n709), .B2(new_n710), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT94), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(new_n718), .A3(new_n714), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  NAND3_X1  g535(.A1(new_n597), .A2(new_n706), .A3(new_n638), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT95), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n597), .A2(new_n706), .A3(KEYINPUT95), .A4(new_n638), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n685), .A2(new_n683), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n697), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G125), .ZN(G27));
  NAND3_X1  g543(.A1(new_n698), .A2(KEYINPUT97), .A3(new_n469), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n614), .B1(new_n282), .B2(new_n285), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n685), .A2(new_n683), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT97), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n733), .B1(new_n688), .B2(new_n470), .ZN(new_n734));
  INV_X1    g548(.A(new_n527), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT96), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n524), .B(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n521), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(G469), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n519), .A2(new_n520), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n735), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n730), .A2(new_n732), .A3(new_n734), .A4(new_n741), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n689), .A2(new_n741), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n685), .A2(new_n683), .ZN(new_n744));
  INV_X1    g558(.A(new_n731), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n744), .A2(KEYINPUT42), .A3(new_n745), .ZN(new_n746));
  AOI22_X1  g560(.A1(new_n742), .A2(KEYINPUT42), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G131), .ZN(G33));
  NOR3_X1   g562(.A1(new_n745), .A2(new_n688), .A3(new_n470), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n647), .A3(new_n741), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  NAND3_X1  g565(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n610), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT43), .ZN(new_n754));
  INV_X1    g568(.A(new_n570), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n529), .B1(new_n574), .B2(new_n187), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n754), .B(new_n638), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT98), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n738), .A2(KEYINPUT45), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n521), .B1(new_n510), .B2(new_n523), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n762), .A2(KEYINPUT45), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n761), .A2(G469), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT46), .B1(new_n764), .B2(new_n520), .ZN(new_n765));
  INV_X1    g579(.A(new_n519), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT46), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n764), .A2(new_n520), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n527), .A3(new_n654), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(new_n758), .B2(new_n757), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n760), .A2(new_n731), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G137), .ZN(G39));
  INV_X1    g588(.A(KEYINPUT47), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n769), .A2(new_n768), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n776), .A2(new_n766), .A3(new_n765), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n775), .B1(new_n777), .B2(new_n735), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n770), .A2(KEYINPUT47), .A3(new_n527), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR4_X1   g594(.A1(new_n744), .A2(new_n698), .A3(new_n469), .A4(new_n745), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G140), .ZN(G42));
  NOR4_X1   g597(.A1(new_n688), .A2(new_n648), .A3(new_n646), .A4(new_n528), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n744), .B1(new_n724), .B2(new_n725), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n784), .B1(new_n785), .B2(new_n697), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT100), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n712), .A2(new_n644), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n632), .A2(new_n637), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n668), .A3(new_n789), .A4(new_n741), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n786), .A2(new_n787), .A3(new_n686), .A4(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n728), .A2(new_n650), .A3(new_n686), .A4(new_n790), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT100), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n791), .A2(KEYINPUT52), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT52), .B1(new_n791), .B2(new_n793), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n726), .A2(new_n727), .A3(new_n741), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n789), .A2(new_n437), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n593), .A2(new_n798), .A3(new_n645), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n745), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT99), .ZN(new_n802));
  NOR4_X1   g616(.A1(new_n598), .A2(new_n286), .A3(new_n470), .A4(new_n625), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n802), .B1(new_n803), .B2(new_n640), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n755), .A2(new_n756), .A3(new_n528), .ZN(new_n805));
  INV_X1    g619(.A(new_n286), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(new_n806), .A3(new_n469), .A4(new_n626), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n805), .A2(new_n701), .A3(new_n806), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(KEYINPUT99), .A3(new_n808), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n804), .A2(new_n809), .B1(new_n593), .B2(new_n471), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n805), .A2(new_n806), .A3(new_n469), .A4(new_n613), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n801), .A2(new_n810), .A3(new_n750), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n694), .A2(new_n702), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n716), .B2(new_n719), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n747), .A3(new_n699), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n796), .A2(KEYINPUT53), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT102), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n792), .A2(KEYINPUT52), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n791), .A2(new_n793), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n816), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n826), .A2(KEYINPUT101), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT101), .B1(new_n826), .B2(new_n827), .ZN(new_n829));
  OAI22_X1  g643(.A1(new_n819), .A2(new_n820), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT54), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n754), .A2(KEYINPUT105), .A3(new_n289), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT105), .B1(new_n754), .B2(new_n289), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT106), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n745), .A2(new_n692), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n836), .B1(new_n835), .B2(new_n837), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n730), .A2(new_n734), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT48), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT48), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n841), .A2(new_n845), .A3(new_n842), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n711), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n834), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n697), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n676), .A2(new_n289), .A3(new_n469), .A4(new_n837), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n852), .A2(new_n610), .A3(new_n609), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n691), .A2(new_n735), .A3(new_n519), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n778), .A2(new_n779), .A3(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n855), .A2(new_n731), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n853), .B1(new_n856), .B2(new_n849), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n614), .B(new_n711), .C1(new_n832), .C2(new_n833), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n673), .A2(new_n692), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT50), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n726), .B1(new_n839), .B2(new_n840), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n857), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n851), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n288), .B(KEYINPUT107), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n857), .A2(KEYINPUT51), .A3(new_n861), .A4(new_n862), .ZN(new_n867));
  AND4_X1   g681(.A1(new_n847), .A2(new_n865), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n792), .A2(KEYINPUT100), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n792), .A2(KEYINPUT100), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n824), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n694), .A2(new_n702), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n717), .A2(new_n718), .A3(new_n714), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n718), .B1(new_n717), .B2(new_n714), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n872), .B(new_n699), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n742), .A2(KEYINPUT42), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n743), .A2(new_n746), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n803), .A2(new_n640), .A3(new_n802), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT99), .B1(new_n807), .B2(new_n808), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n594), .B(new_n811), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n750), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n882), .A2(new_n883), .A3(new_n800), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n791), .A2(KEYINPUT52), .A3(new_n793), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n871), .A2(new_n879), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n827), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n827), .B1(new_n815), .B2(KEYINPUT103), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT103), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n814), .A2(new_n747), .A3(new_n889), .A4(new_n699), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n825), .A2(new_n888), .A3(new_n884), .A4(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n887), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT104), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n887), .A2(new_n891), .A3(new_n892), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT104), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n609), .A2(new_n610), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n852), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n831), .A2(new_n868), .A3(new_n898), .A4(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT108), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(G952), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n287), .ZN(new_n905));
  AOI22_X1  g719(.A1(new_n830), .A2(KEYINPUT54), .B1(new_n895), .B2(new_n897), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n906), .A2(KEYINPUT108), .A3(new_n868), .A4(new_n900), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n903), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n669), .A2(new_n614), .ZN(new_n909));
  INV_X1    g723(.A(new_n691), .ZN(new_n910));
  OR3_X1    g724(.A1(new_n910), .A2(KEYINPUT49), .A3(new_n766), .ZN(new_n911));
  OAI21_X1  g725(.A(KEYINPUT49), .B1(new_n910), .B2(new_n766), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n911), .A2(new_n753), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n673), .A2(new_n470), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n909), .A2(new_n913), .A3(new_n914), .A4(new_n527), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n908), .A2(new_n915), .ZN(G75));
  AOI21_X1  g730(.A(KEYINPUT53), .B1(new_n796), .B2(new_n816), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n871), .A2(new_n821), .A3(new_n890), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT103), .B1(new_n875), .B2(new_n878), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n884), .A3(KEYINPUT53), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(new_n187), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(G210), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n279), .B(new_n271), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT109), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT55), .Z(new_n927));
  XNOR2_X1  g741(.A(KEYINPUT110), .B(KEYINPUT56), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n924), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT56), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n927), .B1(new_n924), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n904), .A2(G953), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT111), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n929), .A2(new_n931), .A3(new_n934), .ZN(G51));
  XOR2_X1   g749(.A(new_n520), .B(KEYINPUT57), .Z(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(KEYINPUT54), .B1(new_n917), .B2(new_n921), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n937), .B1(new_n938), .B2(new_n896), .ZN(new_n939));
  INV_X1    g753(.A(new_n517), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT112), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n892), .B1(new_n887), .B2(new_n891), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n936), .B1(new_n893), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT112), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n943), .A2(new_n944), .A3(new_n517), .ZN(new_n945));
  OR3_X1    g759(.A1(new_n922), .A2(new_n187), .A3(new_n764), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n941), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n933), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT113), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n947), .A2(KEYINPUT113), .A3(new_n933), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(G54));
  AND2_X1   g766(.A1(new_n923), .A2(KEYINPUT58), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n433), .B1(new_n953), .B2(G475), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n923), .A2(KEYINPUT58), .A3(G475), .A4(new_n433), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT114), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  AOI211_X1 g772(.A(new_n934), .B(new_n954), .C1(new_n957), .C2(new_n958), .ZN(G60));
  NAND2_X1  g773(.A1(new_n604), .A2(new_n605), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n608), .B(KEYINPUT59), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n960), .B(new_n961), .C1(new_n893), .C2(new_n942), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(KEYINPUT115), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n938), .A2(new_n896), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT115), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n964), .A2(new_n965), .A3(new_n960), .A4(new_n961), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT116), .B1(new_n967), .B2(new_n933), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT116), .ZN(new_n969));
  AOI211_X1 g783(.A(new_n969), .B(new_n934), .C1(new_n963), .C2(new_n966), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n831), .A2(new_n898), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n960), .B1(new_n971), .B2(new_n961), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n968), .A2(new_n970), .A3(new_n972), .ZN(G63));
  XNOR2_X1  g787(.A(KEYINPUT117), .B(KEYINPUT60), .ZN(new_n974));
  NAND2_X1  g788(.A1(G217), .A2(G902), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n922), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n458), .A2(new_n461), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n933), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n980), .B1(new_n635), .B2(new_n977), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT61), .ZN(G66));
  OAI21_X1  g796(.A(G953), .B1(new_n292), .B2(new_n255), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n875), .A2(new_n882), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n983), .B1(new_n984), .B2(G953), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT118), .Z(new_n986));
  OAI21_X1  g800(.A(new_n268), .B1(G898), .B2(new_n287), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n986), .B(new_n987), .Z(G69));
  INV_X1    g802(.A(new_n773), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT62), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n728), .A2(new_n650), .A3(new_n686), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT120), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n680), .A2(KEYINPUT121), .A3(new_n990), .A4(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT121), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n993), .A2(new_n675), .A3(new_n679), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n995), .B1(new_n996), .B2(KEYINPUT62), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n989), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(KEYINPUT122), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT122), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n996), .A2(new_n1001), .A3(KEYINPUT62), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n899), .B1(new_n417), .B2(new_n610), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT123), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1005), .A2(new_n658), .A3(new_n749), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n998), .A2(new_n1003), .A3(new_n782), .A4(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(KEYINPUT119), .B1(new_n1007), .B2(new_n287), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n567), .B(new_n424), .Z(new_n1009));
  OR2_X1    g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(G953), .B1(new_n501), .B2(new_n643), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT119), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1013), .B1(new_n1007), .B2(new_n287), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT125), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n883), .B1(new_n780), .B2(new_n781), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n773), .A2(new_n993), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n842), .A2(new_n713), .ZN(new_n1018));
  OR2_X1    g832(.A1(new_n771), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n747), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1015), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(new_n1022));
  NOR3_X1   g836(.A1(new_n1017), .A2(new_n1015), .A3(new_n1020), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n287), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n643), .A2(G953), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT124), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1024), .A2(new_n1009), .A3(new_n1027), .ZN(new_n1028));
  OR2_X1    g842(.A1(new_n1014), .A2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1030));
  OAI211_X1 g844(.A(new_n1010), .B(new_n1012), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  NOR3_X1   g845(.A1(new_n1014), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1011), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1031), .A2(new_n1034), .ZN(G72));
  NAND2_X1  g849(.A1(G472), .A2(G902), .ZN(new_n1036));
  XOR2_X1   g850(.A(new_n1036), .B(KEYINPUT63), .Z(new_n1037));
  INV_X1    g851(.A(new_n984), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1037), .B1(new_n1007), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g853(.A(KEYINPUT126), .ZN(new_n1040));
  AND2_X1   g854(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1042));
  INV_X1    g856(.A(new_n663), .ZN(new_n1043));
  NOR3_X1   g857(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  AND2_X1   g858(.A1(new_n568), .A2(new_n555), .ZN(new_n1045));
  OAI211_X1 g859(.A(new_n830), .B(new_n1037), .C1(new_n1045), .C2(new_n580), .ZN(new_n1046));
  INV_X1    g860(.A(new_n1023), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1047), .A2(new_n984), .A3(new_n1021), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1048), .A2(new_n1037), .ZN(new_n1049));
  OAI211_X1 g863(.A(new_n547), .B(new_n664), .C1(new_n1049), .C2(KEYINPUT127), .ZN(new_n1050));
  AND2_X1   g864(.A1(new_n1049), .A2(KEYINPUT127), .ZN(new_n1051));
  OAI211_X1 g865(.A(new_n933), .B(new_n1046), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g866(.A1(new_n1044), .A2(new_n1052), .ZN(G57));
endmodule


