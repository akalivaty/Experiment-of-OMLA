//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n192), .A3(new_n195), .A4(new_n190), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(KEYINPUT0), .A2(G128), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT0), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT65), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT0), .A3(G128), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n198), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT67), .B1(new_n205), .B2(G143), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G146), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n208), .B2(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n205), .A2(KEYINPUT66), .A3(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n204), .B1(new_n210), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G143), .B(G146), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT0), .A3(G128), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n197), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT68), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n190), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n188), .A2(G137), .ZN(new_n222));
  OAI21_X1  g036(.A(G131), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n205), .A2(G143), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n200), .B1(new_n224), .B2(KEYINPUT1), .ZN(new_n225));
  INV_X1    g039(.A(new_n214), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n206), .A2(new_n209), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n216), .A2(G128), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n223), .B(new_n196), .C1(new_n228), .C2(new_n230), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n197), .A2(new_n215), .A3(KEYINPUT68), .A4(new_n217), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n220), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  XOR2_X1   g047(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n234));
  AND3_X1   g048(.A1(new_n233), .A2(KEYINPUT69), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT69), .B1(new_n233), .B2(new_n234), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n231), .A2(KEYINPUT30), .A3(new_n218), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NOR3_X1   g052(.A1(new_n235), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT70), .ZN(new_n240));
  XOR2_X1   g054(.A(G116), .B(G119), .Z(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT2), .B(G113), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n241), .B(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n239), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n233), .A2(new_n234), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n233), .A2(KEYINPUT69), .A3(new_n234), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n247), .A2(new_n243), .A3(new_n237), .A4(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT70), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n244), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G237), .ZN(new_n252));
  INV_X1    g066(.A(G953), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(G210), .ZN(new_n254));
  XOR2_X1   g068(.A(new_n254), .B(G101), .Z(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n256));
  XOR2_X1   g070(.A(new_n255), .B(new_n256), .Z(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n243), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n231), .A2(new_n259), .A3(new_n218), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n251), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n260), .B(KEYINPUT28), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n233), .A2(new_n243), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n257), .B1(new_n265), .B2(KEYINPUT29), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT29), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G902), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n231), .A2(new_n218), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n243), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n263), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n268), .B1(new_n266), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(G472), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n260), .A2(new_n257), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n240), .B1(new_n239), .B2(new_n243), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n249), .A2(KEYINPUT70), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT31), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n265), .A2(new_n258), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n280), .B(KEYINPUT71), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT31), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n251), .A2(new_n282), .A3(new_n275), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n279), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(G472), .A2(G902), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT32), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT32), .ZN(new_n289));
  AOI211_X1 g103(.A(KEYINPUT72), .B(new_n289), .C1(new_n284), .C2(new_n285), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n273), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(G125), .B(G140), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT16), .ZN(new_n293));
  INV_X1    g107(.A(G125), .ZN(new_n294));
  OR3_X1    g108(.A1(new_n294), .A2(KEYINPUT16), .A3(G140), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n205), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n293), .A2(G146), .A3(new_n295), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n200), .A2(G119), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g116(.A1(new_n200), .A2(G119), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G110), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n303), .A2(new_n300), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT24), .B(G110), .Z(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n299), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  XOR2_X1   g124(.A(KEYINPUT74), .B(G110), .Z(new_n311));
  OAI22_X1  g125(.A1(new_n307), .A2(new_n308), .B1(new_n305), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n292), .A2(new_n205), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n298), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT22), .B(G137), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n316), .B(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G221), .ZN(new_n319));
  INV_X1    g133(.A(G234), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n319), .A2(new_n320), .A3(G953), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n318), .B(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n315), .B(new_n322), .ZN(new_n323));
  OR3_X1    g137(.A1(new_n323), .A2(KEYINPUT25), .A3(G902), .ZN(new_n324));
  XOR2_X1   g138(.A(KEYINPUT73), .B(G217), .Z(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n320), .B2(G902), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT25), .B1(new_n323), .B2(G902), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n324), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  OR2_X1    g143(.A1(new_n329), .A2(KEYINPUT77), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(KEYINPUT77), .ZN(new_n331));
  INV_X1    g145(.A(new_n323), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(new_n268), .A3(new_n326), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT90), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n297), .A2(new_n298), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n252), .A2(new_n253), .A3(G214), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(G143), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(new_n195), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT17), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n339), .B(new_n195), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n337), .B(new_n341), .C1(new_n342), .C2(KEYINPUT17), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(KEYINPUT18), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT18), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n339), .B1(new_n345), .B2(new_n195), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n292), .B(new_n205), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(G113), .B(G122), .ZN(new_n350));
  INV_X1    g164(.A(G104), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n350), .B(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n336), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n343), .A2(KEYINPUT90), .A3(new_n352), .A4(new_n348), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n292), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT19), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n292), .B1(KEYINPUT87), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT88), .B1(new_n361), .B2(G146), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT88), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n358), .A2(new_n363), .A3(new_n205), .A4(new_n360), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n342), .A2(new_n362), .A3(new_n298), .A4(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n348), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT89), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n365), .A2(KEYINPUT89), .A3(new_n348), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n353), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n356), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G475), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(new_n268), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT20), .ZN(new_n374));
  AOI21_X1  g188(.A(G475), .B1(new_n356), .B2(new_n370), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT20), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(new_n268), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT91), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n352), .B1(new_n349), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n379), .B1(new_n378), .B2(new_n349), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n356), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n268), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n374), .A2(new_n377), .B1(G475), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G116), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(KEYINPUT14), .A3(G122), .ZN(new_n385));
  XOR2_X1   g199(.A(G116), .B(G122), .Z(new_n386));
  OAI211_X1 g200(.A(G107), .B(new_n385), .C1(new_n386), .C2(KEYINPUT14), .ZN(new_n387));
  OR2_X1    g201(.A1(new_n387), .A2(KEYINPUT92), .ZN(new_n388));
  OR2_X1    g202(.A1(new_n386), .A2(G107), .ZN(new_n389));
  XNOR2_X1  g203(.A(G128), .B(G143), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(new_n188), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n387), .A2(KEYINPUT92), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n388), .A2(new_n389), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n386), .A2(G107), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n390), .A2(new_n188), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n188), .B1(new_n390), .B2(KEYINPUT13), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n208), .A2(G128), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n397), .B1(KEYINPUT13), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n395), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n393), .A2(new_n400), .ZN(new_n401));
  XOR2_X1   g215(.A(KEYINPUT9), .B(G234), .Z(new_n402));
  NAND3_X1  g216(.A1(new_n325), .A2(new_n402), .A3(new_n253), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n403), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n268), .ZN(new_n407));
  INV_X1    g221(.A(G478), .ZN(new_n408));
  OR2_X1    g222(.A1(new_n408), .A2(KEYINPUT15), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n407), .B(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(G234), .A2(G237), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(G952), .A3(new_n253), .ZN(new_n412));
  XOR2_X1   g226(.A(new_n412), .B(KEYINPUT93), .Z(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  XOR2_X1   g228(.A(KEYINPUT21), .B(G898), .Z(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n411), .A2(G902), .A3(G953), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n414), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n383), .A2(new_n410), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n351), .A2(G107), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT78), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n422), .B(new_n423), .ZN(new_n424));
  XOR2_X1   g238(.A(KEYINPUT79), .B(G101), .Z(new_n425));
  OAI21_X1  g239(.A(KEYINPUT3), .B1(new_n351), .B2(G107), .ZN(new_n426));
  OR3_X1    g240(.A1(new_n351), .A2(KEYINPUT3), .A3(G107), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n424), .A2(new_n425), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n422), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n351), .A2(G107), .ZN(new_n430));
  OAI21_X1  g244(.A(G101), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n228), .A2(new_n230), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT81), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n225), .A2(new_n216), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n428), .B(new_n431), .C1(new_n230), .C2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT81), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n432), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n435), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n197), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT12), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n215), .A2(new_n217), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n444));
  AOI22_X1  g258(.A1(KEYINPUT4), .A2(new_n428), .B1(new_n444), .B2(G101), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n444), .A2(KEYINPUT4), .A3(G101), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n428), .A2(new_n431), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n448), .B(KEYINPUT10), .C1(new_n228), .C2(new_n230), .ZN(new_n449));
  INV_X1    g263(.A(new_n197), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT80), .B(KEYINPUT10), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n437), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n447), .A2(new_n449), .A3(new_n450), .A4(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(G110), .B(G140), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n253), .A2(G227), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n454), .B(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT12), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n440), .A2(new_n457), .A3(new_n197), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n442), .A2(new_n453), .A3(new_n456), .A4(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n447), .A2(new_n449), .A3(new_n452), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n197), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n453), .ZN(new_n462));
  INV_X1    g276(.A(new_n456), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G469), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n268), .ZN(new_n467));
  NAND2_X1  g281(.A1(G469), .A2(G902), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n461), .A2(new_n453), .A3(new_n456), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n442), .A2(new_n453), .A3(new_n458), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n469), .B1(new_n470), .B2(new_n456), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n467), .B(new_n468), .C1(new_n466), .C2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n319), .B1(new_n402), .B2(new_n268), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n443), .A2(new_n294), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n433), .A2(new_n294), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n253), .A2(G224), .ZN(new_n479));
  XOR2_X1   g293(.A(new_n478), .B(new_n479), .Z(new_n480));
  INV_X1    g294(.A(G113), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n384), .A2(G119), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n484), .B1(new_n241), .B2(new_n482), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(KEYINPUT83), .ZN(new_n486));
  OR2_X1    g300(.A1(new_n241), .A2(new_n242), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n487), .A3(new_n448), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n243), .B1(new_n445), .B2(new_n446), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XOR2_X1   g304(.A(G110), .B(G122), .Z(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n491), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n488), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(KEYINPUT6), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n490), .A2(new_n496), .A3(new_n491), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n480), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n479), .A2(KEYINPUT7), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n478), .A2(new_n499), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n500), .A2(KEYINPUT86), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n476), .A2(KEYINPUT7), .A3(new_n479), .A4(new_n477), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n494), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n486), .A2(new_n487), .A3(new_n432), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT5), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n484), .B1(new_n505), .B2(new_n241), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT85), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n506), .A2(new_n507), .A3(new_n487), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n507), .B1(new_n506), .B2(new_n487), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n448), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT84), .B(KEYINPUT8), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n491), .B(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n504), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n500), .A2(KEYINPUT86), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n501), .A2(new_n503), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n498), .A2(new_n515), .A3(new_n268), .ZN(new_n516));
  OAI21_X1  g330(.A(G210), .B1(G237), .B2(G902), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n498), .A2(new_n515), .A3(new_n268), .A4(new_n517), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(G214), .B1(G237), .B2(G902), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n421), .A2(new_n475), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n291), .A2(new_n335), .A3(new_n524), .ZN(new_n525));
  XOR2_X1   g339(.A(new_n525), .B(new_n425), .Z(G3));
  INV_X1    g340(.A(G472), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n527), .B1(new_n284), .B2(new_n268), .ZN(new_n528));
  INV_X1    g342(.A(new_n285), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n282), .B1(new_n251), .B2(new_n275), .ZN(new_n530));
  AOI211_X1 g344(.A(KEYINPUT31), .B(new_n274), .C1(new_n244), .C2(new_n250), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n529), .B1(new_n532), .B2(new_n281), .ZN(new_n533));
  NOR4_X1   g347(.A1(new_n528), .A2(new_n533), .A3(new_n334), .A4(new_n475), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n407), .A2(new_n408), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n401), .A2(KEYINPUT95), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT95), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n393), .A2(new_n538), .A3(new_n400), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n403), .A3(new_n539), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n540), .A2(KEYINPUT96), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n404), .B1(new_n540), .B2(KEYINPUT96), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT33), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n406), .A2(KEYINPUT33), .ZN(new_n544));
  AOI21_X1  g358(.A(G902), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n536), .B1(new_n545), .B2(G478), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n382), .A2(G475), .ZN(new_n548));
  INV_X1    g362(.A(new_n377), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n376), .B1(new_n375), .B2(new_n268), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT94), .B1(new_n521), .B2(new_n522), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT94), .ZN(new_n554));
  INV_X1    g368(.A(new_n522), .ZN(new_n555));
  AOI211_X1 g369(.A(new_n554), .B(new_n555), .C1(new_n519), .C2(new_n520), .ZN(new_n556));
  NOR4_X1   g370(.A1(new_n552), .A2(new_n553), .A3(new_n556), .A4(new_n419), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n534), .A2(new_n557), .ZN(new_n558));
  XOR2_X1   g372(.A(KEYINPUT34), .B(G104), .Z(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(G6));
  INV_X1    g374(.A(KEYINPUT97), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n374), .A2(new_n561), .A3(new_n377), .ZN(new_n562));
  INV_X1    g376(.A(new_n410), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n550), .A2(KEYINPUT97), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n562), .A2(new_n563), .A3(new_n548), .A4(new_n564), .ZN(new_n565));
  NOR4_X1   g379(.A1(new_n553), .A2(new_n556), .A3(new_n565), .A4(new_n419), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n534), .A2(new_n566), .ZN(new_n567));
  XOR2_X1   g381(.A(KEYINPUT35), .B(G107), .Z(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(G9));
  NOR2_X1   g383(.A1(new_n322), .A2(KEYINPUT36), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(new_n315), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(new_n268), .A3(new_n326), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n330), .A2(new_n331), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(G902), .B1(new_n532), .B2(new_n281), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n286), .B(new_n573), .C1(new_n574), .C2(new_n527), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT98), .ZN(new_n576));
  INV_X1    g390(.A(new_n528), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT98), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n577), .A2(new_n578), .A3(new_n286), .A4(new_n573), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n576), .A2(new_n524), .A3(new_n579), .ZN(new_n580));
  XOR2_X1   g394(.A(KEYINPUT37), .B(G110), .Z(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT99), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n580), .B(new_n582), .ZN(G12));
  NAND3_X1  g397(.A1(new_n573), .A2(new_n474), .A3(new_n472), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n584), .A2(new_n553), .A3(new_n556), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n291), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G900), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n414), .B1(new_n587), .B2(new_n418), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n565), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G128), .ZN(G30));
  XNOR2_X1  g405(.A(new_n588), .B(KEYINPUT39), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n475), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT40), .ZN(new_n594));
  INV_X1    g408(.A(new_n573), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n258), .B1(new_n251), .B2(new_n260), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n261), .A2(new_n270), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n268), .ZN(new_n598));
  OAI21_X1  g412(.A(G472), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n599), .B1(new_n288), .B2(new_n290), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n521), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n551), .A2(new_n563), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n602), .A2(new_n555), .A3(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n594), .A2(new_n595), .A3(new_n600), .A4(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G143), .ZN(G45));
  NOR2_X1   g420(.A1(new_n552), .A2(new_n588), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n586), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G146), .ZN(G48));
  INV_X1    g423(.A(new_n465), .ZN(new_n610));
  OAI21_X1  g424(.A(G469), .B1(new_n610), .B2(G902), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n611), .A2(new_n467), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n474), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n291), .A2(new_n557), .A3(new_n335), .A4(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT41), .B(G113), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT101), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n615), .B(new_n617), .ZN(G15));
  NAND4_X1  g432(.A1(new_n291), .A2(new_n335), .A3(new_n566), .A4(new_n614), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G116), .ZN(G18));
  NOR2_X1   g434(.A1(new_n595), .A2(new_n421), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n613), .A2(new_n553), .A3(new_n556), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n291), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G119), .ZN(G21));
  NOR4_X1   g438(.A1(new_n553), .A2(new_n556), .A3(new_n603), .A4(new_n419), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n271), .A2(new_n258), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n279), .A2(new_n283), .A3(new_n626), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n627), .A2(KEYINPUT102), .A3(new_n285), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT102), .B1(new_n627), .B2(new_n285), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n628), .A2(new_n528), .A3(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n625), .A2(new_n630), .A3(new_n335), .A4(new_n614), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G122), .ZN(G24));
  NAND4_X1  g446(.A1(new_n630), .A2(new_n573), .A3(new_n607), .A4(new_n622), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G125), .ZN(G27));
  NAND2_X1  g448(.A1(new_n471), .A2(KEYINPUT103), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n469), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n467), .B(new_n468), .C1(new_n638), .C2(new_n466), .ZN(new_n639));
  INV_X1    g453(.A(new_n521), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n473), .A2(new_n555), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n291), .A2(new_n335), .A3(new_n607), .A4(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT42), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n642), .A2(new_n552), .A3(new_n588), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n648), .B1(new_n533), .B2(KEYINPUT32), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n533), .A2(KEYINPUT32), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n286), .A2(KEYINPUT104), .A3(new_n289), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n649), .A2(new_n273), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n647), .A2(new_n652), .A3(KEYINPUT42), .A4(new_n335), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT105), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n646), .A2(KEYINPUT105), .A3(new_n653), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G131), .ZN(G33));
  NAND4_X1  g473(.A1(new_n291), .A2(new_n335), .A3(new_n589), .A4(new_n643), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G134), .ZN(G36));
  INV_X1    g475(.A(KEYINPUT45), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n471), .A2(new_n662), .ZN(new_n663));
  OAI211_X1 g477(.A(G469), .B(new_n663), .C1(new_n638), .C2(new_n662), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n468), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT46), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n664), .A2(KEYINPUT46), .A3(new_n468), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n667), .A2(new_n467), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n474), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n592), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n546), .A2(new_n551), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n672), .A2(KEYINPUT43), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(KEYINPUT43), .ZN(new_n674));
  OAI221_X1 g488(.A(new_n573), .B1(new_n533), .B2(new_n528), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n521), .A2(new_n555), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n671), .A2(new_n677), .A3(new_n678), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G137), .ZN(G39));
  OAI21_X1  g495(.A(new_n670), .B1(KEYINPUT106), .B2(KEYINPUT47), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n291), .A2(new_n335), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n669), .A2(new_n474), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n679), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n552), .A2(new_n687), .A3(new_n588), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n682), .A2(new_n683), .A3(new_n686), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G140), .ZN(G42));
  AND2_X1   g504(.A1(new_n647), .A2(KEYINPUT42), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n652), .A2(new_n335), .ZN(new_n692));
  AOI22_X1  g506(.A1(new_n691), .A2(new_n692), .B1(new_n644), .B2(new_n645), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n615), .A2(new_n619), .A3(new_n623), .A4(new_n631), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT53), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n547), .A2(new_n697), .A3(new_n551), .ZN(new_n698));
  OAI21_X1  g512(.A(KEYINPUT107), .B1(new_n546), .B2(new_n383), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n698), .B(new_n699), .C1(new_n410), .C2(new_n551), .ZN(new_n700));
  INV_X1    g514(.A(new_n523), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n534), .A2(new_n420), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n702), .A2(new_n525), .A3(new_n580), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n584), .A2(new_n563), .A3(new_n588), .ZN(new_n704));
  AND4_X1   g518(.A1(new_n548), .A2(new_n679), .A3(new_n564), .A4(new_n562), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n291), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n660), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n647), .A2(new_n630), .A3(new_n573), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n703), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n291), .B(new_n585), .C1(new_n589), .C2(new_n607), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n553), .A2(new_n556), .A3(new_n603), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n573), .A2(new_n588), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n712), .A2(new_n639), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n600), .A2(new_n474), .A3(new_n711), .A4(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n710), .A2(new_n714), .A3(new_n633), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT52), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n710), .A2(new_n714), .A3(KEYINPUT52), .A4(new_n633), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n696), .A2(new_n709), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n696), .A2(new_n709), .A3(new_n719), .A4(KEYINPUT109), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n719), .A2(KEYINPUT108), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n709), .ZN(new_n726));
  INV_X1    g540(.A(new_n694), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n717), .A2(new_n728), .A3(new_n718), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n658), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n695), .B1(new_n726), .B2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT54), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n724), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT53), .B1(new_n726), .B2(new_n730), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n703), .A2(new_n707), .A3(new_n708), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n717), .B2(new_n718), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n736), .A2(new_n695), .A3(new_n658), .A4(new_n727), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n734), .A2(KEYINPUT54), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n673), .A2(new_n674), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n614), .A2(new_n414), .A3(new_n679), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n692), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT114), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT48), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n630), .A2(new_n335), .A3(new_n414), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n614), .A2(new_n602), .ZN(new_n748));
  NOR4_X1   g562(.A1(new_n747), .A2(new_n522), .A3(new_n741), .A4(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n750), .A2(KEYINPUT110), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT110), .B1(new_n750), .B2(new_n751), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n750), .A2(KEYINPUT111), .A3(new_n751), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n755), .B1(new_n749), .B2(KEYINPUT50), .ZN(new_n756));
  OAI22_X1  g570(.A1(new_n752), .A2(new_n753), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n747), .A2(new_n741), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n682), .A2(new_n686), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n612), .A2(new_n473), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n600), .A2(new_n742), .A3(new_n334), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n383), .A3(new_n546), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT112), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n762), .A2(new_n679), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n743), .A2(new_n573), .A3(new_n630), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n757), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n757), .A2(new_n768), .A3(KEYINPUT51), .A4(new_n769), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n758), .A2(new_n622), .ZN(new_n774));
  XOR2_X1   g588(.A(new_n774), .B(KEYINPUT113), .Z(new_n775));
  INV_X1    g589(.A(new_n763), .ZN(new_n776));
  OAI211_X1 g590(.A(G952), .B(new_n253), .C1(new_n776), .C2(new_n552), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n772), .A2(new_n773), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n740), .A2(new_n746), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT115), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n740), .A2(new_n779), .A3(new_n782), .A4(new_n746), .ZN(new_n783));
  OR2_X1    g597(.A1(G952), .A2(G953), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n781), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n612), .B(KEYINPUT49), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n786), .A2(new_n641), .A3(new_n672), .ZN(new_n787));
  INV_X1    g601(.A(new_n600), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n787), .A2(new_n788), .A3(new_n335), .A4(new_n602), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n785), .A2(new_n789), .ZN(G75));
  AND2_X1   g604(.A1(new_n724), .A2(new_n731), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n268), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT56), .B1(new_n792), .B2(G210), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n495), .A2(new_n497), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(new_n480), .ZN(new_n795));
  XNOR2_X1  g609(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n795), .B(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n793), .A2(new_n797), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n253), .A2(G952), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(G51));
  XOR2_X1   g615(.A(new_n468), .B(KEYINPUT117), .Z(new_n802));
  XOR2_X1   g616(.A(new_n802), .B(KEYINPUT57), .Z(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT109), .B1(new_n736), .B2(new_n696), .ZN(new_n805));
  INV_X1    g619(.A(new_n723), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n646), .A2(KEYINPUT105), .A3(new_n653), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT105), .B1(new_n646), .B2(new_n653), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n727), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n717), .A2(new_n728), .A3(new_n718), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n735), .B1(new_n719), .B2(KEYINPUT108), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT53), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT54), .B1(new_n807), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n804), .B1(new_n815), .B2(new_n733), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT118), .B1(new_n816), .B2(new_n610), .ZN(new_n817));
  OR3_X1    g631(.A1(new_n791), .A2(new_n268), .A3(new_n664), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n724), .A2(new_n731), .A3(new_n732), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n732), .B1(new_n724), .B2(new_n731), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n803), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n822), .A3(new_n465), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n817), .A2(new_n818), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n800), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(G54));
  NAND3_X1  g640(.A1(new_n792), .A2(KEYINPUT58), .A3(G475), .ZN(new_n827));
  INV_X1    g641(.A(new_n371), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n829), .A2(new_n830), .A3(new_n800), .ZN(G60));
  NAND2_X1  g645(.A1(new_n543), .A2(new_n544), .ZN(new_n832));
  NAND2_X1  g646(.A1(G478), .A2(G902), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT59), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n832), .B1(new_n739), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n832), .A2(new_n834), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n815), .B2(new_n733), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n835), .A2(new_n837), .A3(new_n800), .ZN(G63));
  NAND2_X1  g652(.A1(G217), .A2(G902), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT60), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n724), .B2(new_n731), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n825), .B1(new_n841), .B2(new_n332), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n724), .A2(new_n731), .ZN(new_n843));
  INV_X1    g657(.A(new_n840), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n843), .A2(new_n571), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT120), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n323), .B1(new_n791), .B2(new_n840), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n841), .A2(new_n571), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n847), .A2(new_n848), .A3(new_n825), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT61), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n846), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n852), .B1(new_n846), .B2(new_n850), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(G66));
  AOI21_X1  g669(.A(new_n253), .B1(new_n415), .B2(G224), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n727), .A2(new_n703), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n856), .B1(new_n857), .B2(new_n253), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n794), .B1(G898), .B2(new_n253), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n858), .B(new_n859), .Z(G69));
  AOI21_X1  g674(.A(new_n253), .B1(G227), .B2(G900), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n239), .B(new_n361), .Z(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n658), .A2(new_n633), .A3(new_n710), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n680), .A2(new_n689), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n671), .A2(new_n711), .A3(new_n692), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n864), .A2(new_n660), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n253), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n587), .A2(G953), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT125), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT125), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n868), .A2(new_n872), .A3(new_n869), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n863), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n291), .A2(new_n335), .A3(new_n700), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n593), .A3(new_n679), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n605), .A2(new_n633), .A3(new_n710), .ZN(new_n877));
  AND2_X1   g691(.A1(KEYINPUT121), .A2(KEYINPUT62), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(KEYINPUT121), .A2(KEYINPUT62), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n877), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n865), .A2(new_n876), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n882), .A2(KEYINPUT122), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(KEYINPUT122), .ZN(new_n884));
  AOI21_X1  g698(.A(G953), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(new_n862), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n861), .B1(new_n874), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n873), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n872), .B1(new_n868), .B2(new_n869), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n862), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n891), .B1(new_n885), .B2(new_n862), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n886), .A2(KEYINPUT123), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n890), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n861), .B(KEYINPUT124), .Z(new_n895));
  OAI21_X1  g709(.A(new_n887), .B1(new_n894), .B2(new_n895), .ZN(G72));
  NAND2_X1  g710(.A1(G472), .A2(G902), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT63), .Z(new_n898));
  NAND2_X1  g712(.A1(new_n883), .A2(new_n884), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n898), .B1(new_n899), .B2(new_n857), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n596), .ZN(new_n901));
  INV_X1    g715(.A(new_n596), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n902), .A2(new_n262), .A3(new_n898), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT127), .Z(new_n904));
  NAND3_X1  g718(.A1(new_n734), .A2(new_n737), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n898), .B1(new_n867), .B2(new_n857), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n262), .B(KEYINPUT126), .Z(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AND4_X1   g722(.A1(new_n825), .A2(new_n901), .A3(new_n905), .A4(new_n908), .ZN(G57));
endmodule


