//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n585, new_n586, new_n587,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n604, new_n605, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n644,
    new_n645, new_n648, new_n650, new_n651, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1261;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT66), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT67), .B(G2105), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI211_X1 g042(.A(new_n460), .B(new_n461), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n467), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT67), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(KEYINPUT68), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n461), .A2(G137), .ZN(new_n477));
  INV_X1    g052(.A(new_n463), .ZN(new_n478));
  XNOR2_X1  g053(.A(KEYINPUT69), .B(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n464), .A2(KEYINPUT69), .ZN(new_n484));
  OAI211_X1 g059(.A(G101), .B(new_n470), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(KEYINPUT70), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n464), .A2(KEYINPUT69), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n482), .A2(G2104), .ZN(new_n489));
  AOI21_X1  g064(.A(G2105), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n487), .B1(new_n490), .B2(G101), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n481), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n476), .A2(new_n492), .ZN(G160));
  NAND2_X1  g068(.A1(new_n479), .A2(KEYINPUT3), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(new_n463), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n480), .A2(KEYINPUT71), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n461), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G124), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n480), .A2(KEYINPUT71), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n480), .A2(KEYINPUT71), .ZN(new_n502));
  OAI211_X1 g077(.A(G136), .B(new_n470), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(G100), .A2(G2105), .ZN(new_n504));
  XNOR2_X1  g079(.A(new_n504), .B(KEYINPUT72), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n505), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n500), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G162));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n471), .A2(new_n473), .A3(G138), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n463), .A2(new_n465), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g087(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n513));
  INV_X1    g088(.A(G114), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n513), .B1(new_n514), .B2(G2105), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT4), .A2(G138), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n461), .A2(new_n518), .B1(G126), .B2(G2105), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n512), .B(new_n516), .C1(new_n495), .C2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(G164));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n523));
  AND3_X1   g098(.A1(new_n523), .A2(KEYINPUT5), .A3(G543), .ZN(new_n524));
  AOI21_X1  g099(.A(G543), .B1(new_n523), .B2(KEYINPUT5), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G62), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n522), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  OAI21_X1  g105(.A(G543), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n528), .A2(G651), .B1(G50), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT6), .B(G651), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n534), .B1(new_n524), .B2(new_n525), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G543), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT5), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n539), .B2(KEYINPUT73), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n523), .A2(KEYINPUT5), .A3(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n542), .A2(KEYINPUT74), .A3(new_n534), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n537), .A2(G88), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n533), .A2(new_n544), .ZN(G303));
  INV_X1    g120(.A(G303), .ZN(G166));
  NAND3_X1  g121(.A1(new_n537), .A2(G89), .A3(new_n543), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n531), .A2(KEYINPUT75), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n549));
  OAI211_X1 g124(.A(new_n549), .B(G543), .C1(new_n529), .C2(new_n530), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G51), .ZN(new_n552));
  AND2_X1   g127(.A1(G63), .A2(G651), .ZN(new_n553));
  NAND3_X1  g128(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n554), .A2(KEYINPUT7), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(KEYINPUT7), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n542), .A2(new_n553), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AND3_X1   g132(.A1(new_n547), .A2(new_n552), .A3(new_n557), .ZN(G168));
  NAND3_X1  g133(.A1(new_n537), .A2(G90), .A3(new_n543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n551), .A2(G52), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(G64), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n540), .B2(new_n541), .ZN(new_n565));
  AND2_X1   g140(.A1(G77), .A2(G543), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g144(.A(KEYINPUT76), .B(G651), .C1(new_n565), .C2(new_n566), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n559), .A2(KEYINPUT77), .A3(new_n560), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n563), .A2(new_n571), .A3(new_n572), .ZN(G301));
  INV_X1    g148(.A(G301), .ZN(G171));
  NAND3_X1  g149(.A1(new_n537), .A2(G81), .A3(new_n543), .ZN(new_n575));
  NAND2_X1  g150(.A1(G68), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G56), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n526), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G651), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n551), .A2(G43), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n575), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G860), .ZN(G153));
  NAND4_X1  g158(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g159(.A1(G1), .A2(G3), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT8), .ZN(new_n586));
  NAND4_X1  g161(.A1(G319), .A2(G483), .A3(G661), .A4(new_n586), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT78), .ZN(G188));
  AND3_X1   g163(.A1(new_n542), .A2(KEYINPUT74), .A3(new_n534), .ZN(new_n589));
  AOI21_X1  g164(.A(KEYINPUT74), .B1(new_n542), .B2(new_n534), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT80), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT80), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n537), .A2(new_n592), .A3(new_n543), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n593), .A3(G91), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G53), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT9), .B1(new_n531), .B2(new_n596), .ZN(new_n597));
  OR3_X1    g172(.A1(new_n531), .A2(KEYINPUT9), .A3(new_n596), .ZN(new_n598));
  NAND2_X1  g173(.A1(G78), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G65), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n526), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n597), .A2(new_n598), .B1(new_n601), .B2(G651), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n594), .A2(new_n602), .ZN(G299));
  NAND2_X1  g178(.A1(new_n537), .A2(new_n543), .ZN(new_n604));
  INV_X1    g179(.A(G89), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n552), .B(new_n557), .C1(new_n604), .C2(new_n605), .ZN(G286));
  NAND3_X1  g181(.A1(new_n591), .A2(new_n593), .A3(G87), .ZN(new_n607));
  OAI21_X1  g182(.A(G651), .B1(new_n542), .B2(G74), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(KEYINPUT81), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n610), .B(G651), .C1(new_n542), .C2(G74), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n609), .A2(new_n611), .B1(G49), .B2(new_n532), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n607), .A2(new_n612), .ZN(G288));
  NAND3_X1  g188(.A1(new_n591), .A2(new_n593), .A3(G86), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n532), .A2(G48), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n542), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n616));
  INV_X1    g191(.A(G651), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n614), .A2(new_n619), .ZN(G305));
  NAND2_X1  g195(.A1(new_n551), .A2(G47), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n542), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT82), .B(G85), .Z(new_n623));
  OAI221_X1 g198(.A(new_n621), .B1(new_n617), .B2(new_n622), .C1(new_n604), .C2(new_n623), .ZN(G290));
  NAND2_X1  g199(.A1(G301), .A2(G868), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n591), .A2(new_n593), .A3(G92), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(KEYINPUT10), .ZN(new_n627));
  NAND2_X1  g202(.A1(G79), .A2(G543), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT84), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT85), .B(G66), .Z(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n526), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G651), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n548), .A2(KEYINPUT83), .A3(new_n550), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G54), .ZN(new_n634));
  AOI21_X1  g209(.A(KEYINPUT83), .B1(new_n548), .B2(new_n550), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT10), .ZN(new_n638));
  NAND4_X1  g213(.A1(new_n591), .A2(new_n593), .A3(new_n638), .A4(G92), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n627), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n625), .B1(new_n641), .B2(G868), .ZN(G284));
  OAI21_X1  g217(.A(new_n625), .B1(new_n641), .B2(G868), .ZN(G321));
  NAND2_X1  g218(.A1(G286), .A2(G868), .ZN(new_n644));
  AND2_X1   g219(.A1(new_n594), .A2(new_n602), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n644), .B1(new_n645), .B2(G868), .ZN(G297));
  OAI21_X1  g221(.A(new_n644), .B1(new_n645), .B2(G868), .ZN(G280));
  INV_X1    g222(.A(G559), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n641), .B1(new_n648), .B2(G860), .ZN(G148));
  NAND2_X1  g224(.A1(new_n641), .A2(new_n648), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(G868), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(G868), .B2(new_n582), .ZN(G323));
  XNOR2_X1  g227(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g228(.A1(new_n499), .A2(G123), .ZN(new_n654));
  OAI211_X1 g229(.A(G135), .B(new_n470), .C1(new_n501), .C2(new_n502), .ZN(new_n655));
  OAI221_X1 g230(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n461), .C2(G111), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n657), .A2(G2096), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(G2096), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT3), .B(G2104), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n490), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT13), .B(G2100), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n658), .A2(new_n659), .A3(new_n665), .ZN(G156));
  XOR2_X1   g241(.A(G2451), .B(G2454), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT16), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1341), .B(G1348), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT14), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2427), .B(G2438), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2430), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT15), .B(G2435), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n674), .B2(new_n673), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n670), .B(new_n676), .Z(new_n677));
  XNOR2_X1  g252(.A(G2443), .B(G2446), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n679), .A2(new_n680), .A3(G14), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT87), .Z(G401));
  XNOR2_X1  g257(.A(G2072), .B(G2078), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT17), .ZN(new_n684));
  XNOR2_X1  g259(.A(G2067), .B(G2678), .ZN(new_n685));
  XOR2_X1   g260(.A(G2084), .B(G2090), .Z(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n684), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT88), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n684), .A2(new_n685), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n690), .B(new_n687), .C1(new_n683), .C2(new_n685), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n686), .A2(new_n683), .A3(new_n685), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT18), .Z(new_n693));
  NAND3_X1  g268(.A1(new_n689), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(G2096), .Z(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT89), .B(G2100), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G227));
  XOR2_X1   g273(.A(G1971), .B(G1976), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT19), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1956), .B(G2474), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(G1961), .B(G1966), .Z(new_n703));
  AND2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT20), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n702), .A2(new_n703), .ZN(new_n707));
  NOR3_X1   g282(.A1(new_n700), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n700), .B2(new_n707), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(G1991), .B(G1996), .Z(new_n711));
  XOR2_X1   g286(.A(new_n710), .B(new_n711), .Z(new_n712));
  XOR2_X1   g287(.A(G1981), .B(G1986), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT90), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n712), .B(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(G229));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G26), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT28), .Z(new_n721));
  NAND2_X1  g296(.A1(new_n499), .A2(G128), .ZN(new_n722));
  OAI221_X1 g297(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n461), .C2(G116), .ZN(new_n723));
  INV_X1    g298(.A(G140), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n470), .B1(new_n501), .B2(new_n502), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n722), .B(new_n723), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n721), .B1(new_n726), .B2(G29), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G2067), .ZN(new_n728));
  INV_X1    g303(.A(G16), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G20), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT23), .Z(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G299), .B2(G16), .ZN(new_n732));
  INV_X1    g307(.A(G1956), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G19), .ZN(new_n735));
  OR3_X1    g310(.A1(new_n735), .A2(KEYINPUT96), .A3(G16), .ZN(new_n736));
  OAI21_X1  g311(.A(KEYINPUT96), .B1(new_n735), .B2(G16), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n736), .B(new_n737), .C1(new_n582), .C2(new_n729), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1341), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n734), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n500), .A2(G29), .A3(new_n503), .A4(new_n506), .ZN(new_n741));
  OR2_X1    g316(.A1(G29), .A2(G35), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(KEYINPUT29), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G2090), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n743), .A2(KEYINPUT29), .ZN(new_n747));
  AND3_X1   g322(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n746), .B1(new_n745), .B2(new_n747), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n728), .B(new_n740), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G4), .A2(G16), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT94), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n640), .B2(new_n729), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(KEYINPUT95), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(KEYINPUT95), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G1348), .ZN(new_n757));
  INV_X1    g332(.A(G1348), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n754), .A2(new_n758), .A3(new_n755), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n750), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  OAI211_X1 g335(.A(G139), .B(new_n470), .C1(new_n501), .C2(new_n502), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n762));
  NAND2_X1  g337(.A1(G103), .A2(G2104), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n474), .B2(new_n763), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n461), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n765));
  NAND2_X1  g340(.A1(G115), .A2(G2104), .ZN(new_n766));
  INV_X1    g341(.A(G127), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n511), .B2(new_n767), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n764), .A2(new_n765), .B1(new_n768), .B2(new_n474), .ZN(new_n769));
  AND3_X1   g344(.A1(new_n761), .A2(KEYINPUT97), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(KEYINPUT97), .B1(new_n761), .B2(new_n769), .ZN(new_n771));
  OAI21_X1  g346(.A(KEYINPUT98), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n761), .A2(new_n769), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT97), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT98), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n761), .A2(KEYINPUT97), .A3(new_n769), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n772), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G29), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n719), .A2(G33), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n780), .A2(G2072), .A3(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G2072), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n719), .B1(new_n772), .B2(new_n778), .ZN(new_n784));
  INV_X1    g359(.A(new_n781), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(G301), .A2(G16), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n729), .A2(G5), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(G1961), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n654), .A2(G29), .A3(new_n655), .A4(new_n656), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT30), .B(G28), .ZN(new_n793));
  OR2_X1    g368(.A1(KEYINPUT31), .A2(G11), .ZN(new_n794));
  NAND2_X1  g369(.A1(KEYINPUT31), .A2(G11), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n793), .A2(new_n719), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  OR3_X1    g372(.A1(G286), .A2(KEYINPUT102), .A3(new_n729), .ZN(new_n798));
  OR2_X1    g373(.A1(G16), .A2(G21), .ZN(new_n799));
  OAI211_X1 g374(.A(KEYINPUT102), .B(new_n799), .C1(G286), .C2(new_n729), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n797), .B1(new_n801), .B2(G1966), .ZN(new_n802));
  INV_X1    g377(.A(G1966), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n798), .A2(new_n803), .A3(new_n800), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n791), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT103), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g382(.A(G141), .B(new_n470), .C1(new_n501), .C2(new_n502), .ZN(new_n808));
  OAI211_X1 g383(.A(G129), .B(new_n474), .C1(new_n501), .C2(new_n502), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n490), .A2(G105), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(KEYINPUT99), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT99), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n490), .A2(new_n812), .A3(G105), .ZN(new_n813));
  NAND3_X1  g388(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n814), .A2(KEYINPUT100), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(KEYINPUT100), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(KEYINPUT26), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT26), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n815), .A2(new_n819), .A3(new_n816), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n811), .A2(new_n813), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n808), .A2(new_n809), .A3(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT101), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n823), .A2(new_n824), .A3(G29), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT27), .B(G1996), .Z(new_n826));
  OAI21_X1  g401(.A(new_n824), .B1(G29), .B2(G32), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n822), .B2(new_n719), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(G1961), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n788), .A2(new_n830), .A3(new_n789), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT104), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n719), .A2(G27), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n520), .B2(G29), .ZN(new_n835));
  INV_X1    g410(.A(G2078), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n835), .A2(new_n836), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n833), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n839), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n841), .A2(KEYINPUT104), .A3(new_n837), .ZN(new_n842));
  AND2_X1   g417(.A1(KEYINPUT24), .A2(G34), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n719), .B1(KEYINPUT24), .B2(G34), .ZN(new_n844));
  OAI22_X1  g419(.A1(G160), .A2(new_n719), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(G2084), .ZN(new_n846));
  INV_X1    g421(.A(G2084), .ZN(new_n847));
  OAI221_X1 g422(.A(new_n847), .B1(new_n843), .B2(new_n844), .C1(G160), .C2(new_n719), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n840), .A2(new_n842), .A3(new_n846), .A4(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n826), .B1(new_n825), .B2(new_n828), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n832), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n791), .A2(new_n802), .A3(KEYINPUT103), .A4(new_n804), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n787), .A2(new_n807), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT105), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n853), .A2(new_n854), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n760), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT106), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n853), .B(new_n854), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT106), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n860), .A3(new_n760), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n729), .A2(G6), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(G305), .B2(G16), .ZN(new_n863));
  XNOR2_X1  g438(.A(KEYINPUT32), .B(G1981), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n729), .A2(G23), .ZN(new_n866));
  XOR2_X1   g441(.A(KEYINPUT33), .B(G1976), .Z(new_n867));
  AOI211_X1 g442(.A(new_n866), .B(new_n867), .C1(G288), .C2(G16), .ZN(new_n868));
  NAND2_X1  g443(.A1(G303), .A2(G16), .ZN(new_n869));
  INV_X1    g444(.A(G1971), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n729), .A2(G22), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n870), .B1(new_n869), .B2(new_n871), .ZN(new_n873));
  NOR3_X1   g448(.A1(new_n868), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n607), .A2(new_n612), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n875), .A2(new_n729), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n867), .B1(new_n876), .B2(new_n866), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n865), .A2(new_n874), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT92), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT34), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT34), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n865), .A2(new_n874), .A3(new_n882), .A4(new_n877), .ZN(new_n883));
  XOR2_X1   g458(.A(KEYINPUT35), .B(G1991), .Z(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n499), .A2(G119), .ZN(new_n886));
  OAI211_X1 g461(.A(G131), .B(new_n470), .C1(new_n501), .C2(new_n502), .ZN(new_n887));
  OAI221_X1 g462(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n461), .C2(G107), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT91), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT91), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n886), .A2(new_n891), .A3(new_n887), .A4(new_n888), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n719), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n719), .A2(G25), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n885), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n890), .A2(new_n892), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n894), .B(new_n884), .C1(new_n897), .C2(new_n719), .ZN(new_n898));
  MUX2_X1   g473(.A(G24), .B(G290), .S(G16), .Z(new_n899));
  XOR2_X1   g474(.A(new_n899), .B(G1986), .Z(new_n900));
  NAND4_X1  g475(.A1(new_n883), .A2(new_n896), .A3(new_n898), .A4(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n879), .B1(new_n878), .B2(KEYINPUT34), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n881), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT93), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT36), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AND4_X1   g480(.A1(new_n883), .A2(new_n896), .A3(new_n898), .A4(new_n900), .ZN(new_n906));
  INV_X1    g481(.A(new_n902), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n907), .A3(new_n880), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT36), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(KEYINPUT93), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n903), .A2(new_n904), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n858), .A2(new_n861), .B1(new_n911), .B2(new_n912), .ZN(G311));
  NOR3_X1   g488(.A1(new_n903), .A2(new_n904), .A3(KEYINPUT36), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n909), .B1(new_n908), .B2(KEYINPUT93), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n857), .A2(KEYINPUT106), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n860), .B1(new_n859), .B2(new_n760), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(G150));
  NOR2_X1   g494(.A1(new_n640), .A2(new_n648), .ZN(new_n920));
  XNOR2_X1  g495(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n920), .B(new_n921), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n578), .A2(G651), .B1(new_n551), .B2(G43), .ZN(new_n923));
  NAND2_X1  g498(.A1(G80), .A2(G543), .ZN(new_n924));
  INV_X1    g499(.A(G67), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n924), .B1(new_n526), .B2(new_n925), .ZN(new_n926));
  AOI22_X1  g501(.A1(new_n926), .A2(G651), .B1(new_n551), .B2(G55), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n537), .A2(G93), .A3(new_n543), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n923), .A2(new_n927), .A3(new_n575), .A4(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n926), .A2(G651), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n551), .A2(G55), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n581), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n922), .B(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n935), .A2(KEYINPUT39), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(KEYINPUT108), .ZN(new_n937));
  AOI21_X1  g512(.A(G860), .B1(new_n935), .B2(KEYINPUT39), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n932), .A2(G860), .ZN(new_n940));
  XOR2_X1   g515(.A(new_n940), .B(KEYINPUT37), .Z(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(G145));
  XOR2_X1   g517(.A(new_n889), .B(KEYINPUT109), .Z(new_n943));
  NAND2_X1  g518(.A1(new_n499), .A2(G130), .ZN(new_n944));
  OAI221_X1 g519(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n461), .C2(G118), .ZN(new_n945));
  INV_X1    g520(.A(G142), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n944), .B(new_n945), .C1(new_n946), .C2(new_n725), .ZN(new_n947));
  INV_X1    g522(.A(new_n663), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n943), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n949), .A2(new_n950), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n889), .B(KEYINPUT109), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n726), .A2(G164), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n725), .A2(new_n724), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n957), .A2(new_n520), .A3(new_n722), .A4(new_n723), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n823), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n956), .A2(new_n823), .A3(new_n958), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n779), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n961), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n770), .A2(new_n771), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n963), .A2(new_n959), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n955), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n772), .B(new_n778), .C1(new_n963), .C2(new_n959), .ZN(new_n967));
  INV_X1    g542(.A(new_n964), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n960), .A2(new_n968), .A3(new_n961), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n967), .A2(new_n969), .A3(new_n951), .A4(new_n954), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n966), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  XOR2_X1   g547(.A(new_n507), .B(new_n657), .Z(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(G160), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G37), .ZN(new_n976));
  INV_X1    g551(.A(new_n974), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n966), .A2(new_n970), .A3(new_n977), .A4(new_n971), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g555(.A1(new_n929), .A2(new_n933), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n650), .B(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n640), .A2(G299), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n636), .B1(KEYINPUT10), .B2(new_n626), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n984), .A2(new_n645), .A3(new_n639), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n982), .A2(new_n986), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n983), .A2(new_n985), .A3(KEYINPUT41), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT41), .B1(new_n983), .B2(new_n985), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n987), .B1(new_n982), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g566(.A(KEYINPUT111), .B(KEYINPUT42), .Z(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(G288), .B(G303), .ZN(new_n994));
  XNOR2_X1  g569(.A(G305), .B(G290), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n994), .B(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n992), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n987), .B(new_n998), .C1(new_n982), .C2(new_n990), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n993), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n997), .B1(new_n993), .B2(new_n999), .ZN(new_n1001));
  OAI21_X1  g576(.A(G868), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n932), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1002), .B1(G868), .B2(new_n1003), .ZN(G295));
  OAI21_X1  g579(.A(new_n1002), .B1(G868), .B2(new_n1003), .ZN(G331));
  NAND2_X1  g580(.A1(new_n572), .A2(new_n571), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT77), .B1(new_n559), .B2(new_n560), .ZN(new_n1007));
  OAI21_X1  g582(.A(G286), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n563), .A2(G168), .A3(new_n571), .A4(new_n572), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n981), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n934), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT41), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n640), .A2(G299), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n645), .B1(new_n984), .B2(new_n639), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n983), .A2(new_n985), .A3(KEYINPUT41), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1013), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1012), .A2(KEYINPUT112), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n934), .A2(new_n1022), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1020), .A2(new_n1021), .A3(new_n1011), .A4(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1019), .A2(new_n1024), .A3(new_n996), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1027));
  AOI21_X1  g602(.A(G37), .B1(new_n1027), .B2(new_n997), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1026), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n996), .B1(new_n1019), .B2(new_n1024), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT113), .B1(new_n1031), .B2(G37), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT43), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1020), .A2(new_n1011), .A3(new_n1023), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n990), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n934), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(new_n986), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1037), .A2(new_n1012), .ZN(new_n1038));
  OAI211_X1 g613(.A(KEYINPUT114), .B(new_n997), .C1(new_n1035), .C2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n990), .A2(new_n1034), .B1(new_n1012), .B2(new_n1037), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(new_n996), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1025), .A2(new_n976), .ZN(new_n1043));
  AND4_X1   g618(.A1(KEYINPUT43), .A2(new_n1039), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT44), .B1(new_n1033), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT44), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT43), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1048));
  AND4_X1   g623(.A1(new_n1047), .A2(new_n1039), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1046), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1045), .A2(new_n1050), .ZN(G397));
  INV_X1    g626(.A(G8), .ZN(new_n1052));
  INV_X1    g627(.A(new_n467), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1053), .B1(new_n660), .B2(G125), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n460), .B1(new_n1054), .B2(new_n461), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n469), .A2(KEYINPUT68), .A3(new_n474), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n485), .A2(KEYINPUT70), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n490), .A2(new_n487), .A3(G101), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1058), .A2(new_n1059), .B1(new_n480), .B2(new_n477), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1057), .A2(new_n1060), .A3(G40), .ZN(new_n1061));
  INV_X1    g636(.A(G1384), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n520), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT45), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1061), .A2(new_n1065), .A3(KEYINPUT118), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1057), .A2(new_n1060), .A3(G40), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT45), .B1(new_n520), .B2(new_n1062), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G126), .A2(G2105), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n474), .B2(new_n517), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n515), .B1(new_n1072), .B2(new_n480), .ZN(new_n1073));
  AOI21_X1  g648(.A(G1384), .B1(new_n1073), .B2(new_n512), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT45), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1066), .A2(new_n1070), .A3(new_n1075), .ZN(new_n1076));
  AOI211_X1 g651(.A(KEYINPUT50), .B(G1384), .C1(new_n1073), .C2(new_n512), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT50), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1078), .B1(new_n520), .B2(new_n1062), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n1077), .A2(new_n1068), .A3(new_n1079), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1076), .A2(new_n803), .B1(new_n847), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1052), .B1(new_n1081), .B2(G168), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT51), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1076), .A2(new_n803), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1080), .A2(new_n847), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(G286), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1083), .B1(new_n1082), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT62), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(G8), .B1(new_n1088), .B2(G286), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1081), .A2(G168), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT51), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT62), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1094), .A2(new_n1095), .A3(new_n1084), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT55), .ZN(new_n1098));
  AOI211_X1 g673(.A(new_n1098), .B(new_n1052), .C1(new_n533), .C2(new_n544), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1061), .A2(new_n1065), .A3(new_n1075), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1080), .A2(new_n746), .B1(new_n1101), .B2(new_n870), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1100), .B1(new_n1102), .B2(new_n1052), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1061), .A2(new_n1065), .A3(new_n1075), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1079), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1074), .A2(new_n1078), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n1061), .A3(new_n1106), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n1104), .A2(G1971), .B1(new_n1107), .B2(G2090), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1100), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(new_n1109), .A3(G8), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1103), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n875), .A2(G1976), .ZN(new_n1112));
  INV_X1    g687(.A(G1976), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT52), .B1(G288), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(G8), .B1(new_n1068), .B2(new_n1063), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1112), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(G288), .A2(new_n1113), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT52), .B1(new_n1118), .B2(new_n1115), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G1981), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n614), .A2(new_n1121), .A3(new_n619), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n537), .A2(G86), .A3(new_n543), .ZN(new_n1123));
  OAI21_X1  g698(.A(G1981), .B1(new_n1123), .B2(new_n618), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT49), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT116), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1115), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT116), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1122), .A2(new_n1124), .A3(new_n1129), .A4(KEYINPUT49), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1127), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1120), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1133), .B1(new_n1101), .B2(G2078), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT126), .B(G1961), .Z(new_n1135));
  NAND2_X1  g710(.A1(new_n1107), .A2(new_n1135), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1133), .A2(G2078), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1066), .A2(new_n1070), .A3(new_n1075), .A4(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(G301), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1111), .A2(new_n1132), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1091), .A2(new_n1096), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT117), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1122), .ZN(new_n1144));
  NOR2_X1   g719(.A1(G288), .A2(G1976), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1144), .B1(new_n1131), .B2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1146), .A2(new_n1115), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1102), .A2(new_n1052), .A3(new_n1100), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1148), .A2(new_n1131), .A3(new_n1120), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1143), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1148), .A2(new_n1131), .A3(new_n1120), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1151), .B(KEYINPUT117), .C1(new_n1115), .C2(new_n1146), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT119), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1153), .A2(KEYINPUT63), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1103), .A2(new_n1120), .A3(new_n1110), .A4(new_n1131), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1088), .A2(G8), .A3(G168), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1154), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1081), .A2(new_n1052), .A3(G286), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1111), .A2(new_n1132), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  AOI22_X1  g735(.A1(new_n1150), .A2(new_n1152), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(KEYINPUT56), .B(G2072), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1061), .A2(new_n1065), .A3(new_n1075), .A4(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1163), .B1(new_n1080), .B2(G1956), .ZN(new_n1164));
  NAND2_X1  g739(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT57), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n594), .A2(new_n1166), .A3(new_n602), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1168), .A2(KEYINPUT121), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1170), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1164), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1164), .A2(new_n1168), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n641), .ZN(new_n1174));
  NAND4_X1  g749(.A1(G160), .A2(KEYINPUT120), .A3(G40), .A4(new_n1074), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT120), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1176), .B1(new_n1068), .B2(new_n1063), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(G2067), .ZN(new_n1179));
  AOI22_X1  g754(.A1(new_n1178), .A2(new_n1179), .B1(new_n758), .B2(new_n1107), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1172), .B1(new_n1174), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT59), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1182), .A2(KEYINPUT123), .ZN(new_n1183));
  XOR2_X1   g758(.A(KEYINPUT58), .B(G1341), .Z(new_n1184));
  NAND3_X1  g759(.A1(new_n1175), .A2(new_n1177), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT122), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1175), .A2(new_n1177), .A3(KEYINPUT122), .A4(new_n1184), .ZN(new_n1188));
  INV_X1    g763(.A(G1996), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1061), .A2(new_n1065), .A3(new_n1075), .A4(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n582), .B(new_n1183), .C1(new_n1187), .C2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n582), .B1(new_n1187), .B2(new_n1191), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1183), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1172), .A2(new_n1173), .A3(KEYINPUT61), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT61), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT124), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1164), .A2(new_n1198), .A3(new_n1168), .ZN(new_n1199));
  OAI21_X1  g774(.A(KEYINPUT124), .B1(new_n1164), .B2(new_n1168), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1107), .A2(new_n733), .ZN(new_n1201));
  AOI22_X1  g776(.A1(new_n1201), .A2(new_n1163), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1202));
  OAI211_X1 g777(.A(new_n1197), .B(new_n1199), .C1(new_n1200), .C2(new_n1202), .ZN(new_n1203));
  AND4_X1   g778(.A1(new_n1192), .A2(new_n1195), .A3(new_n1196), .A4(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n641), .B1(new_n1180), .B2(KEYINPUT60), .ZN(new_n1205));
  INV_X1    g780(.A(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT125), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1180), .A2(new_n1207), .A3(KEYINPUT60), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1207), .B1(new_n1180), .B2(KEYINPUT60), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1206), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1210), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1212), .A2(new_n1205), .A3(new_n1208), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1181), .B1(new_n1204), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1137), .A2(G301), .A3(new_n1139), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT54), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT115), .ZN(new_n1218));
  AOI21_X1  g793(.A(KEYINPUT45), .B1(new_n1063), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1219), .B1(new_n1218), .B2(new_n1063), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1138), .A2(G40), .ZN(new_n1221));
  AOI211_X1 g796(.A(new_n1221), .B(new_n492), .C1(new_n474), .C2(new_n469), .ZN(new_n1222));
  NAND3_X1  g797(.A1(new_n1220), .A2(new_n1075), .A3(new_n1222), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1223), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1217), .B1(new_n1224), .B2(G171), .ZN(new_n1225));
  AOI21_X1  g800(.A(new_n1155), .B1(new_n1216), .B2(new_n1225), .ZN(new_n1226));
  NOR2_X1   g801(.A1(new_n1224), .A2(G171), .ZN(new_n1227));
  OAI21_X1  g802(.A(new_n1217), .B1(new_n1140), .B2(new_n1227), .ZN(new_n1228));
  OAI211_X1 g803(.A(new_n1226), .B(new_n1228), .C1(new_n1090), .C2(new_n1085), .ZN(new_n1229));
  OAI211_X1 g804(.A(new_n1142), .B(new_n1161), .C1(new_n1215), .C2(new_n1229), .ZN(new_n1230));
  XNOR2_X1  g805(.A(new_n726), .B(new_n1179), .ZN(new_n1231));
  XNOR2_X1  g806(.A(new_n822), .B(new_n1189), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NOR2_X1   g808(.A1(new_n1220), .A2(new_n1068), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  XNOR2_X1  g810(.A(new_n889), .B(new_n885), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1236), .A2(new_n1234), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  XNOR2_X1  g813(.A(G290), .B(G1986), .ZN(new_n1239));
  AOI21_X1  g814(.A(new_n1238), .B1(new_n1234), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1230), .A2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g816(.A1(new_n1235), .A2(new_n897), .A3(new_n884), .ZN(new_n1242));
  OR2_X1    g817(.A1(new_n726), .A2(G2067), .ZN(new_n1243));
  NAND3_X1  g818(.A1(new_n1242), .A2(KEYINPUT127), .A3(new_n1243), .ZN(new_n1244));
  NAND2_X1  g819(.A1(new_n1244), .A2(new_n1234), .ZN(new_n1245));
  AOI21_X1  g820(.A(KEYINPUT127), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1246));
  NOR2_X1   g821(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g822(.A1(new_n1234), .A2(new_n1189), .ZN(new_n1248));
  OR2_X1    g823(.A1(new_n1248), .A2(KEYINPUT46), .ZN(new_n1249));
  NAND2_X1  g824(.A1(new_n1248), .A2(KEYINPUT46), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1231), .A2(new_n823), .ZN(new_n1251));
  AOI22_X1  g826(.A1(new_n1249), .A2(new_n1250), .B1(new_n1251), .B2(new_n1234), .ZN(new_n1252));
  XNOR2_X1  g827(.A(new_n1252), .B(KEYINPUT47), .ZN(new_n1253));
  NOR2_X1   g828(.A1(G290), .A2(G1986), .ZN(new_n1254));
  NAND2_X1  g829(.A1(new_n1234), .A2(new_n1254), .ZN(new_n1255));
  XOR2_X1   g830(.A(new_n1255), .B(KEYINPUT48), .Z(new_n1256));
  NOR2_X1   g831(.A1(new_n1256), .A2(new_n1238), .ZN(new_n1257));
  NOR3_X1   g832(.A1(new_n1247), .A2(new_n1253), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g833(.A1(new_n1241), .A2(new_n1258), .ZN(G329));
  assign    G231 = 1'b0;
  AND4_X1   g834(.A1(G319), .A2(new_n697), .A3(new_n681), .A4(new_n717), .ZN(new_n1261));
  OAI211_X1 g835(.A(new_n979), .B(new_n1261), .C1(new_n1048), .C2(new_n1049), .ZN(G225));
  INV_X1    g836(.A(G225), .ZN(G308));
endmodule


