

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744;

  INV_X1 U369 ( .A(n610), .ZN(n718) );
  XNOR2_X1 U370 ( .A(n374), .B(n606), .ZN(n610) );
  NAND2_X1 U371 ( .A1(n376), .A2(n375), .ZN(n374) );
  XNOR2_X1 U372 ( .A(n580), .B(n579), .ZN(n647) );
  AND2_X1 U373 ( .A1(n523), .A2(n667), .ZN(n560) );
  BUF_X1 U374 ( .A(n578), .Z(n491) );
  AND2_X1 U375 ( .A1(n521), .A2(n520), .ZN(n544) );
  XNOR2_X1 U376 ( .A(n561), .B(KEYINPUT19), .ZN(n379) );
  NAND2_X1 U377 ( .A1(n497), .A2(n687), .ZN(n561) );
  OR2_X1 U378 ( .A1(n622), .A2(n406), .ZN(n411) );
  XNOR2_X1 U379 ( .A(n353), .B(n464), .ZN(n714) );
  XNOR2_X1 U380 ( .A(G101), .B(G140), .ZN(n474) );
  INV_X1 U381 ( .A(G953), .ZN(n419) );
  AND2_X2 U382 ( .A1(n491), .A2(n490), .ZN(n581) );
  XNOR2_X1 U383 ( .A(n732), .B(n349), .ZN(n631) );
  XNOR2_X1 U384 ( .A(n475), .B(n476), .ZN(n349) );
  XNOR2_X1 U385 ( .A(n498), .B(KEYINPUT39), .ZN(n530) );
  NAND2_X1 U386 ( .A1(n550), .A2(n688), .ZN(n498) );
  XNOR2_X2 U387 ( .A(KEYINPUT18), .B(G125), .ZN(n388) );
  NOR2_X2 U388 ( .A1(n494), .A2(n677), .ZN(n495) );
  XNOR2_X2 U389 ( .A(n552), .B(KEYINPUT85), .ZN(n559) );
  XNOR2_X2 U390 ( .A(n471), .B(n470), .ZN(n359) );
  XNOR2_X2 U391 ( .A(n396), .B(n395), .ZN(n723) );
  XNOR2_X2 U392 ( .A(G110), .B(G107), .ZN(n396) );
  XNOR2_X1 U393 ( .A(n566), .B(n565), .ZN(n742) );
  NOR2_X2 U394 ( .A1(n373), .A2(n383), .ZN(n612) );
  AND2_X1 U395 ( .A1(n363), .A2(n406), .ZN(n381) );
  NOR2_X1 U396 ( .A1(n567), .A2(n742), .ZN(n568) );
  XNOR2_X1 U397 ( .A(n411), .B(n410), .ZN(n497) );
  XNOR2_X2 U398 ( .A(G125), .B(G140), .ZN(n438) );
  NOR2_X1 U399 ( .A1(n631), .A2(G902), .ZN(n351) );
  BUF_X1 U400 ( .A(n649), .Z(n350) );
  XNOR2_X1 U401 ( .A(n532), .B(n531), .ZN(n649) );
  XNOR2_X2 U402 ( .A(n351), .B(n352), .ZN(n589) );
  XOR2_X1 U403 ( .A(n479), .B(n478), .Z(n352) );
  OR2_X1 U404 ( .A1(n656), .A2(n671), .ZN(n365) );
  XNOR2_X1 U405 ( .A(G116), .B(G113), .ZN(n399) );
  NAND2_X1 U406 ( .A1(n688), .A2(n687), .ZN(n691) );
  XNOR2_X1 U407 ( .A(G902), .B(KEYINPUT95), .ZN(n405) );
  XOR2_X1 U408 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n606) );
  AND2_X1 U409 ( .A1(n354), .A2(n377), .ZN(n376) );
  INV_X1 U410 ( .A(KEYINPUT30), .ZN(n357) );
  XNOR2_X1 U411 ( .A(n418), .B(KEYINPUT0), .ZN(n506) );
  XNOR2_X1 U412 ( .A(n446), .B(n445), .ZN(n519) );
  BUF_X1 U413 ( .A(n506), .Z(n592) );
  NAND2_X1 U414 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U415 ( .A(n365), .B(n593), .ZN(n596) );
  INV_X1 U416 ( .A(G237), .ZN(n407) );
  XNOR2_X1 U417 ( .A(G101), .B(KEYINPUT73), .ZN(n398) );
  XNOR2_X1 U418 ( .A(n421), .B(n420), .ZN(n453) );
  XNOR2_X1 U419 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n420) );
  NAND2_X1 U420 ( .A1(n406), .A2(KEYINPUT2), .ZN(n382) );
  NAND2_X1 U421 ( .A1(n381), .A2(n718), .ZN(n380) );
  INV_X1 U422 ( .A(n687), .ZN(n370) );
  INV_X1 U423 ( .A(n533), .ZN(n688) );
  BUF_X1 U424 ( .A(n497), .Z(n528) );
  INV_X1 U425 ( .A(G902), .ZN(n444) );
  XNOR2_X1 U426 ( .A(G137), .B(G146), .ZN(n461) );
  XOR2_X1 U427 ( .A(G107), .B(KEYINPUT9), .Z(n423) );
  NAND2_X1 U428 ( .A1(G234), .A2(G237), .ZN(n413) );
  NAND2_X1 U429 ( .A1(n718), .A2(n611), .ZN(n373) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n706) );
  INV_X1 U431 ( .A(KEYINPUT41), .ZN(n371) );
  NAND2_X1 U432 ( .A1(n688), .A2(n369), .ZN(n372) );
  NOR2_X1 U433 ( .A1(n690), .A2(n370), .ZN(n369) );
  XNOR2_X1 U434 ( .A(n496), .B(n357), .ZN(n356) );
  XNOR2_X1 U435 ( .A(n631), .B(n634), .ZN(n635) );
  AND2_X1 U436 ( .A1(n618), .A2(G953), .ZN(n717) );
  XNOR2_X1 U437 ( .A(n373), .B(KEYINPUT2), .ZN(n710) );
  XNOR2_X1 U438 ( .A(n367), .B(n366), .ZN(n671) );
  INV_X1 U439 ( .A(KEYINPUT31), .ZN(n366) );
  NOR2_X1 U440 ( .A1(n592), .A2(n682), .ZN(n367) );
  XNOR2_X1 U441 ( .A(n368), .B(KEYINPUT100), .ZN(n656) );
  NOR2_X1 U442 ( .A1(n592), .A2(n591), .ZN(n368) );
  XNOR2_X1 U443 ( .A(n528), .B(KEYINPUT38), .ZN(n533) );
  BUF_X1 U444 ( .A(n419), .Z(n738) );
  XOR2_X1 U445 ( .A(n454), .B(n731), .Z(n353) );
  AND2_X1 U446 ( .A1(n598), .A2(n597), .ZN(n354) );
  INV_X1 U447 ( .A(KEYINPUT2), .ZN(n383) );
  XNOR2_X2 U448 ( .A(n355), .B(KEYINPUT81), .ZN(n550) );
  NAND2_X1 U449 ( .A1(n358), .A2(n356), .ZN(n355) );
  XNOR2_X1 U450 ( .A(n495), .B(KEYINPUT82), .ZN(n358) );
  XNOR2_X2 U451 ( .A(n472), .B(n359), .ZN(n732) );
  XNOR2_X2 U452 ( .A(n361), .B(n360), .ZN(n471) );
  XNOR2_X2 U453 ( .A(KEYINPUT68), .B(KEYINPUT69), .ZN(n360) );
  XNOR2_X2 U454 ( .A(G146), .B(G131), .ZN(n361) );
  XNOR2_X2 U455 ( .A(n425), .B(G134), .ZN(n472) );
  XNOR2_X2 U456 ( .A(n362), .B(n392), .ZN(n425) );
  XNOR2_X2 U457 ( .A(G143), .B(KEYINPUT84), .ZN(n362) );
  XNOR2_X1 U458 ( .A(n609), .B(KEYINPUT79), .ZN(n363) );
  NAND2_X1 U459 ( .A1(n364), .A2(n574), .ZN(n609) );
  XNOR2_X1 U460 ( .A(n571), .B(n570), .ZN(n364) );
  XNOR2_X2 U461 ( .A(n430), .B(n429), .ZN(n520) );
  NOR2_X2 U462 ( .A1(n637), .A2(n717), .ZN(n639) );
  NOR2_X2 U463 ( .A1(n643), .A2(n717), .ZN(n646) );
  NOR2_X2 U464 ( .A1(n619), .A2(n717), .ZN(n621) );
  NOR2_X2 U465 ( .A1(n628), .A2(n717), .ZN(n630) );
  XNOR2_X2 U466 ( .A(n608), .B(KEYINPUT65), .ZN(n613) );
  NAND2_X1 U467 ( .A1(n378), .A2(n605), .ZN(n375) );
  NAND2_X1 U468 ( .A1(n585), .A2(KEYINPUT44), .ZN(n377) );
  NAND2_X1 U469 ( .A1(n603), .A2(n604), .ZN(n378) );
  NAND2_X1 U470 ( .A1(n379), .A2(n386), .ZN(n418) );
  AND2_X1 U471 ( .A1(n379), .A2(n540), .ZN(n541) );
  NAND2_X1 U472 ( .A1(n380), .A2(n382), .ZN(n608) );
  BUF_X1 U473 ( .A(n650), .Z(n713) );
  XOR2_X1 U474 ( .A(KEYINPUT77), .B(KEYINPUT22), .Z(n384) );
  AND2_X1 U475 ( .A1(n493), .A2(n492), .ZN(n385) );
  AND2_X1 U476 ( .A1(n493), .A2(n417), .ZN(n386) );
  INV_X1 U477 ( .A(n581), .ZN(n582) );
  INV_X1 U478 ( .A(KEYINPUT102), .ZN(n433) );
  AND2_X1 U479 ( .A1(n673), .A2(n385), .ZN(n515) );
  XNOR2_X1 U480 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U481 ( .A(n436), .B(n435), .ZN(n439) );
  INV_X1 U482 ( .A(KEYINPUT10), .ZN(n437) );
  XNOR2_X1 U483 ( .A(n640), .B(KEYINPUT62), .ZN(n641) );
  BUF_X1 U484 ( .A(n647), .Z(n648) );
  XNOR2_X2 U485 ( .A(G146), .B(KEYINPUT17), .ZN(n387) );
  XNOR2_X1 U486 ( .A(n388), .B(n387), .ZN(n391) );
  NAND2_X1 U487 ( .A1(n419), .A2(G224), .ZN(n389) );
  XNOR2_X1 U488 ( .A(n389), .B(KEYINPUT4), .ZN(n390) );
  XNOR2_X1 U489 ( .A(n391), .B(n390), .ZN(n394) );
  INV_X1 U490 ( .A(G128), .ZN(n392) );
  INV_X1 U491 ( .A(n425), .ZN(n393) );
  XNOR2_X1 U492 ( .A(n394), .B(n393), .ZN(n397) );
  INV_X1 U493 ( .A(G104), .ZN(n395) );
  XNOR2_X1 U494 ( .A(n723), .B(KEYINPUT74), .ZN(n476) );
  XNOR2_X1 U495 ( .A(n397), .B(n476), .ZN(n403) );
  XNOR2_X1 U496 ( .A(n399), .B(n398), .ZN(n401) );
  XNOR2_X1 U497 ( .A(KEYINPUT3), .B(G119), .ZN(n400) );
  XNOR2_X1 U498 ( .A(n401), .B(n400), .ZN(n484) );
  XNOR2_X1 U499 ( .A(KEYINPUT16), .B(G122), .ZN(n402) );
  XNOR2_X1 U500 ( .A(n484), .B(n402), .ZN(n726) );
  XNOR2_X1 U501 ( .A(n403), .B(n726), .ZN(n622) );
  INV_X1 U502 ( .A(KEYINPUT15), .ZN(n404) );
  XNOR2_X1 U503 ( .A(n405), .B(n404), .ZN(n607) );
  INV_X1 U504 ( .A(n607), .ZN(n406) );
  NAND2_X1 U505 ( .A1(n407), .A2(n444), .ZN(n412) );
  NAND2_X1 U506 ( .A1(n412), .A2(G210), .ZN(n409) );
  XNOR2_X1 U507 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n408) );
  XNOR2_X1 U508 ( .A(n409), .B(n408), .ZN(n410) );
  NAND2_X1 U509 ( .A1(n412), .A2(G214), .ZN(n687) );
  XNOR2_X1 U510 ( .A(n413), .B(KEYINPUT14), .ZN(n701) );
  INV_X1 U511 ( .A(G952), .ZN(n618) );
  NAND2_X1 U512 ( .A1(n738), .A2(n618), .ZN(n415) );
  OR2_X1 U513 ( .A1(n738), .A2(G902), .ZN(n414) );
  AND2_X1 U514 ( .A1(n415), .A2(n414), .ZN(n416) );
  AND2_X1 U515 ( .A1(n701), .A2(n416), .ZN(n493) );
  NAND2_X1 U516 ( .A1(G953), .A2(G898), .ZN(n417) );
  NAND2_X1 U517 ( .A1(n419), .A2(G234), .ZN(n421) );
  NAND2_X1 U518 ( .A1(G217), .A2(n453), .ZN(n422) );
  XNOR2_X1 U519 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U520 ( .A(n424), .B(KEYINPUT7), .ZN(n428) );
  XNOR2_X1 U521 ( .A(G116), .B(G122), .ZN(n426) );
  XOR2_X1 U522 ( .A(n472), .B(n426), .Z(n427) );
  XNOR2_X1 U523 ( .A(n427), .B(n428), .ZN(n651) );
  NAND2_X1 U524 ( .A1(n651), .A2(n444), .ZN(n430) );
  INV_X1 U525 ( .A(G478), .ZN(n429) );
  XOR2_X1 U526 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n432) );
  XNOR2_X1 U527 ( .A(G143), .B(G104), .ZN(n431) );
  XNOR2_X1 U528 ( .A(n432), .B(n431), .ZN(n436) );
  XNOR2_X1 U529 ( .A(G113), .B(G122), .ZN(n434) );
  XNOR2_X2 U530 ( .A(n438), .B(n437), .ZN(n731) );
  XNOR2_X1 U531 ( .A(n439), .B(n731), .ZN(n443) );
  NOR2_X2 U532 ( .A1(G237), .A2(G953), .ZN(n440) );
  XNOR2_X1 U533 ( .A(KEYINPUT80), .B(n440), .ZN(n480) );
  NAND2_X1 U534 ( .A1(n480), .A2(G214), .ZN(n441) );
  XNOR2_X1 U535 ( .A(n471), .B(n441), .ZN(n442) );
  XNOR2_X1 U536 ( .A(n443), .B(n442), .ZN(n615) );
  NAND2_X1 U537 ( .A1(n615), .A2(n444), .ZN(n446) );
  XNOR2_X1 U538 ( .A(KEYINPUT13), .B(G475), .ZN(n445) );
  NAND2_X1 U539 ( .A1(n520), .A2(n519), .ZN(n690) );
  NAND2_X1 U540 ( .A1(G234), .A2(n607), .ZN(n447) );
  XNOR2_X1 U541 ( .A(KEYINPUT20), .B(n447), .ZN(n465) );
  AND2_X1 U542 ( .A1(n465), .A2(G221), .ZN(n449) );
  XNOR2_X1 U543 ( .A(KEYINPUT98), .B(KEYINPUT21), .ZN(n448) );
  XNOR2_X1 U544 ( .A(n449), .B(n448), .ZN(n673) );
  INV_X1 U545 ( .A(n673), .ZN(n450) );
  OR2_X1 U546 ( .A1(n690), .A2(n450), .ZN(n451) );
  NOR2_X2 U547 ( .A1(n506), .A2(n451), .ZN(n452) );
  XNOR2_X1 U548 ( .A(n452), .B(n384), .ZN(n578) );
  NAND2_X1 U549 ( .A1(G221), .A2(n453), .ZN(n454) );
  XNOR2_X1 U550 ( .A(G119), .B(G128), .ZN(n460) );
  INV_X1 U551 ( .A(G110), .ZN(n455) );
  NAND2_X1 U552 ( .A1(KEYINPUT23), .A2(n455), .ZN(n458) );
  INV_X1 U553 ( .A(KEYINPUT23), .ZN(n456) );
  NAND2_X1 U554 ( .A1(n456), .A2(G110), .ZN(n457) );
  NAND2_X1 U555 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X1 U556 ( .A(n460), .B(n459), .ZN(n463) );
  XNOR2_X1 U557 ( .A(n461), .B(KEYINPUT24), .ZN(n462) );
  XOR2_X1 U558 ( .A(n463), .B(n462), .Z(n464) );
  NOR2_X2 U559 ( .A1(n714), .A2(G902), .ZN(n468) );
  NAND2_X1 U560 ( .A1(n465), .A2(G217), .ZN(n466) );
  XNOR2_X1 U561 ( .A(KEYINPUT25), .B(n466), .ZN(n467) );
  XNOR2_X2 U562 ( .A(n468), .B(n467), .ZN(n514) );
  INV_X1 U563 ( .A(KEYINPUT103), .ZN(n469) );
  XNOR2_X1 U564 ( .A(n514), .B(n469), .ZN(n674) );
  XNOR2_X1 U565 ( .A(KEYINPUT4), .B(G137), .ZN(n470) );
  NAND2_X1 U566 ( .A1(n738), .A2(G227), .ZN(n473) );
  XNOR2_X1 U567 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U568 ( .A(KEYINPUT72), .B(G469), .ZN(n479) );
  INV_X1 U569 ( .A(KEYINPUT71), .ZN(n478) );
  XNOR2_X1 U570 ( .A(n589), .B(KEYINPUT1), .ZN(n587) );
  INV_X1 U571 ( .A(n587), .ZN(n678) );
  NAND2_X1 U572 ( .A1(n674), .A2(n678), .ZN(n487) );
  NAND2_X1 U573 ( .A1(n480), .A2(G210), .ZN(n482) );
  XNOR2_X1 U574 ( .A(KEYINPUT99), .B(KEYINPUT5), .ZN(n481) );
  XNOR2_X1 U575 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U576 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U577 ( .A(n732), .B(n485), .ZN(n640) );
  OR2_X2 U578 ( .A1(n640), .A2(G902), .ZN(n486) );
  XNOR2_X2 U579 ( .A(n486), .B(G472), .ZN(n534) );
  XNOR2_X1 U580 ( .A(n534), .B(KEYINPUT6), .ZN(n518) );
  INV_X1 U581 ( .A(n518), .ZN(n575) );
  NOR2_X1 U582 ( .A1(n487), .A2(n575), .ZN(n488) );
  NAND2_X1 U583 ( .A1(n491), .A2(n488), .ZN(n597) );
  XNOR2_X1 U584 ( .A(n597), .B(G101), .ZN(G3) );
  OR2_X1 U585 ( .A1(n514), .A2(n534), .ZN(n489) );
  NOR2_X1 U586 ( .A1(n587), .A2(n489), .ZN(n490) );
  XOR2_X1 U587 ( .A(G110), .B(n581), .Z(G12) );
  NAND2_X1 U588 ( .A1(G953), .A2(G900), .ZN(n492) );
  NAND2_X1 U589 ( .A1(n589), .A2(n385), .ZN(n494) );
  NAND2_X1 U590 ( .A1(n514), .A2(n673), .ZN(n677) );
  NAND2_X1 U591 ( .A1(n534), .A2(n687), .ZN(n496) );
  INV_X1 U592 ( .A(n520), .ZN(n499) );
  AND2_X1 U593 ( .A1(n499), .A2(n519), .ZN(n670) );
  NAND2_X1 U594 ( .A1(n530), .A2(n670), .ZN(n572) );
  XOR2_X1 U595 ( .A(G134), .B(KEYINPUT113), .Z(n500) );
  XNOR2_X1 U596 ( .A(n572), .B(n500), .ZN(G36) );
  XNOR2_X1 U597 ( .A(G122), .B(KEYINPUT127), .ZN(n513) );
  INV_X1 U598 ( .A(n677), .ZN(n501) );
  AND2_X1 U599 ( .A1(n501), .A2(n587), .ZN(n502) );
  NAND2_X1 U600 ( .A1(n502), .A2(n575), .ZN(n505) );
  XNOR2_X1 U601 ( .A(KEYINPUT104), .B(KEYINPUT33), .ZN(n503) );
  XNOR2_X1 U602 ( .A(n503), .B(KEYINPUT75), .ZN(n504) );
  XNOR2_X1 U603 ( .A(n505), .B(n504), .ZN(n705) );
  NOR2_X1 U604 ( .A1(n705), .A2(n592), .ZN(n509) );
  XNOR2_X1 U605 ( .A(KEYINPUT83), .B(KEYINPUT34), .ZN(n507) );
  XNOR2_X1 U606 ( .A(n507), .B(KEYINPUT76), .ZN(n508) );
  XNOR2_X1 U607 ( .A(n509), .B(n508), .ZN(n510) );
  OR2_X1 U608 ( .A1(n520), .A2(n519), .ZN(n548) );
  NOR2_X1 U609 ( .A1(n510), .A2(n548), .ZN(n512) );
  XNOR2_X1 U610 ( .A(KEYINPUT88), .B(KEYINPUT35), .ZN(n511) );
  XNOR2_X1 U611 ( .A(n512), .B(n511), .ZN(n605) );
  XOR2_X1 U612 ( .A(n513), .B(n605), .Z(G24) );
  INV_X1 U613 ( .A(n514), .ZN(n516) );
  NAND2_X1 U614 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U615 ( .A(n517), .B(KEYINPUT70), .ZN(n535) );
  NOR2_X1 U616 ( .A1(n535), .A2(n518), .ZN(n523) );
  INV_X1 U617 ( .A(n519), .ZN(n521) );
  INV_X1 U618 ( .A(KEYINPUT105), .ZN(n522) );
  XNOR2_X2 U619 ( .A(n544), .B(n522), .ZN(n667) );
  NAND2_X1 U620 ( .A1(n560), .A2(n687), .ZN(n524) );
  XOR2_X1 U621 ( .A(KEYINPUT106), .B(n524), .Z(n525) );
  AND2_X1 U622 ( .A1(n525), .A2(n678), .ZN(n527) );
  XNOR2_X1 U623 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n526) );
  XNOR2_X1 U624 ( .A(n527), .B(n526), .ZN(n529) );
  INV_X1 U625 ( .A(n528), .ZN(n547) );
  NAND2_X1 U626 ( .A1(n529), .A2(n547), .ZN(n573) );
  XNOR2_X1 U627 ( .A(n573), .B(G140), .ZN(G42) );
  NAND2_X1 U628 ( .A1(n530), .A2(n544), .ZN(n532) );
  INV_X1 U629 ( .A(KEYINPUT40), .ZN(n531) );
  INV_X1 U630 ( .A(n534), .ZN(n586) );
  NOR2_X2 U631 ( .A1(n535), .A2(n586), .ZN(n536) );
  XNOR2_X1 U632 ( .A(n536), .B(KEYINPUT28), .ZN(n542) );
  XNOR2_X1 U633 ( .A(n589), .B(KEYINPUT108), .ZN(n540) );
  NAND2_X1 U634 ( .A1(n542), .A2(n540), .ZN(n537) );
  NOR2_X1 U635 ( .A1(n706), .A2(n537), .ZN(n538) );
  XNOR2_X1 U636 ( .A(n538), .B(KEYINPUT42), .ZN(n744) );
  NOR2_X2 U637 ( .A1(n649), .A2(n744), .ZN(n539) );
  XNOR2_X1 U638 ( .A(n539), .B(KEYINPUT46), .ZN(n569) );
  NAND2_X1 U639 ( .A1(n542), .A2(n541), .ZN(n661) );
  NAND2_X1 U640 ( .A1(n661), .A2(KEYINPUT47), .ZN(n543) );
  XNOR2_X1 U641 ( .A(n543), .B(KEYINPUT86), .ZN(n546) );
  NOR2_X1 U642 ( .A1(n670), .A2(n544), .ZN(n692) );
  NAND2_X1 U643 ( .A1(n692), .A2(KEYINPUT47), .ZN(n545) );
  NAND2_X1 U644 ( .A1(n546), .A2(n545), .ZN(n551) );
  NOR2_X1 U645 ( .A1(n548), .A2(n547), .ZN(n549) );
  AND2_X1 U646 ( .A1(n550), .A2(n549), .ZN(n664) );
  OR2_X2 U647 ( .A1(n551), .A2(n664), .ZN(n552) );
  INV_X1 U648 ( .A(KEYINPUT87), .ZN(n553) );
  XNOR2_X1 U649 ( .A(n692), .B(n553), .ZN(n594) );
  XNOR2_X1 U650 ( .A(KEYINPUT47), .B(KEYINPUT66), .ZN(n554) );
  OR2_X1 U651 ( .A1(n594), .A2(n554), .ZN(n555) );
  NOR2_X1 U652 ( .A1(n661), .A2(n555), .ZN(n557) );
  INV_X1 U653 ( .A(KEYINPUT78), .ZN(n556) );
  XNOR2_X1 U654 ( .A(n557), .B(n556), .ZN(n558) );
  NAND2_X1 U655 ( .A1(n559), .A2(n558), .ZN(n567) );
  XNOR2_X1 U656 ( .A(n560), .B(KEYINPUT109), .ZN(n562) );
  NOR2_X1 U657 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U658 ( .A(n563), .B(KEYINPUT36), .ZN(n564) );
  NAND2_X1 U659 ( .A1(n564), .A2(n587), .ZN(n566) );
  INV_X1 U660 ( .A(KEYINPUT110), .ZN(n565) );
  NAND2_X1 U661 ( .A1(n569), .A2(n568), .ZN(n571) );
  INV_X1 U662 ( .A(KEYINPUT48), .ZN(n570) );
  AND2_X1 U663 ( .A1(n573), .A2(n572), .ZN(n574) );
  OR2_X1 U664 ( .A1(n674), .A2(n678), .ZN(n576) );
  NOR2_X1 U665 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U666 ( .A1(n578), .A2(n577), .ZN(n580) );
  INV_X1 U667 ( .A(KEYINPUT32), .ZN(n579) );
  INV_X1 U668 ( .A(n647), .ZN(n583) );
  XNOR2_X2 U669 ( .A(n584), .B(KEYINPUT91), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n600), .A2(n605), .ZN(n585) );
  NOR2_X1 U671 ( .A1(n677), .A2(n586), .ZN(n588) );
  NAND2_X1 U672 ( .A1(n588), .A2(n587), .ZN(n682) );
  NOR2_X1 U673 ( .A1(n677), .A2(n534), .ZN(n590) );
  NAND2_X1 U674 ( .A1(n590), .A2(n589), .ZN(n591) );
  INV_X1 U675 ( .A(KEYINPUT101), .ZN(n593) );
  INV_X1 U676 ( .A(n594), .ZN(n595) );
  NAND2_X1 U677 ( .A1(n596), .A2(n595), .ZN(n598) );
  NOR2_X1 U678 ( .A1(n601), .A2(KEYINPUT44), .ZN(n599) );
  NAND2_X1 U679 ( .A1(n600), .A2(n599), .ZN(n604) );
  INV_X1 U680 ( .A(n600), .ZN(n602) );
  INV_X1 U681 ( .A(KEYINPUT90), .ZN(n601) );
  NAND2_X1 U682 ( .A1(n602), .A2(n601), .ZN(n603) );
  INV_X1 U683 ( .A(n609), .ZN(n611) );
  NOR2_X4 U684 ( .A1(n613), .A2(n612), .ZN(n650) );
  NAND2_X1 U685 ( .A1(n650), .A2(G475), .ZN(n617) );
  XNOR2_X1 U686 ( .A(KEYINPUT120), .B(KEYINPUT59), .ZN(n614) );
  XNOR2_X1 U687 ( .A(n615), .B(n614), .ZN(n616) );
  XNOR2_X1 U688 ( .A(n617), .B(n616), .ZN(n619) );
  XOR2_X1 U689 ( .A(KEYINPUT121), .B(KEYINPUT60), .Z(n620) );
  XNOR2_X1 U690 ( .A(n621), .B(n620), .ZN(G60) );
  NAND2_X1 U691 ( .A1(n650), .A2(G210), .ZN(n627) );
  BUF_X1 U692 ( .A(n622), .Z(n625) );
  XNOR2_X1 U693 ( .A(KEYINPUT93), .B(KEYINPUT54), .ZN(n623) );
  XNOR2_X1 U694 ( .A(n623), .B(KEYINPUT55), .ZN(n624) );
  XNOR2_X1 U695 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U696 ( .A(n627), .B(n626), .ZN(n628) );
  XOR2_X1 U697 ( .A(KEYINPUT89), .B(KEYINPUT56), .Z(n629) );
  XNOR2_X1 U698 ( .A(n630), .B(n629), .ZN(G51) );
  NAND2_X1 U699 ( .A1(n650), .A2(G469), .ZN(n636) );
  XNOR2_X1 U700 ( .A(KEYINPUT118), .B(KEYINPUT57), .ZN(n633) );
  XNOR2_X1 U701 ( .A(KEYINPUT58), .B(KEYINPUT117), .ZN(n632) );
  XNOR2_X1 U702 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U703 ( .A(n636), .B(n635), .ZN(n637) );
  INV_X1 U704 ( .A(KEYINPUT119), .ZN(n638) );
  XNOR2_X1 U705 ( .A(n639), .B(n638), .ZN(G54) );
  NAND2_X1 U706 ( .A1(n650), .A2(G472), .ZN(n642) );
  XNOR2_X1 U707 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U708 ( .A(KEYINPUT94), .B(KEYINPUT63), .ZN(n644) );
  XOR2_X1 U709 ( .A(n644), .B(KEYINPUT92), .Z(n645) );
  XNOR2_X1 U710 ( .A(n646), .B(n645), .ZN(G57) );
  XOR2_X1 U711 ( .A(n648), .B(G119), .Z(G21) );
  XOR2_X1 U712 ( .A(G131), .B(n350), .Z(G33) );
  NAND2_X1 U713 ( .A1(n713), .A2(G478), .ZN(n653) );
  XOR2_X1 U714 ( .A(n651), .B(KEYINPUT122), .Z(n652) );
  XNOR2_X1 U715 ( .A(n653), .B(n652), .ZN(n654) );
  NOR2_X1 U716 ( .A1(n654), .A2(n717), .ZN(G63) );
  NAND2_X1 U717 ( .A1(n656), .A2(n667), .ZN(n655) );
  XNOR2_X1 U718 ( .A(n655), .B(G104), .ZN(G6) );
  XOR2_X1 U719 ( .A(KEYINPUT26), .B(KEYINPUT111), .Z(n658) );
  NAND2_X1 U720 ( .A1(n670), .A2(n656), .ZN(n657) );
  XNOR2_X1 U721 ( .A(n658), .B(n657), .ZN(n660) );
  XOR2_X1 U722 ( .A(G107), .B(KEYINPUT27), .Z(n659) );
  XNOR2_X1 U723 ( .A(n660), .B(n659), .ZN(G9) );
  XOR2_X1 U724 ( .A(G128), .B(KEYINPUT29), .Z(n663) );
  INV_X1 U725 ( .A(n661), .ZN(n665) );
  NAND2_X1 U726 ( .A1(n665), .A2(n670), .ZN(n662) );
  XNOR2_X1 U727 ( .A(n663), .B(n662), .ZN(G30) );
  XOR2_X1 U728 ( .A(G143), .B(n664), .Z(G45) );
  NAND2_X1 U729 ( .A1(n665), .A2(n667), .ZN(n666) );
  XNOR2_X1 U730 ( .A(n666), .B(G146), .ZN(G48) );
  NAND2_X1 U731 ( .A1(n671), .A2(n667), .ZN(n668) );
  XNOR2_X1 U732 ( .A(n668), .B(KEYINPUT112), .ZN(n669) );
  XNOR2_X1 U733 ( .A(G113), .B(n669), .ZN(G15) );
  NAND2_X1 U734 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U735 ( .A(n672), .B(G116), .ZN(G18) );
  NOR2_X1 U736 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U737 ( .A(KEYINPUT49), .B(n675), .Z(n676) );
  NOR2_X1 U738 ( .A1(n676), .A2(n534), .ZN(n681) );
  NAND2_X1 U739 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U740 ( .A(n679), .B(KEYINPUT50), .ZN(n680) );
  NAND2_X1 U741 ( .A1(n681), .A2(n680), .ZN(n683) );
  NAND2_X1 U742 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U743 ( .A(KEYINPUT51), .B(n684), .ZN(n685) );
  NOR2_X1 U744 ( .A1(n706), .A2(n685), .ZN(n686) );
  XOR2_X1 U745 ( .A(KEYINPUT114), .B(n686), .Z(n699) );
  NOR2_X1 U746 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U747 ( .A1(n690), .A2(n689), .ZN(n694) );
  NOR2_X1 U748 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U749 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U750 ( .A(KEYINPUT115), .B(n695), .ZN(n697) );
  INV_X1 U751 ( .A(n705), .ZN(n696) );
  NAND2_X1 U752 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U753 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U754 ( .A(KEYINPUT52), .B(n700), .Z(n703) );
  NAND2_X1 U755 ( .A1(G952), .A2(n701), .ZN(n702) );
  NOR2_X1 U756 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U757 ( .A1(G953), .A2(n704), .ZN(n708) );
  OR2_X1 U758 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U759 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U760 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U761 ( .A(n711), .B(KEYINPUT53), .ZN(n712) );
  XNOR2_X1 U762 ( .A(n712), .B(KEYINPUT116), .ZN(G75) );
  NAND2_X1 U763 ( .A1(n713), .A2(G217), .ZN(n715) );
  XNOR2_X1 U764 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U765 ( .A1(n717), .A2(n716), .ZN(G66) );
  NAND2_X1 U766 ( .A1(n718), .A2(n738), .ZN(n722) );
  NAND2_X1 U767 ( .A1(G953), .A2(G224), .ZN(n719) );
  XNOR2_X1 U768 ( .A(KEYINPUT61), .B(n719), .ZN(n720) );
  NAND2_X1 U769 ( .A1(n720), .A2(G898), .ZN(n721) );
  NAND2_X1 U770 ( .A1(n722), .A2(n721), .ZN(n730) );
  XNOR2_X1 U771 ( .A(KEYINPUT124), .B(KEYINPUT123), .ZN(n724) );
  XOR2_X1 U772 ( .A(n724), .B(n723), .Z(n725) );
  XNOR2_X1 U773 ( .A(n726), .B(n725), .ZN(n728) );
  NOR2_X1 U774 ( .A1(n738), .A2(G898), .ZN(n727) );
  NOR2_X1 U775 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U776 ( .A(n730), .B(n729), .ZN(G69) );
  XNOR2_X1 U777 ( .A(n732), .B(n731), .ZN(n737) );
  XOR2_X1 U778 ( .A(KEYINPUT125), .B(n737), .Z(n733) );
  XNOR2_X1 U779 ( .A(G227), .B(n733), .ZN(n734) );
  NAND2_X1 U780 ( .A1(n734), .A2(G900), .ZN(n735) );
  NAND2_X1 U781 ( .A1(n735), .A2(G953), .ZN(n736) );
  XNOR2_X1 U782 ( .A(n736), .B(KEYINPUT126), .ZN(n741) );
  XNOR2_X1 U783 ( .A(n609), .B(n737), .ZN(n739) );
  NAND2_X1 U784 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U785 ( .A1(n741), .A2(n740), .ZN(G72) );
  XNOR2_X1 U786 ( .A(G125), .B(KEYINPUT37), .ZN(n743) );
  XNOR2_X1 U787 ( .A(n743), .B(n742), .ZN(G27) );
  XOR2_X1 U788 ( .A(G137), .B(n744), .Z(G39) );
endmodule

