//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923;
  NAND2_X1  g000(.A1(G85gat), .A2(G92gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT7), .ZN(new_n203));
  INV_X1    g002(.A(G99gat), .ZN(new_n204));
  INV_X1    g003(.A(G106gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT8), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(KEYINPUT99), .B(G85gat), .Z(new_n207));
  OAI211_X1 g006(.A(new_n203), .B(new_n206), .C1(G92gat), .C2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G99gat), .B(G106gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT91), .B(G50gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n212), .B1(new_n213), .B2(G43gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(G43gat), .B(G50gat), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n215), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n216));
  NOR3_X1   g015(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(KEYINPUT92), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n214), .B(new_n216), .C1(new_n218), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G29gat), .A2(G36gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(new_n220), .B2(new_n217), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(KEYINPUT15), .A3(new_n215), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT17), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n221), .A2(KEYINPUT17), .A3(new_n224), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(G232gat), .A2(G233gat), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n210), .A2(new_n225), .B1(KEYINPUT41), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n232), .B(G190gat), .ZN(new_n233));
  INV_X1    g032(.A(G218gat), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT98), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(new_n234), .B2(new_n233), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n230), .A2(KEYINPUT41), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n236), .A2(new_n237), .ZN(new_n240));
  XOR2_X1   g039(.A(G134gat), .B(G162gat), .Z(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NOR3_X1   g041(.A1(new_n239), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n242), .B1(new_n239), .B2(new_n240), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OR2_X1    g045(.A1(G57gat), .A2(G64gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(G57gat), .A2(G64gat), .ZN(new_n248));
  AND2_X1   g047(.A1(G71gat), .A2(G78gat), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n247), .B(new_n248), .C1(new_n249), .C2(KEYINPUT9), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT96), .ZN(new_n251));
  NOR2_X1   g050(.A1(G71gat), .A2(G78gat), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n249), .A2(new_n252), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n255), .A2(KEYINPUT21), .ZN(new_n256));
  NAND2_X1  g055(.A1(G231gat), .A2(G233gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G127gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(G183gat), .B(G211gat), .Z(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G8gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(G15gat), .B(G22gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT16), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n264), .B1(new_n265), .B2(G1gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT93), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n263), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(G1gat), .B2(new_n264), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n270), .B1(KEYINPUT21), .B2(new_n255), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT97), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(G155gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n272), .B(new_n274), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n262), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n262), .A2(new_n275), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n246), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT100), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n208), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n255), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n211), .B(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G230gat), .ZN(new_n284));
  INV_X1    g083(.A(G233gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n287), .B(KEYINPUT101), .Z(new_n288));
  NAND3_X1  g087(.A1(new_n210), .A2(KEYINPUT10), .A3(new_n255), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(new_n283), .B2(KEYINPUT10), .ZN(new_n290));
  INV_X1    g089(.A(new_n286), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OR2_X1    g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  XOR2_X1   g092(.A(G120gat), .B(G148gat), .Z(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT102), .ZN(new_n295));
  XNOR2_X1  g094(.A(G176gat), .B(G204gat), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n295), .B(new_n296), .Z(new_n297));
  OR2_X1    g096(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n293), .A2(new_n297), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n279), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G1gat), .B(G29gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n304), .B(KEYINPUT0), .ZN(new_n305));
  XNOR2_X1  g104(.A(G57gat), .B(G85gat), .ZN(new_n306));
  XOR2_X1   g105(.A(new_n305), .B(new_n306), .Z(new_n307));
  NAND2_X1  g106(.A1(G225gat), .A2(G233gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  AND2_X1   g108(.A1(G113gat), .A2(G120gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(G113gat), .A2(G120gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT67), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT1), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G134gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n259), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G127gat), .A2(G134gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(G127gat), .A2(G134gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(G127gat), .A2(G134gat), .ZN(new_n322));
  NOR3_X1   g121(.A1(new_n321), .A2(new_n322), .A3(KEYINPUT66), .ZN(new_n323));
  XNOR2_X1  g122(.A(G113gat), .B(G120gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n314), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT66), .B1(new_n312), .B2(new_n313), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n320), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G155gat), .B(G162gat), .ZN(new_n328));
  INV_X1    g127(.A(G141gat), .ZN(new_n329));
  INV_X1    g128(.A(G148gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G141gat), .A2(G148gat), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n328), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT77), .B(G155gat), .ZN(new_n334));
  INV_X1    g133(.A(G162gat), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT2), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT76), .B1(G155gat), .B2(G162gat), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n337), .B1(new_n328), .B2(KEYINPUT76), .ZN(new_n338));
  NAND2_X1  g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT2), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(new_n331), .A3(new_n332), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n333), .A2(new_n336), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n327), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT66), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n317), .A2(new_n344), .A3(new_n318), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT1), .B1(new_n345), .B2(new_n312), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n344), .B1(new_n324), .B2(KEYINPUT67), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n346), .A2(new_n347), .B1(new_n315), .B2(new_n319), .ZN(new_n348));
  AND2_X1   g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(G155gat), .A2(G162gat), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT76), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n337), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n341), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT2), .ZN(new_n354));
  INV_X1    g153(.A(G155gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT77), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G155gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n354), .B1(new_n359), .B2(G162gat), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n328), .A2(new_n331), .A3(new_n332), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n353), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n348), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n309), .B1(new_n343), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT79), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT79), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n366), .B(new_n309), .C1(new_n343), .C2(new_n363), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n362), .A2(KEYINPUT3), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT3), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n353), .B(new_n370), .C1(new_n360), .C2(new_n361), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(new_n371), .A3(new_n348), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n348), .A2(new_n362), .A3(KEYINPUT4), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT4), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n374), .B1(new_n327), .B2(new_n342), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n308), .B(new_n372), .C1(new_n373), .C2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT78), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n374), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT4), .B1(new_n348), .B2(new_n362), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n381), .A2(KEYINPUT78), .A3(new_n308), .A4(new_n372), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n368), .A2(new_n378), .A3(new_n382), .A4(KEYINPUT5), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT5), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n381), .A2(new_n384), .A3(new_n308), .A4(new_n372), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n307), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  XOR2_X1   g185(.A(KEYINPUT80), .B(KEYINPUT6), .Z(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n383), .A2(new_n385), .ZN(new_n390));
  INV_X1    g189(.A(new_n307), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n385), .A2(new_n307), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n388), .B1(new_n383), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n392), .B1(KEYINPUT81), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(KEYINPUT81), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n389), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(G211gat), .A2(G218gat), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT22), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(G197gat), .A2(G204gat), .ZN(new_n402));
  AND2_X1   g201(.A1(G197gat), .A2(G204gat), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(G211gat), .B(G218gat), .Z(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G211gat), .B(G218gat), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n407), .B(new_n401), .C1(new_n402), .C2(new_n403), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(G226gat), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n411), .A2(new_n285), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT65), .ZN(new_n413));
  INV_X1    g212(.A(G190gat), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT27), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n413), .B(new_n414), .C1(new_n415), .C2(G183gat), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT28), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(G183gat), .ZN(new_n419));
  AOI21_X1  g218(.A(G190gat), .B1(new_n419), .B2(KEYINPUT27), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n415), .A2(G183gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n420), .A2(KEYINPUT65), .A3(new_n417), .A4(new_n421), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n425), .B1(G169gat), .B2(G176gat), .ZN(new_n426));
  NOR2_X1   g225(.A1(G169gat), .A2(G176gat), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n427), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n423), .A2(new_n424), .A3(new_n426), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G183gat), .A2(G190gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT24), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT24), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n432), .A2(G183gat), .A3(G190gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n414), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT64), .ZN(new_n436));
  NOR2_X1   g235(.A1(G183gat), .A2(G190gat), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT64), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n434), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(G169gat), .ZN(new_n441));
  INV_X1    g240(.A(G176gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT23), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT23), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n444), .B1(G169gat), .B2(G176gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(G169gat), .A2(G176gat), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT25), .B1(new_n440), .B2(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n443), .A2(new_n445), .A3(KEYINPUT25), .A4(new_n446), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n434), .B2(new_n435), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n429), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT73), .B(KEYINPUT29), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n412), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n412), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n434), .A2(new_n435), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n455), .A2(new_n447), .A3(KEYINPUT25), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n437), .B(KEYINPUT64), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n457), .B1(new_n458), .B2(new_n434), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n456), .B1(new_n459), .B2(KEYINPUT25), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n454), .B1(new_n460), .B2(new_n429), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n410), .B1(new_n453), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n451), .A2(new_n412), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT29), .B1(new_n460), .B2(new_n429), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n409), .B(new_n463), .C1(new_n464), .C2(new_n412), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(G8gat), .B(G36gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n467), .B(KEYINPUT74), .ZN(new_n468));
  XNOR2_X1  g267(.A(G64gat), .B(G92gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(KEYINPUT75), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n462), .A2(new_n465), .A3(new_n470), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT30), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n398), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT83), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n409), .A2(new_n452), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n342), .B1(new_n480), .B2(new_n370), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n409), .B1(new_n371), .B2(new_n452), .ZN(new_n482));
  INV_X1    g281(.A(G228gat), .ZN(new_n483));
  OAI22_X1  g282(.A1(new_n481), .A2(new_n482), .B1(new_n483), .B2(new_n285), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n371), .A2(new_n452), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n410), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n483), .A2(new_n285), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT29), .B1(new_n406), .B2(new_n408), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n362), .B1(new_n488), .B2(KEYINPUT3), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n484), .A2(new_n490), .A3(G22gat), .ZN(new_n491));
  XOR2_X1   g290(.A(G78gat), .B(G106gat), .Z(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(KEYINPUT82), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT31), .B(G50gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(G22gat), .B1(new_n484), .B2(new_n490), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n479), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n484), .A2(new_n490), .ZN(new_n499));
  INV_X1    g298(.A(G22gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n501), .A2(KEYINPUT83), .A3(new_n495), .A4(new_n491), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n499), .ZN(new_n504));
  NAND2_X1  g303(.A1(KEYINPUT84), .A2(G22gat), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n495), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n506), .B1(new_n504), .B2(new_n505), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n478), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT37), .ZN(new_n511));
  OR3_X1    g310(.A1(new_n453), .A2(new_n461), .A3(new_n410), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n512), .A2(KEYINPUT88), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n463), .B1(new_n464), .B2(new_n412), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n512), .A2(KEYINPUT88), .B1(new_n514), .B2(new_n410), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n511), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT38), .ZN(new_n517));
  XOR2_X1   g316(.A(KEYINPUT89), .B(KEYINPUT37), .Z(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n517), .B(new_n471), .C1(new_n466), .C2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n474), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n466), .A2(new_n519), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n522), .A2(new_n470), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n466), .A2(KEYINPUT37), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n517), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT86), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n392), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n386), .A2(KEYINPUT86), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n394), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n526), .A2(new_n530), .A3(new_n389), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT85), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n372), .B1(new_n373), .B2(new_n375), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n532), .B1(new_n533), .B2(new_n309), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n533), .A2(new_n532), .A3(new_n309), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT39), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n391), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT87), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n343), .A2(new_n363), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n538), .B1(new_n541), .B2(new_n308), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n535), .A2(new_n536), .A3(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n539), .A2(new_n540), .A3(KEYINPUT40), .A4(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n536), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n538), .B1(new_n545), .B2(new_n534), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n546), .A2(new_n543), .A3(KEYINPUT40), .A4(new_n307), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT87), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n386), .B(new_n527), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n546), .A2(new_n543), .A3(new_n307), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT40), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n473), .A2(new_n475), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n549), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n531), .A2(new_n554), .A3(new_n508), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT34), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT68), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n327), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n348), .A2(KEYINPUT68), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(new_n451), .A3(new_n559), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n460), .A2(KEYINPUT68), .A3(new_n348), .A4(new_n429), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G227gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n563), .A2(new_n285), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n556), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  AOI211_X1 g365(.A(KEYINPUT34), .B(new_n564), .C1(new_n560), .C2(new_n561), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n560), .A2(new_n564), .A3(new_n561), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT32), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT69), .B(KEYINPUT33), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G15gat), .B(G43gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(G71gat), .B(G99gat), .Z(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n570), .A2(new_n572), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n577), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n569), .B(KEYINPUT32), .C1(new_n571), .C2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n568), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT72), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n568), .A2(new_n578), .A3(KEYINPUT72), .A4(new_n580), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n566), .ZN(new_n586));
  INV_X1    g385(.A(new_n567), .ZN(new_n587));
  AOI22_X1  g386(.A1(new_n578), .A2(new_n580), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT36), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n510), .A2(new_n555), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT35), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n588), .B1(new_n503), .B2(new_n507), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(new_n585), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT90), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT90), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n595), .A2(new_n585), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n383), .A2(new_n393), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n387), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT81), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n604), .A2(new_n392), .A3(new_n396), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n476), .B1(new_n605), .B2(new_n389), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n594), .B1(new_n600), .B2(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n530), .A2(new_n389), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n477), .A2(new_n594), .A3(new_n585), .A4(new_n595), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n593), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n270), .B(new_n225), .ZN(new_n612));
  XOR2_X1   g411(.A(KEYINPUT94), .B(KEYINPUT13), .Z(new_n613));
  NAND2_X1  g412(.A1(G229gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n616), .B(KEYINPUT95), .Z(new_n617));
  AOI21_X1  g416(.A(new_n270), .B1(new_n226), .B2(new_n225), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n618), .A2(new_n228), .B1(new_n270), .B2(new_n225), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n619), .A2(new_n614), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n620), .A2(KEYINPUT18), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(KEYINPUT18), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G113gat), .B(G141gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(G197gat), .ZN(new_n625));
  XOR2_X1   g424(.A(KEYINPUT11), .B(G169gat), .Z(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n627), .B(KEYINPUT12), .Z(new_n628));
  OR2_X1    g427(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n623), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n611), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n398), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n303), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g434(.A1(new_n303), .A2(new_n632), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n636), .A2(new_n477), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n637), .A2(new_n263), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n638), .B(KEYINPUT103), .Z(new_n639));
  XOR2_X1   g438(.A(KEYINPUT16), .B(G8gat), .Z(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT42), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(G1325gat));
  OAI21_X1  g442(.A(G15gat), .B1(new_n636), .B2(new_n592), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n590), .A2(G15gat), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n303), .A2(new_n632), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(G1326gat));
  NOR2_X1   g446(.A1(new_n636), .A2(new_n508), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT104), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT43), .B(G22gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(G1327gat));
  INV_X1    g450(.A(G29gat), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n653), .B1(new_n611), .B2(new_n246), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT106), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n607), .A2(new_n655), .A3(new_n610), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n595), .A2(new_n585), .A3(new_n598), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n598), .B1(new_n595), .B2(new_n585), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT35), .B1(new_n659), .B2(new_n478), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n608), .A2(new_n609), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT106), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n593), .B1(new_n656), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT107), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n246), .A2(new_n653), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n663), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n510), .A2(new_n555), .A3(new_n592), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n655), .B1(new_n607), .B2(new_n610), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n660), .A2(KEYINPUT106), .A3(new_n661), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT107), .B1(new_n671), .B2(new_n665), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n654), .B1(new_n667), .B2(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n278), .B(KEYINPUT105), .Z(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(new_n631), .A3(new_n301), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT108), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT108), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(new_n673), .B2(new_n675), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n633), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n652), .B1(new_n680), .B2(KEYINPUT109), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n681), .B1(KEYINPUT109), .B2(new_n680), .ZN(new_n682));
  INV_X1    g481(.A(new_n246), .ZN(new_n683));
  INV_X1    g482(.A(new_n278), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n683), .A2(new_n684), .A3(new_n300), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n632), .A2(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n686), .A2(G29gat), .A3(new_n398), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT45), .Z(new_n688));
  NAND2_X1  g487(.A1(new_n682), .A2(new_n688), .ZN(G1328gat));
  NAND3_X1  g488(.A1(new_n677), .A2(new_n476), .A3(new_n679), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(G36gat), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n686), .A2(G36gat), .A3(new_n477), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT46), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(G1329gat));
  NOR3_X1   g493(.A1(new_n686), .A2(G43gat), .A3(new_n590), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n676), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT112), .B1(new_n697), .B2(new_n592), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(G43gat), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n697), .A2(KEYINPUT112), .A3(new_n592), .ZN(new_n700));
  OAI211_X1 g499(.A(KEYINPUT47), .B(new_n696), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n592), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n677), .A2(new_n702), .A3(new_n679), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n703), .A2(KEYINPUT111), .A3(G43gat), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT111), .B1(new_n703), .B2(G43gat), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n704), .A2(new_n705), .A3(new_n695), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n701), .B1(new_n706), .B2(new_n707), .ZN(G1330gat));
  OAI21_X1  g507(.A(new_n213), .B1(new_n697), .B2(new_n508), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n686), .A2(new_n508), .A3(new_n213), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n709), .A2(KEYINPUT48), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n677), .A2(new_n509), .A3(new_n679), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n710), .B1(new_n713), .B2(new_n213), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n712), .B1(new_n714), .B2(new_n715), .ZN(G1331gat));
  INV_X1    g515(.A(new_n631), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n663), .A2(new_n717), .A3(new_n279), .A4(new_n300), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n718), .A2(KEYINPUT114), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(KEYINPUT114), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n633), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g523(.A1(new_n721), .A2(new_n477), .ZN(new_n725));
  NOR2_X1   g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  AND2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n725), .B2(new_n726), .ZN(G1333gat));
  OAI21_X1  g528(.A(G71gat), .B1(new_n721), .B2(new_n592), .ZN(new_n730));
  OR2_X1    g529(.A1(new_n590), .A2(G71gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n721), .B2(new_n731), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g532(.A1(new_n722), .A2(new_n509), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g534(.A1(new_n684), .A2(new_n631), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n300), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n667), .A2(new_n672), .ZN(new_n738));
  INV_X1    g537(.A(new_n654), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n207), .B1(new_n741), .B2(new_n398), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT51), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n663), .A2(new_n743), .A3(new_n246), .A4(new_n736), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n246), .A2(new_n736), .ZN(new_n745));
  OAI21_X1  g544(.A(KEYINPUT51), .B1(new_n671), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n744), .A2(new_n300), .A3(new_n746), .ZN(new_n747));
  OR3_X1    g546(.A1(new_n747), .A2(new_n398), .A3(new_n207), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n742), .A2(new_n748), .ZN(G1336gat));
  OAI21_X1  g548(.A(G92gat), .B1(new_n741), .B2(new_n477), .ZN(new_n750));
  OR3_X1    g549(.A1(new_n747), .A2(G92gat), .A3(new_n477), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT115), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n753), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n752), .B(new_n755), .ZN(G1337gat));
  NOR3_X1   g555(.A1(new_n741), .A2(new_n204), .A3(new_n592), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n747), .A2(new_n590), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n757), .B1(new_n204), .B2(new_n758), .ZN(G1338gat));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n508), .A2(G106gat), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n744), .A2(new_n746), .A3(new_n300), .A4(new_n761), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n673), .A2(new_n508), .A3(new_n737), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n760), .B(new_n762), .C1(new_n763), .C2(new_n205), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT117), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n205), .B1(new_n740), .B2(new_n509), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n760), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n762), .A2(KEYINPUT116), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n763), .B2(new_n205), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n765), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n738), .A2(new_n739), .ZN(new_n772));
  INV_X1    g571(.A(new_n737), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(new_n509), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(new_n767), .A3(G106gat), .ZN(new_n775));
  AND4_X1   g574(.A1(new_n765), .A2(new_n770), .A3(KEYINPUT53), .A4(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n764), .B1(new_n771), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT118), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g578(.A(KEYINPUT118), .B(new_n764), .C1(new_n771), .C2(new_n776), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(G1339gat));
  NOR2_X1   g580(.A1(new_n302), .A2(new_n631), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n292), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n291), .B2(new_n290), .ZN(new_n786));
  INV_X1    g585(.A(new_n297), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n787), .B1(new_n292), .B2(new_n784), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n786), .A2(KEYINPUT55), .A3(new_n788), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n298), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT119), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n298), .A2(new_n791), .A3(KEYINPUT119), .A4(new_n792), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n631), .A3(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n619), .A2(new_n614), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n612), .A2(new_n615), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n627), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n629), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n300), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n246), .B1(new_n797), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n246), .A2(new_n801), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n795), .A2(new_n796), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n674), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n398), .B1(new_n783), .B2(new_n807), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n808), .A2(new_n477), .A3(new_n600), .ZN(new_n809));
  AOI21_X1  g608(.A(G113gat), .B1(new_n809), .B2(new_n631), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n783), .A2(new_n807), .ZN(new_n811));
  INV_X1    g610(.A(new_n596), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n398), .A2(new_n476), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n631), .A2(G113gat), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n810), .B1(new_n816), .B2(new_n817), .ZN(G1340gat));
  AOI21_X1  g617(.A(G120gat), .B1(new_n809), .B2(new_n300), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n300), .A2(G120gat), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n816), .B2(new_n820), .ZN(G1341gat));
  INV_X1    g620(.A(new_n816), .ZN(new_n822));
  OAI21_X1  g621(.A(G127gat), .B1(new_n822), .B2(new_n674), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n809), .A2(new_n259), .A3(new_n684), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(G1342gat));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n316), .A3(new_n246), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n826), .A2(KEYINPUT56), .ZN(new_n827));
  OAI21_X1  g626(.A(G134gat), .B1(new_n822), .B2(new_n683), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(KEYINPUT56), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(G1343gat));
  INV_X1    g629(.A(new_n806), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n802), .B1(new_n793), .B2(new_n717), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n683), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n684), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n509), .B1(new_n834), .B2(new_n782), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT57), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n508), .B1(new_n783), .B2(new_n807), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n702), .A2(new_n815), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n836), .A2(new_n839), .A3(new_n631), .A4(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n329), .B1(new_n841), .B2(KEYINPUT121), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n842), .B1(KEYINPUT121), .B2(new_n841), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844));
  AND4_X1   g643(.A1(new_n477), .A2(new_n808), .A3(new_n509), .A4(new_n592), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(new_n329), .A3(new_n631), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n841), .A2(G141gat), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n846), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n849), .A2(KEYINPUT120), .A3(KEYINPUT58), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT120), .B1(new_n849), .B2(KEYINPUT58), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n847), .B1(new_n850), .B2(new_n851), .ZN(G1344gat));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n839), .A3(new_n840), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n853), .B(G148gat), .C1(new_n854), .C2(new_n301), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT122), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n804), .A2(new_n793), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n684), .B1(new_n857), .B2(new_n833), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n838), .B(new_n509), .C1(new_n858), .C2(new_n782), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n301), .A2(new_n702), .A3(new_n815), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n859), .B(new_n860), .C1(new_n837), .C2(new_n838), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(G148gat), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n856), .B1(new_n862), .B2(KEYINPUT59), .ZN(new_n863));
  AOI211_X1 g662(.A(KEYINPUT122), .B(new_n853), .C1(new_n861), .C2(G148gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n855), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n845), .A2(new_n330), .A3(new_n300), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1345gat));
  OAI21_X1  g666(.A(new_n359), .B1(new_n854), .B2(new_n674), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n845), .A2(new_n334), .A3(new_n684), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1346gat));
  NOR3_X1   g669(.A1(new_n854), .A2(new_n335), .A3(new_n683), .ZN(new_n871));
  AOI21_X1  g670(.A(G162gat), .B1(new_n845), .B2(new_n246), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(G1347gat));
  NAND2_X1  g672(.A1(new_n398), .A2(new_n476), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT123), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n811), .A2(new_n812), .A3(new_n875), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n876), .A2(new_n441), .A3(new_n717), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n633), .B1(new_n783), .B2(new_n807), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n878), .A2(new_n476), .A3(new_n600), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n631), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n877), .B1(new_n880), .B2(new_n441), .ZN(G1348gat));
  NOR3_X1   g680(.A1(new_n876), .A2(new_n442), .A3(new_n301), .ZN(new_n882));
  AOI21_X1  g681(.A(G176gat), .B1(new_n879), .B2(new_n300), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n883), .A2(KEYINPUT124), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(KEYINPUT124), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(G1349gat));
  NAND2_X1  g685(.A1(new_n419), .A2(KEYINPUT27), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n879), .A2(new_n887), .A3(new_n421), .A4(new_n684), .ZN(new_n888));
  OAI21_X1  g687(.A(G183gat), .B1(new_n876), .B2(new_n674), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g690(.A(G190gat), .B1(new_n876), .B2(new_n683), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT61), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n879), .A2(new_n414), .A3(new_n246), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1351gat));
  AND4_X1   g694(.A1(new_n476), .A2(new_n878), .A3(new_n509), .A4(new_n592), .ZN(new_n896));
  INV_X1    g695(.A(G197gat), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(new_n897), .A3(new_n631), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n875), .A2(new_n592), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n859), .B(new_n899), .C1(new_n837), .C2(new_n838), .ZN(new_n900));
  OAI21_X1  g699(.A(G197gat), .B1(new_n900), .B2(new_n717), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT125), .ZN(G1352gat));
  INV_X1    g702(.A(G204gat), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n896), .A2(new_n904), .A3(new_n300), .ZN(new_n905));
  XOR2_X1   g704(.A(new_n905), .B(KEYINPUT62), .Z(new_n906));
  OAI21_X1  g705(.A(G204gat), .B1(new_n900), .B2(new_n301), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1353gat));
  OAI21_X1  g707(.A(G211gat), .B1(new_n900), .B2(new_n278), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT126), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT63), .ZN(new_n911));
  OR3_X1    g710(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n909), .A2(new_n911), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT127), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT127), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n909), .A2(new_n915), .A3(new_n911), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n910), .B1(new_n909), .B2(new_n911), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n912), .A2(new_n914), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(G211gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n896), .A2(new_n919), .A3(new_n684), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1354gat));
  NAND3_X1  g720(.A1(new_n896), .A2(new_n234), .A3(new_n246), .ZN(new_n922));
  OAI21_X1  g721(.A(G218gat), .B1(new_n900), .B2(new_n683), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1355gat));
endmodule


