//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n996, new_n997;
  AOI21_X1  g000(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT96), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT98), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n202), .B(KEYINPUT96), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT98), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G71gat), .B(G78gat), .Z(new_n209));
  NAND2_X1  g008(.A1(KEYINPUT97), .A2(G57gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G64gat), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n210), .A2(G64gat), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n205), .A2(new_n208), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT99), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT99), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n205), .A2(new_n208), .A3(new_n216), .A4(new_n213), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(G57gat), .B(G64gat), .Z(new_n219));
  NAND2_X1  g018(.A1(new_n206), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n209), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT21), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G231gat), .A2(G233gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G127gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G183gat), .B(G211gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n226), .B(G127gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n229), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT16), .ZN(new_n235));
  INV_X1    g034(.A(G1gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT88), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT88), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G1gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n235), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n240), .B(KEYINPUT89), .ZN(new_n241));
  XNOR2_X1  g040(.A(G15gat), .B(G22gat), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n242), .A2(KEYINPUT87), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(KEYINPUT87), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n243), .A2(new_n236), .A3(new_n244), .ZN(new_n247));
  XOR2_X1   g046(.A(KEYINPUT90), .B(G8gat), .Z(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT91), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT91), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n246), .A2(new_n251), .A3(new_n247), .A4(new_n248), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n246), .A2(new_n247), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G8gat), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n250), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n255), .B1(new_n223), .B2(new_n222), .ZN(new_n256));
  OR2_X1    g055(.A1(new_n256), .A2(KEYINPUT100), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(KEYINPUT100), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n259));
  INV_X1    g058(.A(G155gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n257), .A2(new_n258), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n262), .B1(new_n257), .B2(new_n258), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n234), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n263), .A2(new_n264), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n267), .A2(new_n230), .A3(new_n233), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G85gat), .A2(G92gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT7), .ZN(new_n271));
  NAND2_X1  g070(.A1(G99gat), .A2(G106gat), .ZN(new_n272));
  INV_X1    g071(.A(G85gat), .ZN(new_n273));
  INV_X1    g072(.A(G92gat), .ZN(new_n274));
  AOI22_X1  g073(.A1(KEYINPUT8), .A2(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G99gat), .B(G106gat), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n276), .B(new_n277), .Z(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(G43gat), .B(G50gat), .Z(new_n280));
  INV_X1    g079(.A(KEYINPUT15), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(G29gat), .A2(G36gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT14), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G43gat), .B(G50gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT15), .ZN(new_n287));
  NAND2_X1  g086(.A1(G29gat), .A2(G36gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(KEYINPUT86), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n282), .A2(new_n285), .A3(new_n287), .A4(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  AOI211_X1 g090(.A(new_n281), .B(new_n280), .C1(new_n285), .C2(new_n289), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(G232gat), .A2(G233gat), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n279), .A2(new_n294), .B1(KEYINPUT41), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT17), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(new_n291), .B2(new_n292), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n289), .A3(new_n285), .ZN(new_n299));
  INV_X1    g098(.A(new_n287), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(KEYINPUT17), .A3(new_n290), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n296), .B1(new_n303), .B2(new_n279), .ZN(new_n304));
  XOR2_X1   g103(.A(G134gat), .B(G162gat), .Z(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(G190gat), .B(G218gat), .Z(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT102), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n295), .A2(KEYINPUT41), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(KEYINPUT101), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n308), .B(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n306), .B(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G230gat), .A2(G233gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(KEYINPUT105), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n221), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n317), .B1(new_n215), .B2(new_n217), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n271), .A2(new_n277), .A3(new_n275), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT103), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n278), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n318), .A2(new_n278), .A3(new_n321), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT10), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT10), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n278), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n318), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT104), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT104), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n318), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n316), .B1(new_n325), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G120gat), .B(G148gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(G176gat), .B(G204gat), .ZN(new_n335));
  XOR2_X1   g134(.A(new_n334), .B(new_n335), .Z(new_n336));
  NAND2_X1  g135(.A1(new_n323), .A2(new_n324), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n333), .B(new_n336), .C1(new_n337), .C2(new_n316), .ZN(new_n338));
  INV_X1    g137(.A(new_n336), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n329), .A2(new_n331), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n318), .A2(new_n278), .A3(new_n321), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n326), .B1(new_n341), .B2(new_n322), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n315), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n337), .A2(new_n316), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n339), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n338), .A2(new_n345), .ZN(new_n346));
  NOR3_X1   g145(.A1(new_n269), .A2(new_n313), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT95), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT71), .ZN(new_n350));
  NOR2_X1   g149(.A1(G169gat), .A2(G176gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(KEYINPUT67), .A3(KEYINPUT26), .ZN(new_n352));
  NAND2_X1  g151(.A1(G183gat), .A2(G190gat), .ZN(new_n353));
  INV_X1    g152(.A(G169gat), .ZN(new_n354));
  INV_X1    g153(.A(G176gat), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n354), .A2(new_n355), .A3(KEYINPUT67), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT26), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n357), .B1(new_n354), .B2(new_n355), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n352), .B(new_n353), .C1(new_n356), .C2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G183gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT27), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT27), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G183gat), .ZN(new_n363));
  INV_X1    g162(.A(G190gat), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n361), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT65), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT66), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT28), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT66), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n368), .B1(new_n365), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n359), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n366), .A2(KEYINPUT66), .A3(new_n368), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT23), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n373), .A2(G169gat), .A3(G176gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n351), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT23), .B1(new_n354), .B2(new_n355), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(G190gat), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n364), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n379), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT64), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n377), .B(new_n383), .C1(new_n384), .C2(KEYINPUT25), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n351), .A2(KEYINPUT23), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n373), .B1(G169gat), .B2(G176gat), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n384), .B(new_n386), .C1(new_n387), .C2(new_n351), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT25), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n386), .B1(new_n387), .B2(new_n351), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n364), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n378), .A2(G190gat), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n391), .B1(new_n392), .B2(new_n381), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n388), .B(new_n389), .C1(new_n390), .C2(new_n393), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n371), .A2(new_n372), .B1(new_n385), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G120gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(G113gat), .ZN(new_n397));
  INV_X1    g196(.A(G113gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(G120gat), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT1), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n227), .A2(G134gat), .ZN(new_n401));
  INV_X1    g200(.A(G134gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(G127gat), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT68), .B1(new_n227), .B2(G134gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n401), .A2(new_n403), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n406), .B1(new_n407), .B2(KEYINPUT68), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n405), .B1(new_n408), .B2(new_n400), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n395), .A2(KEYINPUT69), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n359), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n365), .A2(new_n369), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT28), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n369), .B1(new_n365), .B2(KEYINPUT65), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n372), .B(new_n411), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n394), .A2(new_n385), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OR2_X1    g216(.A1(new_n409), .A2(KEYINPUT69), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n409), .A2(KEYINPUT69), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G227gat), .ZN(new_n421));
  INV_X1    g220(.A(G233gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n410), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT32), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT33), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  XOR2_X1   g226(.A(G15gat), .B(G43gat), .Z(new_n428));
  XNOR2_X1  g227(.A(G71gat), .B(G99gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n425), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n430), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n424), .B(KEYINPUT32), .C1(new_n426), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n423), .B1(new_n410), .B2(new_n420), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT34), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI211_X1 g236(.A(KEYINPUT34), .B(new_n423), .C1(new_n410), .C2(new_n420), .ZN(new_n438));
  OR2_X1    g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n350), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n437), .A2(new_n438), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n441), .A2(new_n431), .A3(KEYINPUT71), .A4(new_n433), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n434), .A2(new_n439), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n445), .A2(KEYINPUT36), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT36), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n434), .A2(KEYINPUT70), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT70), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n431), .A2(new_n449), .A3(new_n433), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n439), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n447), .B1(new_n443), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n446), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT76), .ZN(new_n454));
  INV_X1    g253(.A(G148gat), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n454), .B1(new_n455), .B2(G141gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(G141gat), .ZN(new_n457));
  INV_X1    g256(.A(G141gat), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n458), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n456), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(G155gat), .A2(G162gat), .ZN(new_n461));
  INV_X1    g260(.A(G162gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n260), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n463), .B2(KEYINPUT2), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g264(.A1(G155gat), .A2(G162gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(G155gat), .A2(G162gat), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G141gat), .B(G148gat), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n468), .B1(new_n469), .B2(KEYINPUT2), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(G211gat), .ZN(new_n472));
  INV_X1    g271(.A(G218gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(G197gat), .ZN(new_n475));
  INV_X1    g274(.A(G204gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(G197gat), .A2(G204gat), .ZN(new_n478));
  OAI22_X1  g277(.A1(KEYINPUT22), .A2(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(G211gat), .B(G218gat), .Z(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT29), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  OAI221_X1 g281(.A(new_n480), .B1(KEYINPUT22), .B2(new_n474), .C1(new_n478), .C2(new_n477), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT80), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT3), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n484), .B1(new_n482), .B2(new_n483), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n471), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G228gat), .A2(G233gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n479), .A2(KEYINPUT72), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n480), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT72), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n465), .A2(new_n470), .A3(new_n486), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT77), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT77), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n465), .A2(new_n470), .A3(new_n498), .A4(new_n486), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT29), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n489), .B(new_n490), .C1(new_n495), .C2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n495), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT2), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n455), .A2(G141gat), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n458), .A2(G148gat), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n506), .A2(new_n468), .B1(new_n460), .B2(new_n464), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT29), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n508), .A3(new_n493), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n507), .B1(new_n509), .B2(new_n486), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n502), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n501), .B1(new_n511), .B2(new_n490), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT31), .B(G50gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G78gat), .B(G106gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(G22gat), .ZN(new_n516));
  INV_X1    g315(.A(new_n513), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n501), .B(new_n517), .C1(new_n490), .C2(new_n511), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n514), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n516), .B1(new_n514), .B2(new_n518), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n497), .A2(new_n499), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT68), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n523), .B1(new_n401), .B2(new_n403), .ZN(new_n524));
  XNOR2_X1  g323(.A(G113gat), .B(G120gat), .ZN(new_n525));
  OAI22_X1  g324(.A1(new_n524), .A2(new_n406), .B1(KEYINPUT1), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n471), .A2(KEYINPUT3), .B1(new_n526), .B2(new_n405), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT4), .B1(new_n409), .B2(new_n471), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT4), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n507), .A2(new_n529), .A3(new_n526), .A4(new_n405), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n522), .A2(new_n527), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G225gat), .A2(G233gat), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n409), .A2(new_n471), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n507), .A2(new_n526), .A3(new_n405), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n535), .A3(new_n532), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n536), .A2(KEYINPUT82), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(KEYINPUT82), .ZN(new_n538));
  AND4_X1   g337(.A1(KEYINPUT39), .A2(new_n533), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G1gat), .B(G29gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT0), .ZN(new_n541));
  XNOR2_X1  g340(.A(G57gat), .B(G85gat), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n541), .B(new_n542), .Z(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(new_n533), .B2(KEYINPUT39), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT81), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT81), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n546), .B(new_n543), .C1(new_n533), .C2(KEYINPUT39), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n539), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n548), .A2(KEYINPUT40), .ZN(new_n549));
  NAND2_X1  g348(.A1(G226gat), .A2(G233gat), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n550), .B(KEYINPUT73), .Z(new_n551));
  AOI21_X1  g350(.A(new_n551), .B1(new_n417), .B2(new_n508), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n550), .B1(new_n415), .B2(new_n416), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n494), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT74), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G8gat), .B(G36gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(G64gat), .B(G92gat), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n557), .B(new_n558), .Z(new_n559));
  OAI211_X1 g358(.A(KEYINPUT74), .B(new_n494), .C1(new_n552), .C2(new_n553), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n417), .A2(new_n508), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n550), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n417), .A2(new_n551), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n495), .A3(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n556), .A2(new_n559), .A3(new_n560), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT30), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n561), .A2(new_n550), .B1(new_n551), .B2(new_n417), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n554), .A2(new_n555), .B1(new_n567), .B2(new_n495), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT30), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n568), .A2(new_n569), .A3(new_n559), .A4(new_n560), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT75), .ZN(new_n572));
  INV_X1    g371(.A(new_n551), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(new_n395), .B2(KEYINPUT29), .ZN(new_n574));
  INV_X1    g373(.A(new_n553), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n495), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n564), .B1(new_n576), .B2(KEYINPUT74), .ZN(new_n577));
  INV_X1    g376(.A(new_n560), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n572), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n559), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n568), .A2(KEYINPUT75), .A3(new_n560), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n571), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n498), .B1(new_n507), .B2(new_n486), .ZN(new_n584));
  INV_X1    g383(.A(new_n499), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n527), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n528), .A2(new_n530), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT5), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n586), .A2(new_n587), .A3(new_n588), .A4(new_n532), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT78), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n531), .A2(KEYINPUT78), .A3(new_n588), .A4(new_n532), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n531), .A2(new_n532), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n534), .A2(new_n535), .ZN(new_n595));
  INV_X1    g394(.A(new_n532), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n588), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n543), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n548), .A2(KEYINPUT40), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n549), .A2(new_n583), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  OR3_X1    g402(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT37), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n604), .A2(KEYINPUT38), .A3(new_n580), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n579), .A2(KEYINPUT37), .A3(new_n581), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n567), .A2(new_n494), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n495), .B1(new_n552), .B2(new_n553), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n607), .A2(KEYINPUT37), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n604), .A2(new_n580), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT38), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n605), .A2(new_n606), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n591), .A2(new_n592), .B1(new_n594), .B2(new_n597), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT6), .B1(new_n613), .B2(new_n543), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n601), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n599), .A2(KEYINPUT6), .A3(new_n600), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n565), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n521), .B(new_n603), .C1(new_n612), .C2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n593), .A2(new_n598), .A3(new_n543), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT6), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n613), .A2(new_n543), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n616), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n582), .B(new_n571), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT79), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n521), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n617), .A2(KEYINPUT79), .A3(new_n582), .A4(new_n571), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n453), .A2(new_n620), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NOR4_X1   g433(.A1(new_n445), .A2(new_n627), .A3(new_n630), .A4(KEYINPUT35), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n443), .A2(new_n521), .A3(new_n451), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n571), .A2(new_n582), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT79), .B1(new_n638), .B2(new_n617), .ZN(new_n639));
  INV_X1    g438(.A(new_n631), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT35), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n635), .B1(new_n642), .B2(KEYINPUT83), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT83), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n641), .A2(new_n644), .A3(KEYINPUT35), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n634), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G113gat), .B(G141gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(G169gat), .B(G197gat), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT12), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT85), .ZN(new_n653));
  NAND2_X1  g452(.A1(G229gat), .A2(G233gat), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n250), .A2(new_n252), .A3(new_n254), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n294), .ZN(new_n657));
  INV_X1    g456(.A(new_n303), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n658), .A2(new_n252), .A3(new_n254), .A4(new_n250), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT92), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n255), .A2(KEYINPUT92), .A3(new_n658), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n655), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(KEYINPUT18), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n656), .B(new_n293), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(new_n654), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n663), .A2(KEYINPUT18), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n653), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n668), .B1(KEYINPUT18), .B2(new_n663), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT94), .B1(new_n663), .B2(KEYINPUT18), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT94), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT18), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n656), .A2(new_n660), .A3(new_n303), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT92), .B1(new_n656), .B2(new_n294), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n677), .B1(new_n659), .B2(new_n678), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n675), .B(new_n676), .C1(new_n679), .C2(new_n655), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n673), .A2(new_n674), .A3(new_n652), .A4(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n672), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n349), .B1(new_n646), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n636), .B1(new_n629), .B2(new_n631), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT35), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT83), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n635), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n645), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n633), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(KEYINPUT95), .A3(new_n682), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n348), .B1(new_n684), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n618), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g493(.A(KEYINPUT16), .B(G8gat), .Z(new_n695));
  NAND4_X1  g494(.A1(new_n692), .A2(KEYINPUT42), .A3(new_n583), .A4(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT95), .B1(new_n690), .B2(new_n682), .ZN(new_n698));
  AOI211_X1 g497(.A(new_n349), .B(new_n683), .C1(new_n689), .C2(new_n633), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n583), .B(new_n347), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n695), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n697), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(G8gat), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n696), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT106), .ZN(G1325gat));
  INV_X1    g504(.A(new_n445), .ZN(new_n706));
  AOI21_X1  g505(.A(G15gat), .B1(new_n692), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n453), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G15gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT107), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n707), .B1(new_n692), .B2(new_n710), .ZN(G1326gat));
  NAND2_X1  g510(.A1(new_n692), .A2(new_n630), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT43), .B(G22gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1327gat));
  NAND2_X1  g513(.A1(new_n684), .A2(new_n691), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n346), .B1(new_n266), .B2(new_n268), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n716), .A2(new_n313), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(G29gat), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n719), .A2(new_n720), .A3(new_n618), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT45), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT44), .B1(new_n690), .B2(new_n313), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n725));
  AOI211_X1 g524(.A(new_n725), .B(new_n312), .C1(new_n689), .C2(new_n633), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT108), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n682), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n672), .A2(new_n681), .A3(KEYINPUT108), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n716), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT109), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n727), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(G29gat), .B1(new_n735), .B2(new_n617), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n722), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n723), .A2(new_n736), .A3(new_n737), .ZN(G1328gat));
  INV_X1    g537(.A(G36gat), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n719), .A2(new_n739), .A3(new_n583), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n740), .A2(KEYINPUT46), .ZN(new_n741));
  OAI21_X1  g540(.A(G36gat), .B1(new_n735), .B2(new_n638), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(KEYINPUT46), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(G1329gat));
  OAI21_X1  g543(.A(G43gat), .B1(new_n735), .B2(new_n453), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT47), .B1(new_n745), .B2(KEYINPUT110), .ZN(new_n746));
  OR2_X1    g545(.A1(new_n445), .A2(G43gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n718), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  OAI221_X1 g548(.A(new_n745), .B1(KEYINPUT110), .B2(KEYINPUT47), .C1(new_n718), .C2(new_n747), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(G1330gat));
  OAI21_X1  g550(.A(new_n725), .B1(new_n646), .B2(new_n312), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n312), .B1(new_n689), .B2(new_n633), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT44), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n752), .A2(new_n630), .A3(new_n754), .A4(new_n734), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT111), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n727), .A2(new_n757), .A3(new_n630), .A4(new_n734), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n756), .A2(new_n758), .A3(G50gat), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n521), .A2(G50gat), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n717), .B(new_n760), .C1(new_n698), .C2(new_n699), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT48), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n755), .A2(G50gat), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n761), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT48), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n764), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(G50gat), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n755), .B2(KEYINPUT111), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n762), .B1(new_n772), .B2(new_n758), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT48), .B1(new_n765), .B2(new_n761), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT112), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n770), .A2(new_n775), .ZN(G1331gat));
  INV_X1    g575(.A(new_n269), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n312), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n731), .A2(new_n346), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n646), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n618), .ZN(new_n781));
  XOR2_X1   g580(.A(KEYINPUT113), .B(G57gat), .Z(new_n782));
  XNOR2_X1  g581(.A(new_n781), .B(new_n782), .ZN(G1332gat));
  XNOR2_X1  g582(.A(new_n583), .B(KEYINPUT114), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n786));
  AND2_X1   g585(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(new_n785), .B2(new_n786), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT115), .ZN(G1333gat));
  NAND2_X1  g589(.A1(new_n780), .A2(new_n708), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n445), .A2(G71gat), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n791), .A2(G71gat), .B1(new_n780), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n793), .B(new_n794), .ZN(G1334gat));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n630), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G78gat), .ZN(G1335gat));
  INV_X1    g596(.A(new_n346), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n798), .A2(G85gat), .A3(new_n617), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n732), .A2(new_n777), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n690), .A2(new_n313), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT117), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n753), .A2(KEYINPUT51), .A3(new_n800), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT117), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n805), .A2(new_n807), .A3(KEYINPUT118), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n799), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n779), .A2(new_n777), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n727), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(G85gat), .B1(new_n814), .B2(new_n617), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n815), .ZN(G1336gat));
  AND2_X1   g615(.A1(new_n727), .A2(new_n813), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n583), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n806), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n784), .A2(new_n274), .A3(new_n346), .ZN(new_n820));
  XOR2_X1   g619(.A(new_n820), .B(KEYINPUT119), .Z(new_n821));
  AOI22_X1  g620(.A1(new_n818), .A2(G92gat), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n820), .ZN(new_n824));
  INV_X1    g623(.A(new_n784), .ZN(new_n825));
  OAI21_X1  g624(.A(G92gat), .B1(new_n814), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n823), .ZN(new_n827));
  OAI22_X1  g626(.A1(new_n822), .A2(new_n823), .B1(new_n824), .B2(new_n827), .ZN(G1337gat));
  NOR3_X1   g627(.A1(new_n798), .A2(new_n445), .A3(G99gat), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n810), .B2(new_n811), .ZN(new_n830));
  OAI21_X1  g629(.A(G99gat), .B1(new_n814), .B2(new_n453), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(G1338gat));
  NAND3_X1  g631(.A1(new_n727), .A2(new_n630), .A3(new_n813), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n833), .A2(G106gat), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n798), .A2(G106gat), .A3(new_n521), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n803), .B2(new_n806), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT53), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n819), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n836), .B1(new_n840), .B2(new_n804), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(KEYINPUT120), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT53), .B1(new_n833), .B2(G106gat), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n843), .B1(new_n841), .B2(KEYINPUT120), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n838), .B1(new_n842), .B2(new_n844), .ZN(G1339gat));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n336), .B1(new_n343), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n340), .A2(new_n342), .A3(new_n315), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n333), .A2(new_n848), .A3(KEYINPUT54), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n847), .A2(new_n849), .A3(KEYINPUT55), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n852), .A2(new_n338), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n729), .A2(new_n854), .A3(new_n730), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n661), .A2(new_n662), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT121), .B1(new_n856), .B2(new_n654), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n665), .A2(new_n667), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT122), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT122), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n665), .A2(new_n860), .A3(new_n667), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n857), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n856), .A2(KEYINPUT121), .A3(new_n654), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n651), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n681), .A3(new_n346), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n313), .B1(new_n855), .B2(new_n865), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n864), .A2(new_n681), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n854), .A2(new_n867), .A3(new_n313), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n269), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n347), .A2(new_n731), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n445), .A2(new_n630), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n784), .A2(new_n617), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(new_n398), .A3(new_n683), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n617), .B1(new_n869), .B2(new_n870), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n877), .A2(new_n637), .A3(new_n825), .ZN(new_n878));
  AOI21_X1  g677(.A(G113gat), .B1(new_n878), .B2(new_n732), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n876), .A2(new_n879), .ZN(G1340gat));
  OAI21_X1  g679(.A(G120gat), .B1(new_n875), .B2(new_n798), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n346), .A2(new_n396), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n882), .B(KEYINPUT123), .Z(new_n883));
  NAND2_X1  g682(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n881), .A2(new_n884), .ZN(G1341gat));
  OAI21_X1  g684(.A(G127gat), .B1(new_n875), .B2(new_n269), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n878), .A2(new_n227), .A3(new_n777), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1342gat));
  OAI21_X1  g687(.A(G134gat), .B1(new_n875), .B2(new_n312), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n312), .A2(new_n583), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n877), .A2(new_n402), .A3(new_n637), .A4(new_n890), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n891), .A2(KEYINPUT56), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(KEYINPUT56), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n889), .A2(new_n892), .A3(new_n893), .ZN(G1343gat));
  INV_X1    g693(.A(KEYINPUT126), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT58), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n874), .A2(new_n453), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n852), .A2(new_n338), .A3(new_n853), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n865), .B1(new_n683), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n312), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n854), .A2(new_n867), .A3(new_n313), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n777), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n347), .A2(new_n731), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n630), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n897), .B1(new_n904), .B2(KEYINPUT57), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT57), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n871), .A2(new_n906), .A3(new_n630), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n905), .A2(new_n907), .A3(new_n682), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT58), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n909), .A3(G141gat), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n708), .A2(new_n521), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n911), .B1(new_n877), .B2(KEYINPUT125), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n913));
  AOI211_X1 g712(.A(new_n913), .B(new_n617), .C1(new_n869), .C2(new_n870), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n825), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n683), .A2(G141gat), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n896), .B(new_n910), .C1(new_n916), .C2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n920));
  AOI211_X1 g719(.A(KEYINPUT57), .B(new_n521), .C1(new_n869), .C2(new_n870), .ZN(new_n921));
  INV_X1    g720(.A(new_n897), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n682), .A2(new_n338), .A3(new_n852), .A4(new_n853), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n313), .B1(new_n923), .B2(new_n865), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n269), .B1(new_n924), .B2(new_n868), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n521), .B1(new_n925), .B2(new_n870), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n922), .B1(new_n926), .B2(new_n906), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n920), .B1(new_n921), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n905), .A2(new_n907), .A3(KEYINPUT124), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(new_n929), .A3(new_n732), .ZN(new_n930));
  NOR4_X1   g729(.A1(new_n912), .A2(new_n914), .A3(new_n784), .A4(new_n918), .ZN(new_n931));
  AOI22_X1  g730(.A1(G141gat), .A2(new_n930), .B1(new_n931), .B2(new_n895), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n919), .B1(new_n932), .B2(new_n909), .ZN(G1344gat));
  NAND3_X1  g732(.A1(new_n928), .A2(new_n929), .A3(new_n346), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n455), .A2(KEYINPUT59), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n925), .B1(new_n682), .B2(new_n348), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(new_n906), .A3(new_n630), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n521), .B1(new_n869), .B2(new_n870), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n938), .B(new_n346), .C1(new_n939), .C2(new_n906), .ZN(new_n940));
  OAI21_X1  g739(.A(G148gat), .B1(new_n940), .B2(new_n897), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n941), .A2(KEYINPUT59), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n346), .A2(new_n455), .ZN(new_n943));
  OAI22_X1  g742(.A1(new_n936), .A2(new_n942), .B1(new_n916), .B2(new_n943), .ZN(G1345gat));
  AND3_X1   g743(.A1(new_n928), .A2(new_n929), .A3(new_n777), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n777), .A2(new_n260), .ZN(new_n946));
  OAI22_X1  g745(.A1(new_n945), .A2(new_n260), .B1(new_n916), .B2(new_n946), .ZN(G1346gat));
  NAND3_X1  g746(.A1(new_n915), .A2(new_n462), .A3(new_n890), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n928), .A2(new_n929), .A3(new_n313), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(new_n462), .ZN(G1347gat));
  NOR2_X1   g749(.A1(new_n638), .A2(new_n618), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n873), .A2(new_n951), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n952), .A2(new_n354), .A3(new_n683), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n825), .A2(new_n618), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n871), .A2(new_n637), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(G169gat), .B1(new_n955), .B2(new_n732), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n953), .A2(new_n956), .ZN(G1348gat));
  OAI21_X1  g756(.A(G176gat), .B1(new_n952), .B2(new_n798), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n955), .A2(new_n355), .A3(new_n346), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1349gat));
  OAI21_X1  g759(.A(G183gat), .B1(new_n952), .B2(new_n269), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n777), .A2(new_n361), .A3(new_n363), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n962), .B1(new_n955), .B2(new_n963), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n955), .A2(new_n962), .A3(new_n963), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(KEYINPUT60), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT60), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n961), .B(new_n968), .C1(new_n964), .C2(new_n965), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(G1350gat));
  NAND3_X1  g769(.A1(new_n955), .A2(new_n364), .A3(new_n313), .ZN(new_n971));
  OAI21_X1  g770(.A(G190gat), .B1(new_n952), .B2(new_n312), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n972), .A2(KEYINPUT61), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n972), .A2(KEYINPUT61), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(G1351gat));
  OR2_X1    g774(.A1(new_n939), .A2(new_n906), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n453), .A2(new_n951), .ZN(new_n977));
  INV_X1    g776(.A(new_n977), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n976), .A2(new_n938), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n682), .A2(G197gat), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n871), .A2(new_n911), .A3(new_n954), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n981), .A2(new_n732), .ZN(new_n982));
  OAI22_X1  g781(.A1(new_n979), .A2(new_n980), .B1(new_n982), .B2(G197gat), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(G1352gat));
  NAND3_X1  g783(.A1(new_n981), .A2(new_n476), .A3(new_n346), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n986));
  OAI21_X1  g785(.A(G204gat), .B1(new_n940), .B2(new_n977), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(G1353gat));
  NAND3_X1  g788(.A1(new_n981), .A2(new_n472), .A3(new_n777), .ZN(new_n990));
  NAND4_X1  g789(.A1(new_n976), .A2(new_n777), .A3(new_n938), .A4(new_n978), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n991), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n992));
  INV_X1    g791(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g792(.A(KEYINPUT63), .B1(new_n991), .B2(G211gat), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n990), .B1(new_n993), .B2(new_n994), .ZN(G1354gat));
  OAI21_X1  g794(.A(G218gat), .B1(new_n979), .B2(new_n312), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n981), .A2(new_n473), .A3(new_n313), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n996), .A2(new_n997), .ZN(G1355gat));
endmodule


