

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U551 ( .A(KEYINPUT65), .ZN(n556) );
  NOR2_X1 U552 ( .A1(n806), .A2(n517), .ZN(n516) );
  AND2_X1 U553 ( .A1(n978), .A2(n817), .ZN(n517) );
  OR2_X1 U554 ( .A1(n771), .A2(n770), .ZN(n518) );
  NAND2_X1 U555 ( .A1(n685), .A2(n773), .ZN(n691) );
  OR2_X1 U556 ( .A1(n893), .A2(n697), .ZN(n695) );
  INV_X1 U557 ( .A(KEYINPUT98), .ZN(n700) );
  XNOR2_X1 U558 ( .A(n701), .B(n700), .ZN(n707) );
  INV_X1 U559 ( .A(KEYINPUT29), .ZN(n713) );
  XNOR2_X1 U560 ( .A(n740), .B(KEYINPUT100), .ZN(n741) );
  NAND2_X1 U561 ( .A1(n741), .A2(G8), .ZN(n743) );
  XNOR2_X1 U562 ( .A(n743), .B(n742), .ZN(n756) );
  XNOR2_X1 U563 ( .A(G2104), .B(KEYINPUT64), .ZN(n559) );
  NAND2_X1 U564 ( .A1(n882), .A2(G101), .ZN(n558) );
  XNOR2_X1 U565 ( .A(KEYINPUT66), .B(n553), .ZN(n883) );
  NOR2_X1 U566 ( .A1(G651), .A2(n643), .ZN(n636) );
  AND2_X1 U567 ( .A1(n562), .A2(n561), .ZN(n684) );
  NOR2_X1 U568 ( .A1(G651), .A2(G543), .ZN(n627) );
  NAND2_X1 U569 ( .A1(n627), .A2(G89), .ZN(n519) );
  XNOR2_X1 U570 ( .A(n519), .B(KEYINPUT4), .ZN(n521) );
  XOR2_X1 U571 ( .A(KEYINPUT0), .B(G543), .Z(n643) );
  INV_X1 U572 ( .A(G651), .ZN(n523) );
  NOR2_X1 U573 ( .A1(n643), .A2(n523), .ZN(n630) );
  NAND2_X1 U574 ( .A1(G76), .A2(n630), .ZN(n520) );
  NAND2_X1 U575 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U576 ( .A(n522), .B(KEYINPUT5), .ZN(n530) );
  NOR2_X1 U577 ( .A1(G543), .A2(n523), .ZN(n524) );
  XOR2_X1 U578 ( .A(KEYINPUT1), .B(n524), .Z(n642) );
  NAND2_X1 U579 ( .A1(n642), .A2(G63), .ZN(n525) );
  XNOR2_X1 U580 ( .A(n525), .B(KEYINPUT74), .ZN(n527) );
  NAND2_X1 U581 ( .A1(G51), .A2(n636), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U583 ( .A(KEYINPUT6), .B(n528), .Z(n529) );
  NAND2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U585 ( .A(n531), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U586 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U587 ( .A1(G85), .A2(n627), .ZN(n533) );
  NAND2_X1 U588 ( .A1(G72), .A2(n630), .ZN(n532) );
  NAND2_X1 U589 ( .A1(n533), .A2(n532), .ZN(n537) );
  NAND2_X1 U590 ( .A1(G60), .A2(n642), .ZN(n535) );
  NAND2_X1 U591 ( .A1(G47), .A2(n636), .ZN(n534) );
  NAND2_X1 U592 ( .A1(n535), .A2(n534), .ZN(n536) );
  OR2_X1 U593 ( .A1(n537), .A2(n536), .ZN(G290) );
  NAND2_X1 U594 ( .A1(G64), .A2(n642), .ZN(n539) );
  NAND2_X1 U595 ( .A1(G52), .A2(n636), .ZN(n538) );
  NAND2_X1 U596 ( .A1(n539), .A2(n538), .ZN(n544) );
  NAND2_X1 U597 ( .A1(G90), .A2(n627), .ZN(n541) );
  NAND2_X1 U598 ( .A1(G77), .A2(n630), .ZN(n540) );
  NAND2_X1 U599 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(n542), .Z(n543) );
  NOR2_X1 U601 ( .A1(n544), .A2(n543), .ZN(G171) );
  AND2_X1 U602 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U603 ( .A(G82), .ZN(G220) );
  INV_X1 U604 ( .A(G57), .ZN(G237) );
  INV_X1 U605 ( .A(G69), .ZN(G235) );
  INV_X1 U606 ( .A(G108), .ZN(G238) );
  INV_X1 U607 ( .A(G120), .ZN(G236) );
  NAND2_X1 U608 ( .A1(G65), .A2(n642), .ZN(n546) );
  NAND2_X1 U609 ( .A1(G53), .A2(n636), .ZN(n545) );
  NAND2_X1 U610 ( .A1(n546), .A2(n545), .ZN(n550) );
  NAND2_X1 U611 ( .A1(G91), .A2(n627), .ZN(n548) );
  NAND2_X1 U612 ( .A1(G78), .A2(n630), .ZN(n547) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U614 ( .A1(n550), .A2(n549), .ZN(n708) );
  INV_X1 U615 ( .A(n708), .ZN(G299) );
  XNOR2_X1 U616 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n552) );
  NOR2_X1 U617 ( .A1(G2105), .A2(G2104), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  NAND2_X1 U619 ( .A1(G137), .A2(n883), .ZN(n555) );
  AND2_X1 U620 ( .A1(G2105), .A2(G2104), .ZN(n879) );
  NAND2_X1 U621 ( .A1(n879), .A2(G113), .ZN(n554) );
  NAND2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n682) );
  INV_X1 U623 ( .A(G2105), .ZN(n560) );
  AND2_X1 U624 ( .A1(n559), .A2(n560), .ZN(n557) );
  XNOR2_X2 U625 ( .A(n557), .B(n556), .ZN(n882) );
  XOR2_X1 U626 ( .A(KEYINPUT23), .B(n558), .Z(n562) );
  NOR2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n878) );
  NAND2_X1 U628 ( .A1(n878), .A2(G125), .ZN(n561) );
  INV_X1 U629 ( .A(n684), .ZN(n563) );
  NOR2_X1 U630 ( .A1(n682), .A2(n563), .ZN(G160) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U633 ( .A(G223), .ZN(n822) );
  NAND2_X1 U634 ( .A1(n822), .A2(G567), .ZN(n565) );
  XOR2_X1 U635 ( .A(KEYINPUT11), .B(n565), .Z(G234) );
  XNOR2_X1 U636 ( .A(KEYINPUT13), .B(KEYINPUT71), .ZN(n571) );
  NAND2_X1 U637 ( .A1(G81), .A2(n627), .ZN(n566) );
  XNOR2_X1 U638 ( .A(n566), .B(KEYINPUT70), .ZN(n567) );
  XNOR2_X1 U639 ( .A(n567), .B(KEYINPUT12), .ZN(n569) );
  NAND2_X1 U640 ( .A1(G68), .A2(n630), .ZN(n568) );
  NAND2_X1 U641 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U642 ( .A(n571), .B(n570), .ZN(n575) );
  NAND2_X1 U643 ( .A1(G56), .A2(n642), .ZN(n572) );
  XNOR2_X1 U644 ( .A(n572), .B(KEYINPUT69), .ZN(n573) );
  XNOR2_X1 U645 ( .A(n573), .B(KEYINPUT14), .ZN(n574) );
  NOR2_X1 U646 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U647 ( .A1(n636), .A2(G43), .ZN(n576) );
  NAND2_X1 U648 ( .A1(n577), .A2(n576), .ZN(n981) );
  INV_X1 U649 ( .A(G860), .ZN(n592) );
  OR2_X1 U650 ( .A1(n981), .A2(n592), .ZN(G153) );
  INV_X1 U651 ( .A(G171), .ZN(G301) );
  NAND2_X1 U652 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U653 ( .A1(G92), .A2(n627), .ZN(n578) );
  XNOR2_X1 U654 ( .A(n578), .B(KEYINPUT72), .ZN(n585) );
  NAND2_X1 U655 ( .A1(G79), .A2(n630), .ZN(n580) );
  NAND2_X1 U656 ( .A1(G66), .A2(n642), .ZN(n579) );
  NAND2_X1 U657 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U658 ( .A1(G54), .A2(n636), .ZN(n581) );
  XNOR2_X1 U659 ( .A(KEYINPUT73), .B(n581), .ZN(n582) );
  NOR2_X1 U660 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U661 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U662 ( .A(KEYINPUT15), .B(n586), .ZN(n893) );
  INV_X1 U663 ( .A(n893), .ZN(n965) );
  INV_X1 U664 ( .A(G868), .ZN(n589) );
  NAND2_X1 U665 ( .A1(n965), .A2(n589), .ZN(n587) );
  NAND2_X1 U666 ( .A1(n588), .A2(n587), .ZN(G284) );
  NOR2_X1 U667 ( .A1(G286), .A2(n589), .ZN(n591) );
  NOR2_X1 U668 ( .A1(G868), .A2(G299), .ZN(n590) );
  NOR2_X1 U669 ( .A1(n591), .A2(n590), .ZN(G297) );
  NAND2_X1 U670 ( .A1(n592), .A2(G559), .ZN(n593) );
  NAND2_X1 U671 ( .A1(n593), .A2(n893), .ZN(n594) );
  XNOR2_X1 U672 ( .A(n594), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U673 ( .A1(G868), .A2(n981), .ZN(n595) );
  XOR2_X1 U674 ( .A(KEYINPUT75), .B(n595), .Z(n599) );
  NAND2_X1 U675 ( .A1(n893), .A2(G868), .ZN(n596) );
  NOR2_X1 U676 ( .A1(G559), .A2(n596), .ZN(n597) );
  XNOR2_X1 U677 ( .A(KEYINPUT76), .B(n597), .ZN(n598) );
  NOR2_X1 U678 ( .A1(n599), .A2(n598), .ZN(G282) );
  NAND2_X1 U679 ( .A1(G123), .A2(n878), .ZN(n600) );
  XOR2_X1 U680 ( .A(KEYINPUT18), .B(n600), .Z(n601) );
  XNOR2_X1 U681 ( .A(n601), .B(KEYINPUT77), .ZN(n603) );
  NAND2_X1 U682 ( .A1(G111), .A2(n879), .ZN(n602) );
  NAND2_X1 U683 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U684 ( .A1(n882), .A2(G99), .ZN(n605) );
  NAND2_X1 U685 ( .A1(G135), .A2(n883), .ZN(n604) );
  NAND2_X1 U686 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U687 ( .A1(n607), .A2(n606), .ZN(n922) );
  XNOR2_X1 U688 ( .A(n922), .B(G2096), .ZN(n608) );
  XNOR2_X1 U689 ( .A(n608), .B(KEYINPUT78), .ZN(n610) );
  INV_X1 U690 ( .A(G2100), .ZN(n609) );
  NAND2_X1 U691 ( .A1(n610), .A2(n609), .ZN(G156) );
  NAND2_X1 U692 ( .A1(n893), .A2(G559), .ZN(n654) );
  XNOR2_X1 U693 ( .A(n981), .B(n654), .ZN(n611) );
  NOR2_X1 U694 ( .A1(n611), .A2(G860), .ZN(n619) );
  NAND2_X1 U695 ( .A1(n642), .A2(G67), .ZN(n614) );
  NAND2_X1 U696 ( .A1(G93), .A2(n627), .ZN(n612) );
  XOR2_X1 U697 ( .A(KEYINPUT79), .B(n612), .Z(n613) );
  NAND2_X1 U698 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U699 ( .A1(G80), .A2(n630), .ZN(n616) );
  NAND2_X1 U700 ( .A1(G55), .A2(n636), .ZN(n615) );
  NAND2_X1 U701 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U702 ( .A1(n618), .A2(n617), .ZN(n651) );
  XNOR2_X1 U703 ( .A(n619), .B(n651), .ZN(G145) );
  NAND2_X1 U704 ( .A1(G88), .A2(n627), .ZN(n621) );
  NAND2_X1 U705 ( .A1(G75), .A2(n630), .ZN(n620) );
  NAND2_X1 U706 ( .A1(n621), .A2(n620), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n642), .A2(G62), .ZN(n622) );
  XNOR2_X1 U708 ( .A(n622), .B(KEYINPUT82), .ZN(n624) );
  NAND2_X1 U709 ( .A1(G50), .A2(n636), .ZN(n623) );
  NAND2_X1 U710 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U711 ( .A1(n626), .A2(n625), .ZN(G166) );
  NAND2_X1 U712 ( .A1(G86), .A2(n627), .ZN(n629) );
  NAND2_X1 U713 ( .A1(G61), .A2(n642), .ZN(n628) );
  NAND2_X1 U714 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U715 ( .A1(n630), .A2(G73), .ZN(n631) );
  XOR2_X1 U716 ( .A(KEYINPUT2), .B(n631), .Z(n632) );
  NOR2_X1 U717 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n636), .A2(G48), .ZN(n634) );
  NAND2_X1 U719 ( .A1(n635), .A2(n634), .ZN(G305) );
  NAND2_X1 U720 ( .A1(n636), .A2(G49), .ZN(n637) );
  XNOR2_X1 U721 ( .A(n637), .B(KEYINPUT80), .ZN(n639) );
  NAND2_X1 U722 ( .A1(G74), .A2(G651), .ZN(n638) );
  NAND2_X1 U723 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U724 ( .A(KEYINPUT81), .B(n640), .Z(n641) );
  NOR2_X1 U725 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n643), .A2(G87), .ZN(n644) );
  NAND2_X1 U727 ( .A1(n645), .A2(n644), .ZN(G288) );
  NOR2_X1 U728 ( .A1(G868), .A2(n651), .ZN(n646) );
  XNOR2_X1 U729 ( .A(n646), .B(KEYINPUT83), .ZN(n657) );
  XNOR2_X1 U730 ( .A(KEYINPUT19), .B(G299), .ZN(n647) );
  XNOR2_X1 U731 ( .A(n647), .B(n981), .ZN(n650) );
  XNOR2_X1 U732 ( .A(G166), .B(G305), .ZN(n648) );
  XNOR2_X1 U733 ( .A(n648), .B(G288), .ZN(n649) );
  XNOR2_X1 U734 ( .A(n650), .B(n649), .ZN(n653) );
  XNOR2_X1 U735 ( .A(G290), .B(n651), .ZN(n652) );
  XNOR2_X1 U736 ( .A(n653), .B(n652), .ZN(n894) );
  XOR2_X1 U737 ( .A(n894), .B(n654), .Z(n655) );
  NAND2_X1 U738 ( .A1(G868), .A2(n655), .ZN(n656) );
  NAND2_X1 U739 ( .A1(n657), .A2(n656), .ZN(G295) );
  NAND2_X1 U740 ( .A1(G2078), .A2(G2084), .ZN(n658) );
  XOR2_X1 U741 ( .A(KEYINPUT20), .B(n658), .Z(n659) );
  NAND2_X1 U742 ( .A1(G2090), .A2(n659), .ZN(n660) );
  XNOR2_X1 U743 ( .A(KEYINPUT21), .B(n660), .ZN(n661) );
  NAND2_X1 U744 ( .A1(n661), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U745 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U746 ( .A(KEYINPUT68), .B(G132), .Z(G219) );
  NOR2_X1 U747 ( .A1(G236), .A2(G238), .ZN(n663) );
  NOR2_X1 U748 ( .A1(G235), .A2(G237), .ZN(n662) );
  NAND2_X1 U749 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U750 ( .A(KEYINPUT84), .B(n664), .ZN(n827) );
  NAND2_X1 U751 ( .A1(n827), .A2(G567), .ZN(n665) );
  XOR2_X1 U752 ( .A(KEYINPUT85), .B(n665), .Z(n670) );
  NOR2_X1 U753 ( .A1(G219), .A2(G220), .ZN(n666) );
  XOR2_X1 U754 ( .A(KEYINPUT22), .B(n666), .Z(n667) );
  NOR2_X1 U755 ( .A1(G218), .A2(n667), .ZN(n668) );
  NAND2_X1 U756 ( .A1(G96), .A2(n668), .ZN(n826) );
  NAND2_X1 U757 ( .A1(G2106), .A2(n826), .ZN(n669) );
  NAND2_X1 U758 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U759 ( .A(KEYINPUT86), .B(n671), .Z(G319) );
  INV_X1 U760 ( .A(G319), .ZN(n673) );
  NAND2_X1 U761 ( .A1(G661), .A2(G483), .ZN(n672) );
  NOR2_X1 U762 ( .A1(n673), .A2(n672), .ZN(n825) );
  NAND2_X1 U763 ( .A1(n825), .A2(G36), .ZN(G176) );
  NAND2_X1 U764 ( .A1(n882), .A2(G102), .ZN(n675) );
  NAND2_X1 U765 ( .A1(G138), .A2(n883), .ZN(n674) );
  NAND2_X1 U766 ( .A1(n675), .A2(n674), .ZN(n679) );
  NAND2_X1 U767 ( .A1(G126), .A2(n878), .ZN(n677) );
  NAND2_X1 U768 ( .A1(G114), .A2(n879), .ZN(n676) );
  NAND2_X1 U769 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U770 ( .A1(n679), .A2(n678), .ZN(G164) );
  XNOR2_X1 U771 ( .A(KEYINPUT87), .B(G166), .ZN(G303) );
  NOR2_X1 U772 ( .A1(G1981), .A2(G305), .ZN(n680) );
  XNOR2_X1 U773 ( .A(KEYINPUT24), .B(n680), .ZN(n686) );
  INV_X1 U774 ( .A(G40), .ZN(n681) );
  NOR2_X1 U775 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U776 ( .A1(n684), .A2(n683), .ZN(n772) );
  XNOR2_X1 U777 ( .A(n772), .B(KEYINPUT95), .ZN(n685) );
  NOR2_X1 U778 ( .A1(G164), .A2(G1384), .ZN(n773) );
  NAND2_X1 U779 ( .A1(G8), .A2(n691), .ZN(n759) );
  INV_X1 U780 ( .A(n759), .ZN(n751) );
  NAND2_X1 U781 ( .A1(n686), .A2(n751), .ZN(n749) );
  NOR2_X1 U782 ( .A1(G2084), .A2(n691), .ZN(n719) );
  NAND2_X1 U783 ( .A1(G8), .A2(n719), .ZN(n733) );
  NOR2_X1 U784 ( .A1(G1966), .A2(n759), .ZN(n731) );
  AND2_X1 U785 ( .A1(n703), .A2(G1996), .ZN(n687) );
  XOR2_X1 U786 ( .A(n687), .B(KEYINPUT26), .Z(n690) );
  AND2_X1 U787 ( .A1(n691), .A2(G1341), .ZN(n688) );
  NOR2_X1 U788 ( .A1(n688), .A2(n981), .ZN(n689) );
  AND2_X1 U789 ( .A1(n690), .A2(n689), .ZN(n696) );
  NAND2_X1 U790 ( .A1(G1348), .A2(n691), .ZN(n693) );
  NAND2_X1 U791 ( .A1(n703), .A2(G2067), .ZN(n692) );
  NAND2_X1 U792 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U793 ( .A(n694), .B(KEYINPUT97), .ZN(n697) );
  NAND2_X1 U794 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U795 ( .A1(n697), .A2(n893), .ZN(n698) );
  NAND2_X1 U796 ( .A1(n699), .A2(n698), .ZN(n701) );
  INV_X1 U797 ( .A(n691), .ZN(n703) );
  NAND2_X1 U798 ( .A1(n703), .A2(G2072), .ZN(n702) );
  XNOR2_X1 U799 ( .A(n702), .B(KEYINPUT27), .ZN(n705) );
  XOR2_X1 U800 ( .A(KEYINPUT96), .B(G1956), .Z(n990) );
  NOR2_X1 U801 ( .A1(n703), .A2(n990), .ZN(n704) );
  NOR2_X1 U802 ( .A1(n705), .A2(n704), .ZN(n709) );
  NAND2_X1 U803 ( .A1(n709), .A2(n708), .ZN(n706) );
  NAND2_X1 U804 ( .A1(n707), .A2(n706), .ZN(n712) );
  NOR2_X1 U805 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U806 ( .A(n710), .B(KEYINPUT28), .Z(n711) );
  NAND2_X1 U807 ( .A1(n712), .A2(n711), .ZN(n714) );
  XNOR2_X1 U808 ( .A(n714), .B(n713), .ZN(n718) );
  XNOR2_X1 U809 ( .A(G2078), .B(KEYINPUT25), .ZN(n942) );
  NOR2_X1 U810 ( .A1(n691), .A2(n942), .ZN(n716) );
  AND2_X1 U811 ( .A1(n691), .A2(G1961), .ZN(n715) );
  NOR2_X1 U812 ( .A1(n716), .A2(n715), .ZN(n723) );
  NAND2_X1 U813 ( .A1(G171), .A2(n723), .ZN(n717) );
  NAND2_X1 U814 ( .A1(n718), .A2(n717), .ZN(n729) );
  NOR2_X1 U815 ( .A1(n731), .A2(n719), .ZN(n720) );
  NAND2_X1 U816 ( .A1(G8), .A2(n720), .ZN(n721) );
  XNOR2_X1 U817 ( .A(KEYINPUT30), .B(n721), .ZN(n722) );
  NOR2_X1 U818 ( .A1(G168), .A2(n722), .ZN(n725) );
  NOR2_X1 U819 ( .A1(G171), .A2(n723), .ZN(n724) );
  NOR2_X1 U820 ( .A1(n725), .A2(n724), .ZN(n727) );
  XNOR2_X1 U821 ( .A(KEYINPUT99), .B(KEYINPUT31), .ZN(n726) );
  XNOR2_X1 U822 ( .A(n727), .B(n726), .ZN(n728) );
  NAND2_X1 U823 ( .A1(n729), .A2(n728), .ZN(n734) );
  INV_X1 U824 ( .A(n734), .ZN(n730) );
  NOR2_X1 U825 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U826 ( .A1(n733), .A2(n732), .ZN(n754) );
  NAND2_X1 U827 ( .A1(n734), .A2(G286), .ZN(n739) );
  NOR2_X1 U828 ( .A1(G1971), .A2(n759), .ZN(n736) );
  NOR2_X1 U829 ( .A1(G2090), .A2(n691), .ZN(n735) );
  NOR2_X1 U830 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U831 ( .A1(n737), .A2(G303), .ZN(n738) );
  NAND2_X1 U832 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U833 ( .A(KEYINPUT101), .B(KEYINPUT32), .Z(n742) );
  NAND2_X1 U834 ( .A1(n754), .A2(n756), .ZN(n746) );
  NOR2_X1 U835 ( .A1(G2090), .A2(G303), .ZN(n744) );
  NAND2_X1 U836 ( .A1(G8), .A2(n744), .ZN(n745) );
  NAND2_X1 U837 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U838 ( .A1(n759), .A2(n747), .ZN(n748) );
  NAND2_X1 U839 ( .A1(n749), .A2(n748), .ZN(n771) );
  XNOR2_X1 U840 ( .A(G1981), .B(G305), .ZN(n970) );
  NAND2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n964) );
  INV_X1 U842 ( .A(KEYINPUT33), .ZN(n763) );
  NOR2_X1 U843 ( .A1(G288), .A2(G1976), .ZN(n750) );
  XNOR2_X1 U844 ( .A(n750), .B(KEYINPUT102), .ZN(n976) );
  NAND2_X1 U845 ( .A1(n751), .A2(n976), .ZN(n752) );
  NOR2_X1 U846 ( .A1(n763), .A2(n752), .ZN(n753) );
  XNOR2_X1 U847 ( .A(n753), .B(KEYINPUT103), .ZN(n762) );
  AND2_X1 U848 ( .A1(n964), .A2(n762), .ZN(n757) );
  AND2_X1 U849 ( .A1(n754), .A2(n757), .ZN(n755) );
  NAND2_X1 U850 ( .A1(n756), .A2(n755), .ZN(n768) );
  INV_X1 U851 ( .A(n757), .ZN(n761) );
  NOR2_X1 U852 ( .A1(G1971), .A2(G303), .ZN(n987) );
  NOR2_X1 U853 ( .A1(n976), .A2(n987), .ZN(n758) );
  OR2_X1 U854 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U855 ( .A1(n761), .A2(n760), .ZN(n766) );
  INV_X1 U856 ( .A(n762), .ZN(n764) );
  NOR2_X1 U857 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U858 ( .A1(n766), .A2(n765), .ZN(n767) );
  AND2_X1 U859 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U860 ( .A1(n970), .A2(n769), .ZN(n770) );
  NOR2_X1 U861 ( .A1(n773), .A2(n772), .ZN(n817) );
  NAND2_X1 U862 ( .A1(n878), .A2(G119), .ZN(n775) );
  NAND2_X1 U863 ( .A1(G131), .A2(n883), .ZN(n774) );
  NAND2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n779) );
  NAND2_X1 U865 ( .A1(G95), .A2(n882), .ZN(n777) );
  NAND2_X1 U866 ( .A1(G107), .A2(n879), .ZN(n776) );
  NAND2_X1 U867 ( .A1(n777), .A2(n776), .ZN(n778) );
  OR2_X1 U868 ( .A1(n779), .A2(n778), .ZN(n870) );
  NAND2_X1 U869 ( .A1(G1991), .A2(n870), .ZN(n790) );
  NAND2_X1 U870 ( .A1(n878), .A2(G129), .ZN(n780) );
  XOR2_X1 U871 ( .A(KEYINPUT91), .B(n780), .Z(n782) );
  NAND2_X1 U872 ( .A1(n879), .A2(G117), .ZN(n781) );
  NAND2_X1 U873 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U874 ( .A(KEYINPUT92), .B(n783), .ZN(n786) );
  NAND2_X1 U875 ( .A1(n882), .A2(G105), .ZN(n784) );
  XOR2_X1 U876 ( .A(KEYINPUT38), .B(n784), .Z(n785) );
  NOR2_X1 U877 ( .A1(n786), .A2(n785), .ZN(n788) );
  NAND2_X1 U878 ( .A1(G141), .A2(n883), .ZN(n787) );
  NAND2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n865) );
  NAND2_X1 U880 ( .A1(G1996), .A2(n865), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n927) );
  NAND2_X1 U882 ( .A1(n817), .A2(n927), .ZN(n791) );
  XNOR2_X1 U883 ( .A(KEYINPUT93), .B(n791), .ZN(n809) );
  NAND2_X1 U884 ( .A1(G128), .A2(n878), .ZN(n793) );
  NAND2_X1 U885 ( .A1(G116), .A2(n879), .ZN(n792) );
  NAND2_X1 U886 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U887 ( .A(KEYINPUT35), .B(n794), .ZN(n800) );
  NAND2_X1 U888 ( .A1(n882), .A2(G104), .ZN(n796) );
  NAND2_X1 U889 ( .A1(G140), .A2(n883), .ZN(n795) );
  NAND2_X1 U890 ( .A1(n796), .A2(n795), .ZN(n798) );
  XOR2_X1 U891 ( .A(KEYINPUT88), .B(KEYINPUT34), .Z(n797) );
  XNOR2_X1 U892 ( .A(n798), .B(n797), .ZN(n799) );
  NAND2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n801) );
  XOR2_X1 U894 ( .A(KEYINPUT36), .B(n801), .Z(n866) );
  XNOR2_X1 U895 ( .A(KEYINPUT37), .B(G2067), .ZN(n815) );
  OR2_X1 U896 ( .A1(n866), .A2(n815), .ZN(n802) );
  XNOR2_X1 U897 ( .A(n802), .B(KEYINPUT89), .ZN(n931) );
  NAND2_X1 U898 ( .A1(n817), .A2(n931), .ZN(n803) );
  XNOR2_X1 U899 ( .A(KEYINPUT90), .B(n803), .ZN(n812) );
  INV_X1 U900 ( .A(n812), .ZN(n804) );
  NOR2_X1 U901 ( .A1(n809), .A2(n804), .ZN(n805) );
  XOR2_X1 U902 ( .A(KEYINPUT94), .B(n805), .Z(n806) );
  XNOR2_X1 U903 ( .A(G1986), .B(G290), .ZN(n978) );
  NAND2_X1 U904 ( .A1(n518), .A2(n516), .ZN(n820) );
  NOR2_X1 U905 ( .A1(G1996), .A2(n865), .ZN(n920) );
  NOR2_X1 U906 ( .A1(G1991), .A2(n870), .ZN(n923) );
  NOR2_X1 U907 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U908 ( .A1(n923), .A2(n807), .ZN(n808) );
  NOR2_X1 U909 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U910 ( .A1(n920), .A2(n810), .ZN(n811) );
  XNOR2_X1 U911 ( .A(KEYINPUT39), .B(n811), .ZN(n813) );
  NAND2_X1 U912 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U913 ( .A(n814), .B(KEYINPUT104), .ZN(n816) );
  NAND2_X1 U914 ( .A1(n815), .A2(n866), .ZN(n933) );
  NAND2_X1 U915 ( .A1(n816), .A2(n933), .ZN(n818) );
  NAND2_X1 U916 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U917 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U918 ( .A(n821), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n822), .ZN(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U921 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U923 ( .A1(n825), .A2(n824), .ZN(G188) );
  NOR2_X1 U925 ( .A1(n827), .A2(n826), .ZN(n828) );
  XOR2_X1 U926 ( .A(KEYINPUT105), .B(n828), .Z(G325) );
  XOR2_X1 U927 ( .A(KEYINPUT106), .B(G325), .Z(G261) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  XOR2_X1 U929 ( .A(KEYINPUT107), .B(G2084), .Z(n830) );
  XNOR2_X1 U930 ( .A(G2078), .B(G2072), .ZN(n829) );
  XNOR2_X1 U931 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U932 ( .A(n831), .B(G2100), .Z(n833) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2090), .ZN(n832) );
  XNOR2_X1 U934 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U935 ( .A(G2096), .B(KEYINPUT43), .Z(n835) );
  XNOR2_X1 U936 ( .A(KEYINPUT42), .B(G2678), .ZN(n834) );
  XNOR2_X1 U937 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U938 ( .A(n837), .B(n836), .Z(G227) );
  XNOR2_X1 U939 ( .A(G1956), .B(KEYINPUT108), .ZN(n847) );
  XOR2_X1 U940 ( .A(G1976), .B(G1981), .Z(n839) );
  XNOR2_X1 U941 ( .A(G1966), .B(G1961), .ZN(n838) );
  XNOR2_X1 U942 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U943 ( .A(G1971), .B(G1986), .Z(n841) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1991), .ZN(n840) );
  XNOR2_X1 U945 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U946 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U947 ( .A(G2474), .B(KEYINPUT41), .ZN(n844) );
  XNOR2_X1 U948 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(G229) );
  NAND2_X1 U950 ( .A1(n878), .A2(G124), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n848), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U952 ( .A1(G136), .A2(n883), .ZN(n849) );
  NAND2_X1 U953 ( .A1(n850), .A2(n849), .ZN(n851) );
  XOR2_X1 U954 ( .A(KEYINPUT109), .B(n851), .Z(n857) );
  NAND2_X1 U955 ( .A1(n879), .A2(G112), .ZN(n852) );
  XNOR2_X1 U956 ( .A(n852), .B(KEYINPUT110), .ZN(n854) );
  NAND2_X1 U957 ( .A1(G100), .A2(n882), .ZN(n853) );
  NAND2_X1 U958 ( .A1(n854), .A2(n853), .ZN(n855) );
  XOR2_X1 U959 ( .A(KEYINPUT111), .B(n855), .Z(n856) );
  NOR2_X1 U960 ( .A1(n857), .A2(n856), .ZN(G162) );
  NAND2_X1 U961 ( .A1(n882), .A2(G103), .ZN(n859) );
  NAND2_X1 U962 ( .A1(G139), .A2(n883), .ZN(n858) );
  NAND2_X1 U963 ( .A1(n859), .A2(n858), .ZN(n864) );
  NAND2_X1 U964 ( .A1(G127), .A2(n878), .ZN(n861) );
  NAND2_X1 U965 ( .A1(G115), .A2(n879), .ZN(n860) );
  NAND2_X1 U966 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U967 ( .A(KEYINPUT47), .B(n862), .Z(n863) );
  NOR2_X1 U968 ( .A1(n864), .A2(n863), .ZN(n914) );
  XNOR2_X1 U969 ( .A(n865), .B(n914), .ZN(n868) );
  XOR2_X1 U970 ( .A(G160), .B(n866), .Z(n867) );
  XNOR2_X1 U971 ( .A(n868), .B(n867), .ZN(n872) );
  XOR2_X1 U972 ( .A(G164), .B(n922), .Z(n869) );
  XNOR2_X1 U973 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U974 ( .A(n872), .B(n871), .Z(n877) );
  XOR2_X1 U975 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n874) );
  XNOR2_X1 U976 ( .A(KEYINPUT48), .B(KEYINPUT114), .ZN(n873) );
  XNOR2_X1 U977 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U978 ( .A(KEYINPUT46), .B(n875), .ZN(n876) );
  XNOR2_X1 U979 ( .A(n877), .B(n876), .ZN(n891) );
  NAND2_X1 U980 ( .A1(G130), .A2(n878), .ZN(n881) );
  NAND2_X1 U981 ( .A1(G118), .A2(n879), .ZN(n880) );
  NAND2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n888) );
  NAND2_X1 U983 ( .A1(n882), .A2(G106), .ZN(n885) );
  NAND2_X1 U984 ( .A1(G142), .A2(n883), .ZN(n884) );
  NAND2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U986 ( .A(KEYINPUT45), .B(n886), .Z(n887) );
  NOR2_X1 U987 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U988 ( .A(G162), .B(n889), .Z(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U990 ( .A1(G37), .A2(n892), .ZN(G395) );
  XNOR2_X1 U991 ( .A(n893), .B(G286), .ZN(n895) );
  XNOR2_X1 U992 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n896), .B(G171), .ZN(n897) );
  NOR2_X1 U994 ( .A1(G37), .A2(n897), .ZN(G397) );
  XOR2_X1 U995 ( .A(G2451), .B(G2430), .Z(n899) );
  XNOR2_X1 U996 ( .A(G2438), .B(G2443), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n905) );
  XOR2_X1 U998 ( .A(G2435), .B(G2454), .Z(n901) );
  XNOR2_X1 U999 ( .A(G1341), .B(G1348), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n901), .B(n900), .ZN(n903) );
  XOR2_X1 U1001 ( .A(G2446), .B(G2427), .Z(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1003 ( .A(n905), .B(n904), .Z(n906) );
  NAND2_X1 U1004 ( .A1(G14), .A2(n906), .ZN(n913) );
  NAND2_X1 U1005 ( .A1(n913), .A2(G319), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n907) );
  XOR2_X1 U1007 ( .A(KEYINPUT115), .B(n907), .Z(n908) );
  XNOR2_X1 U1008 ( .A(n908), .B(KEYINPUT49), .ZN(n909) );
  NOR2_X1 U1009 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1011 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(n913), .ZN(G401) );
  XNOR2_X1 U1014 ( .A(G2072), .B(n914), .ZN(n917) );
  XOR2_X1 U1015 ( .A(G164), .B(G2078), .Z(n915) );
  XNOR2_X1 U1016 ( .A(KEYINPUT117), .B(n915), .ZN(n916) );
  NAND2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(n918), .B(KEYINPUT50), .ZN(n936) );
  XOR2_X1 U1019 ( .A(G2090), .B(G162), .Z(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1021 ( .A(KEYINPUT51), .B(n921), .Z(n929) );
  XNOR2_X1 U1022 ( .A(G160), .B(G2084), .ZN(n925) );
  NOR2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(n932), .B(KEYINPUT116), .ZN(n934) );
  NAND2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1031 ( .A(KEYINPUT52), .B(n937), .ZN(n939) );
  INV_X1 U1032 ( .A(KEYINPUT55), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1034 ( .A1(n940), .A2(G29), .ZN(n1022) );
  XNOR2_X1 U1035 ( .A(G2084), .B(G34), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(n941), .B(KEYINPUT54), .ZN(n958) );
  XOR2_X1 U1037 ( .A(G27), .B(n942), .Z(n951) );
  XNOR2_X1 U1038 ( .A(G1996), .B(G32), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(G33), .B(G2072), .ZN(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n949) );
  XOR2_X1 U1041 ( .A(G1991), .B(G25), .Z(n945) );
  NAND2_X1 U1042 ( .A1(n945), .A2(G28), .ZN(n947) );
  XNOR2_X1 U1043 ( .A(G26), .B(G2067), .ZN(n946) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n950) );
  NOR2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(KEYINPUT53), .B(KEYINPUT118), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(n953), .B(n952), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(G35), .B(G2090), .ZN(n954) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(n956), .B(KEYINPUT119), .ZN(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1053 ( .A(KEYINPUT55), .B(n959), .Z(n960) );
  NOR2_X1 U1054 ( .A1(G29), .A2(n960), .ZN(n961) );
  XOR2_X1 U1055 ( .A(KEYINPUT120), .B(n961), .Z(n962) );
  NAND2_X1 U1056 ( .A1(G11), .A2(n962), .ZN(n1020) );
  XOR2_X1 U1057 ( .A(G16), .B(KEYINPUT56), .Z(n989) );
  NAND2_X1 U1058 ( .A1(G1971), .A2(G303), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(G1348), .B(n965), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n974) );
  XNOR2_X1 U1062 ( .A(KEYINPUT122), .B(KEYINPUT57), .ZN(n972) );
  XNOR2_X1 U1063 ( .A(G1966), .B(G168), .ZN(n968) );
  XNOR2_X1 U1064 ( .A(n968), .B(KEYINPUT121), .ZN(n969) );
  NOR2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1066 ( .A(n972), .B(n971), .Z(n973) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n985) );
  XNOR2_X1 U1069 ( .A(G171), .B(G1961), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(G1956), .B(G299), .ZN(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n983) );
  XNOR2_X1 U1073 ( .A(G1341), .B(n981), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n1017) );
  XNOR2_X1 U1078 ( .A(n990), .B(G20), .ZN(n999) );
  XOR2_X1 U1079 ( .A(KEYINPUT124), .B(G4), .Z(n992) );
  XNOR2_X1 U1080 ( .A(G1348), .B(KEYINPUT59), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(n992), .B(n991), .ZN(n997) );
  XNOR2_X1 U1082 ( .A(G1341), .B(G19), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(G1981), .B(G6), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(n995), .B(KEYINPUT123), .ZN(n996) );
  NOR2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(n1000), .B(KEYINPUT60), .ZN(n1008) );
  XNOR2_X1 U1089 ( .A(G1971), .B(G22), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(G23), .B(G1976), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(G1986), .B(KEYINPUT125), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(n1003), .B(G24), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(KEYINPUT58), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(G1966), .B(G21), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(G1961), .B(G5), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(n1013), .B(KEYINPUT61), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(n1014), .B(KEYINPUT126), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(G16), .A2(n1015), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(KEYINPUT127), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1023), .Z(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

