//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G137), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G131), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n191), .A2(new_n193), .A3(new_n197), .A4(new_n194), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT1), .B1(new_n201), .B2(G146), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(G146), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  OAI211_X1 g019(.A(G128), .B(new_n202), .C1(new_n203), .C2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G107), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(G101), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT3), .B1(new_n207), .B2(G107), .ZN(new_n212));
  AOI21_X1  g026(.A(G101), .B1(new_n207), .B2(G107), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT3), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(new_n209), .A3(G104), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n212), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n204), .A2(G143), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n201), .A2(G146), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n217), .B(new_n218), .C1(KEYINPUT1), .C2(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n206), .A2(new_n211), .A3(new_n216), .A4(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT10), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n221), .B(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n207), .A2(G107), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n212), .A2(new_n215), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT79), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n212), .A2(new_n215), .A3(KEYINPUT79), .A4(new_n225), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT80), .B1(new_n230), .B2(G101), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT80), .ZN(new_n232));
  INV_X1    g046(.A(G101), .ZN(new_n233));
  AOI211_X1 g047(.A(new_n232), .B(new_n233), .C1(new_n228), .C2(new_n229), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n216), .A2(KEYINPUT4), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n231), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT0), .A4(G128), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n203), .A2(new_n205), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT0), .B(G128), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT81), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G101), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n242), .B1(new_n230), .B2(new_n245), .ZN(new_n246));
  AOI211_X1 g060(.A(KEYINPUT81), .B(new_n244), .C1(new_n228), .C2(new_n229), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n241), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n200), .B(new_n224), .C1(new_n236), .C2(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(G110), .B(G140), .ZN(new_n250));
  INV_X1    g064(.A(G953), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n251), .A2(G227), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n250), .B(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT83), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n206), .A2(new_n220), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n211), .A2(new_n216), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n220), .A2(new_n206), .B1(new_n211), .B2(new_n216), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n257), .A2(new_n258), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(KEYINPUT83), .A3(new_n221), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(new_n199), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT12), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT84), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT84), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n264), .A2(new_n268), .A3(new_n265), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(KEYINPUT82), .A2(KEYINPUT12), .ZN(new_n271));
  AND2_X1   g085(.A1(KEYINPUT82), .A2(KEYINPUT12), .ZN(new_n272));
  OAI221_X1 g086(.A(new_n199), .B1(new_n271), .B2(new_n272), .C1(new_n259), .C2(new_n260), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n255), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n224), .B1(new_n236), .B2(new_n248), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n199), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n254), .B1(new_n276), .B2(new_n249), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n187), .B(new_n188), .C1(new_n274), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT85), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n264), .A2(new_n268), .A3(new_n265), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n268), .B1(new_n264), .B2(new_n265), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n273), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n230), .A2(new_n245), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT81), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n230), .A2(new_n242), .A3(new_n245), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n240), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n231), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n233), .B1(new_n228), .B2(new_n229), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n235), .B1(new_n288), .B2(KEYINPUT80), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n223), .B1(new_n286), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n253), .B1(new_n291), .B2(new_n200), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n282), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n286), .A2(new_n290), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n200), .B1(new_n294), .B2(new_n224), .ZN(new_n295));
  AOI211_X1 g109(.A(new_n199), .B(new_n223), .C1(new_n286), .C2(new_n290), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n253), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT85), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n298), .A2(new_n299), .A3(new_n187), .A4(new_n188), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n254), .B1(new_n282), .B2(new_n249), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n255), .A2(new_n295), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n188), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n279), .A2(new_n300), .B1(G469), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(G113), .B(G122), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n305), .B(new_n207), .ZN(new_n306));
  INV_X1    g120(.A(G237), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(new_n251), .A3(G214), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n201), .ZN(new_n309));
  NOR2_X1   g123(.A1(G237), .A2(G953), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(G143), .A3(G214), .ZN(new_n311));
  NAND2_X1  g125(.A1(KEYINPUT18), .A2(G131), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(KEYINPUT89), .ZN(new_n314));
  INV_X1    g128(.A(G140), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G125), .ZN(new_n316));
  INV_X1    g130(.A(G125), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G140), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n316), .A2(new_n318), .A3(KEYINPUT77), .ZN(new_n319));
  OR3_X1    g133(.A1(new_n317), .A2(KEYINPUT77), .A3(G140), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(G146), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n316), .A2(new_n318), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n204), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n309), .A2(new_n311), .ZN(new_n324));
  INV_X1    g138(.A(new_n312), .ZN(new_n325));
  AOI22_X1  g139(.A1(new_n321), .A2(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n314), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n309), .A2(new_n197), .A3(new_n311), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT90), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n324), .A2(G131), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT90), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n309), .A2(new_n331), .A3(new_n197), .A4(new_n311), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  OR2_X1    g147(.A1(new_n333), .A2(KEYINPUT17), .ZN(new_n334));
  AND4_X1   g148(.A1(G143), .A2(new_n307), .A3(new_n251), .A4(G214), .ZN(new_n335));
  AOI21_X1  g149(.A(G143), .B1(new_n310), .B2(G214), .ZN(new_n336));
  OAI211_X1 g150(.A(KEYINPUT17), .B(G131), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT92), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT92), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n324), .A2(new_n339), .A3(KEYINPUT17), .A4(G131), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n319), .A2(new_n320), .A3(KEYINPUT16), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT16), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n316), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n204), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n344), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G146), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n341), .A2(KEYINPUT93), .A3(new_n345), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n334), .A2(new_n348), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n342), .A2(new_n204), .A3(new_n344), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n204), .B1(new_n342), .B2(new_n344), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT93), .B1(new_n352), .B2(new_n341), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n306), .B(new_n327), .C1(new_n349), .C2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n341), .A2(new_n345), .A3(new_n347), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT93), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(new_n334), .A3(new_n348), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n306), .B1(new_n359), .B2(new_n327), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n188), .B1(new_n355), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G475), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT19), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(new_n319), .B2(new_n320), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n322), .A2(KEYINPUT19), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n333), .B(new_n347), .C1(G146), .C2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n306), .B1(new_n367), .B2(new_n327), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT91), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI211_X1 g184(.A(KEYINPUT91), .B(new_n306), .C1(new_n367), .C2(new_n327), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n354), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT20), .ZN(new_n373));
  NOR2_X1   g187(.A1(G475), .A2(G902), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n373), .B1(new_n372), .B2(new_n374), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n362), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT73), .B(G217), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT9), .B(G234), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n378), .A2(new_n379), .A3(G953), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n201), .A2(G128), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n219), .A2(G143), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n383), .B(new_n190), .ZN(new_n384));
  XNOR2_X1  g198(.A(G116), .B(G122), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n209), .ZN(new_n386));
  INV_X1    g200(.A(G116), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(KEYINPUT14), .A3(G122), .ZN(new_n388));
  INV_X1    g202(.A(new_n385), .ZN(new_n389));
  OAI211_X1 g203(.A(G107), .B(new_n388), .C1(new_n389), .C2(KEYINPUT14), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n384), .A2(new_n386), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n381), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n392), .A2(KEYINPUT13), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n382), .B1(new_n392), .B2(KEYINPUT13), .ZN(new_n394));
  OAI21_X1  g208(.A(G134), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n383), .A2(new_n190), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n385), .B(new_n209), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n380), .B1(new_n391), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n391), .A2(new_n398), .A3(new_n380), .ZN(new_n401));
  AOI21_X1  g215(.A(G902), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT15), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G478), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n402), .A2(new_n404), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n251), .A2(G952), .ZN(new_n409));
  INV_X1    g223(.A(G234), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n409), .B1(new_n410), .B2(new_n307), .ZN(new_n411));
  INV_X1    g225(.A(G898), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n251), .B1(KEYINPUT21), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n413), .B1(KEYINPUT21), .B2(new_n412), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n188), .B1(G234), .B2(G237), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n411), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  XOR2_X1   g231(.A(new_n417), .B(KEYINPUT94), .Z(new_n418));
  NAND2_X1  g232(.A1(new_n408), .A2(new_n418), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n377), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G221), .ZN(new_n421));
  INV_X1    g235(.A(new_n379), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n421), .B1(new_n422), .B2(new_n188), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n304), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n378), .B1(G234), .B2(new_n188), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G119), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G128), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n219), .A2(G119), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G110), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT24), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT24), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G110), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n432), .A2(new_n434), .A3(KEYINPUT74), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT74), .B1(new_n432), .B2(new_n434), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n430), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT23), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n438), .B1(new_n427), .B2(G128), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n219), .A2(KEYINPUT23), .A3(G119), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n428), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT78), .B(G110), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n437), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(new_n347), .A3(new_n323), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n431), .B1(new_n441), .B2(KEYINPUT75), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT76), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT75), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n439), .A2(new_n440), .A3(new_n447), .A4(new_n428), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n445), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n446), .B1(new_n445), .B2(new_n448), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OR3_X1    g265(.A1(new_n435), .A2(new_n436), .A3(new_n430), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(new_n350), .B2(new_n351), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n444), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT22), .B(G137), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n421), .A2(new_n410), .A3(G953), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n455), .B(new_n456), .Z(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n444), .B(new_n457), .C1(new_n451), .C2(new_n453), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n188), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT25), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n459), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n460), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n426), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n459), .A2(new_n460), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n425), .A2(G902), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT31), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n206), .A2(new_n198), .A3(new_n220), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT64), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n474), .B1(new_n190), .B2(G137), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n192), .A2(KEYINPUT64), .A3(G134), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n194), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT65), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n478), .A3(G131), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(G131), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT65), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n473), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n241), .A2(new_n199), .ZN(new_n483));
  XNOR2_X1  g297(.A(G116), .B(G119), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT2), .B(G113), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n484), .B(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n482), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n479), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n206), .A2(new_n198), .A3(new_n220), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n478), .B1(new_n477), .B2(G131), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n240), .B1(new_n196), .B2(new_n198), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT30), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT30), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n482), .A2(new_n483), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n486), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n488), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT68), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT26), .B(G101), .Z(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n500), .B(KEYINPUT68), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n503), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n310), .A2(G210), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT67), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n508), .B(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n472), .B1(new_n499), .B2(new_n511), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n482), .A2(new_n483), .A3(new_n495), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n495), .B1(new_n482), .B2(new_n483), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n498), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AND4_X1   g329(.A1(new_n472), .A2(new_n515), .A3(new_n487), .A4(new_n511), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT70), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n482), .A2(new_n483), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT69), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT69), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n482), .A2(new_n483), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(new_n486), .A3(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT28), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n498), .B1(new_n492), .B2(new_n493), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n524), .B1(new_n526), .B2(new_n487), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  XOR2_X1   g343(.A(new_n508), .B(new_n510), .Z(new_n530));
  AOI21_X1  g344(.A(new_n518), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI211_X1 g345(.A(KEYINPUT70), .B(new_n511), .C1(new_n525), .C2(new_n528), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n517), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(G472), .A2(G902), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT71), .B(KEYINPUT32), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n534), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT32), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT72), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n542), .B1(new_n526), .B2(new_n487), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n487), .A2(new_n542), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT28), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n511), .A2(KEYINPUT29), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n546), .A3(new_n525), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT29), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n499), .B2(new_n511), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n498), .B1(new_n519), .B2(KEYINPUT69), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT28), .B1(new_n550), .B2(new_n522), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n551), .A2(new_n530), .A3(new_n527), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n547), .B(new_n188), .C1(new_n549), .C2(new_n552), .ZN(new_n553));
  AOI22_X1  g367(.A1(new_n533), .A2(new_n541), .B1(G472), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n471), .B1(new_n538), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(G214), .B1(G237), .B2(G902), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n484), .ZN(new_n558));
  XOR2_X1   g372(.A(KEYINPUT86), .B(KEYINPUT5), .Z(new_n559));
  OR2_X1    g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(G113), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n387), .A2(G119), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n561), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n558), .A2(new_n485), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n258), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n498), .B1(new_n246), .B2(new_n247), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n567), .B1(new_n236), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(G110), .B(G122), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n570), .B(new_n567), .C1(new_n236), .C2(new_n568), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT6), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n257), .A2(new_n317), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n240), .A2(G125), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(G224), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(G953), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n575), .B(new_n576), .C1(new_n578), .C2(G953), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT6), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n569), .A2(new_n583), .A3(new_n571), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n574), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT87), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT87), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n574), .A2(new_n587), .A3(new_n582), .A4(new_n584), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT88), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT5), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n563), .B1(new_n591), .B2(new_n558), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n566), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n565), .B1(new_n560), .B2(new_n563), .ZN(new_n594));
  INV_X1    g408(.A(new_n258), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n570), .B(KEYINPUT8), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n579), .A2(KEYINPUT7), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n577), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n599), .B1(new_n580), .B2(new_n581), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n590), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n602), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n604), .A2(KEYINPUT88), .A3(new_n600), .A4(new_n598), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n603), .A2(new_n605), .A3(new_n573), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n188), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n589), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(G210), .B1(G237), .B2(G902), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n589), .A2(new_n610), .A3(new_n608), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n557), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n424), .A2(new_n555), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  NAND2_X1  g430(.A1(new_n279), .A2(new_n300), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n303), .A2(G469), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n423), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n515), .A2(new_n487), .A3(new_n511), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(KEYINPUT31), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n499), .A2(new_n472), .A3(new_n511), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n551), .A2(new_n527), .ZN(new_n624));
  OAI21_X1  g438(.A(KEYINPUT70), .B1(new_n624), .B2(new_n511), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n529), .A2(new_n518), .A3(new_n530), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(G472), .B1(new_n627), .B2(G902), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n535), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(new_n471), .ZN(new_n630));
  INV_X1    g444(.A(new_n401), .ZN(new_n631));
  OR2_X1    g445(.A1(new_n631), .A2(KEYINPUT96), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(KEYINPUT96), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n632), .A2(KEYINPUT33), .A3(new_n633), .A4(new_n400), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT95), .B(KEYINPUT33), .Z(new_n635));
  OAI21_X1  g449(.A(new_n635), .B1(new_n631), .B2(new_n399), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n188), .A2(G478), .ZN(new_n638));
  OAI22_X1  g452(.A1(new_n637), .A2(new_n638), .B1(G478), .B2(new_n402), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n377), .A2(new_n418), .A3(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n614), .A2(new_n619), .A3(new_n630), .A4(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  INV_X1    g457(.A(new_n300), .ZN(new_n644));
  AOI21_X1  g458(.A(G902), .B1(new_n293), .B2(new_n297), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n299), .B1(new_n645), .B2(new_n187), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n618), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n625), .A2(new_n626), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n539), .B1(new_n648), .B2(new_n517), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n533), .A2(new_n188), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n649), .B1(new_n650), .B2(G472), .ZN(new_n651));
  INV_X1    g465(.A(new_n423), .ZN(new_n652));
  AND4_X1   g466(.A1(new_n470), .A2(new_n647), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n418), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n377), .A2(new_n408), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n610), .B1(new_n589), .B2(new_n608), .ZN(new_n656));
  AOI211_X1 g470(.A(new_n611), .B(new_n607), .C1(new_n586), .C2(new_n588), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n655), .B(new_n556), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT35), .B(G107), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n463), .A2(new_n464), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n425), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n454), .A2(KEYINPUT97), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n458), .A2(KEYINPUT36), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT97), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n668), .B(new_n444), .C1(new_n451), .C2(new_n453), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n666), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n667), .B1(new_n666), .B2(new_n669), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n467), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n665), .A2(KEYINPUT98), .A3(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT98), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n666), .A2(new_n669), .ZN(new_n676));
  INV_X1    g490(.A(new_n667), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n468), .B1(new_n678), .B2(new_n670), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n675), .B1(new_n465), .B2(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n663), .B1(new_n629), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n674), .A2(new_n680), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n651), .A2(KEYINPUT99), .A3(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n424), .A2(new_n614), .A3(new_n682), .A4(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT37), .B(G110), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT100), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n685), .B(new_n687), .ZN(G12));
  NAND2_X1  g502(.A1(new_n647), .A2(new_n652), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n251), .A2(G900), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n415), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n691), .A2(KEYINPUT101), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(KEYINPUT101), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n692), .A2(new_n411), .A3(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n407), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n695), .B1(new_n696), .B2(new_n405), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n362), .B(new_n697), .C1(new_n375), .C2(new_n376), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n553), .A2(G472), .ZN(new_n700));
  INV_X1    g514(.A(new_n541), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n700), .B1(new_n627), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n536), .B1(new_n533), .B2(new_n534), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n699), .B(new_n683), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n689), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(KEYINPUT102), .A3(new_n614), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT102), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n538), .A2(new_n554), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n698), .B1(new_n680), .B2(new_n674), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n708), .A2(new_n709), .A3(new_n647), .A4(new_n652), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n556), .B1(new_n656), .B2(new_n657), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n707), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n706), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G128), .ZN(G30));
  XNOR2_X1  g528(.A(new_n694), .B(KEYINPUT39), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n619), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT40), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n612), .A2(new_n613), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n499), .A2(new_n530), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n543), .A2(new_n544), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n722), .B(new_n188), .C1(new_n511), .C2(new_n723), .ZN(new_n724));
  AOI22_X1  g538(.A1(new_n533), .A2(new_n541), .B1(new_n724), .B2(G472), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n538), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n376), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n728));
  AOI22_X1  g542(.A1(new_n727), .A2(new_n728), .B1(G475), .B2(new_n361), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n408), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n726), .A2(new_n556), .A3(new_n681), .A4(new_n730), .ZN(new_n731));
  OR3_X1    g545(.A1(new_n717), .A2(new_n720), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G143), .ZN(G45));
  INV_X1    g547(.A(KEYINPUT104), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n377), .A2(new_n639), .A3(new_n694), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n734), .B1(new_n711), .B2(new_n735), .ZN(new_n736));
  AND4_X1   g550(.A1(new_n708), .A2(new_n652), .A3(new_n647), .A4(new_n683), .ZN(new_n737));
  INV_X1    g551(.A(new_n735), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n718), .A2(KEYINPUT104), .A3(new_n556), .A4(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n736), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G146), .ZN(G48));
  OR2_X1    g555(.A1(new_n645), .A2(new_n187), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n617), .A2(new_n652), .A3(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n614), .A2(new_n555), .A3(new_n640), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  NAND4_X1  g560(.A1(new_n614), .A2(new_n555), .A3(new_n655), .A4(new_n743), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G116), .ZN(G18));
  NOR2_X1   g562(.A1(new_n377), .A2(new_n419), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n749), .B(new_n683), .C1(new_n702), .C2(new_n703), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n614), .A3(new_n743), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G119), .ZN(G21));
  AOI21_X1  g567(.A(new_n511), .B1(new_n545), .B2(new_n525), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n534), .B1(new_n623), .B2(new_n754), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n628), .A2(new_n470), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n743), .A2(new_n418), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT105), .B1(new_n614), .B2(new_n730), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n730), .B(new_n556), .C1(new_n656), .C2(new_n657), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT105), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n758), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G122), .ZN(G24));
  NAND3_X1  g578(.A1(new_n617), .A2(new_n652), .A3(new_n742), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n711), .A2(new_n765), .ZN(new_n766));
  AND4_X1   g580(.A1(new_n628), .A2(new_n738), .A3(new_n683), .A4(new_n755), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G125), .ZN(G27));
  INV_X1    g583(.A(KEYINPUT42), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n656), .A2(new_n657), .A3(new_n557), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT106), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n772), .B1(new_n304), .B2(new_n423), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n647), .A2(KEYINPUT106), .A3(new_n652), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n771), .A2(new_n773), .A3(new_n774), .A4(new_n555), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n770), .B1(new_n775), .B2(new_n735), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n735), .A2(new_n770), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n649), .A2(KEYINPUT32), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n778), .B(new_n470), .C1(new_n702), .C2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT107), .B1(new_n777), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT107), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n783), .A2(new_n784), .A3(new_n780), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n776), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G131), .ZN(G33));
  NOR2_X1   g601(.A1(new_n775), .A2(new_n698), .ZN(new_n788));
  XNOR2_X1  g602(.A(KEYINPUT108), .B(G134), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n788), .B(new_n789), .ZN(G36));
  INV_X1    g604(.A(KEYINPUT109), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT43), .B1(new_n729), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n729), .A2(new_n639), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n651), .A2(new_n681), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(KEYINPUT44), .A3(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n796), .A2(new_n771), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n794), .A2(new_n795), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n797), .B1(KEYINPUT44), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n301), .A2(new_n302), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n800), .A2(KEYINPUT45), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(KEYINPUT45), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(G469), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(G469), .A2(G902), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT46), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n805), .B1(new_n300), .B2(new_n279), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n803), .A2(KEYINPUT46), .A3(new_n804), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n652), .A3(new_n715), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n799), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(new_n192), .ZN(G39));
  AOI21_X1  g625(.A(new_n423), .B1(new_n806), .B2(new_n807), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT47), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n708), .A2(new_n470), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n738), .A3(new_n771), .ZN(new_n815));
  XOR2_X1   g629(.A(new_n815), .B(KEYINPUT110), .Z(new_n816));
  NAND2_X1  g630(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G140), .ZN(G42));
  INV_X1    g632(.A(new_n411), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n794), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n820), .A2(new_n756), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n557), .A3(new_n720), .A4(new_n743), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT50), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n718), .A2(new_n765), .A3(new_n557), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  AND4_X1   g639(.A1(new_n628), .A2(new_n825), .A3(new_n683), .A4(new_n755), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n726), .A2(new_n471), .A3(new_n411), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n828), .A2(new_n377), .A3(new_n639), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n823), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n617), .A2(new_n742), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n652), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n771), .B(new_n821), .C1(new_n813), .C2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT51), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n470), .B1(new_n779), .B2(new_n702), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n825), .A2(new_n836), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n837), .B(KEYINPUT48), .Z(new_n838));
  NAND2_X1  g652(.A1(new_n377), .A2(new_n639), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n828), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n821), .A2(new_n766), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n409), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n834), .A2(new_n838), .A3(new_n840), .A4(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT111), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n615), .A2(new_n641), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n845), .B1(new_n615), .B2(new_n641), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT99), .B1(new_n651), .B2(new_n683), .ZN(new_n849));
  AND4_X1   g663(.A1(KEYINPUT99), .A2(new_n683), .A3(new_n628), .A4(new_n535), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n647), .A2(new_n652), .A3(new_n749), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n711), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n640), .B(new_n556), .C1(new_n656), .C2(new_n657), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n470), .B1(new_n702), .B2(new_n703), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n765), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n851), .A2(new_n853), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n718), .A2(KEYINPUT112), .A3(new_n556), .A4(new_n655), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT112), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n658), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n861), .A3(new_n653), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n766), .A2(new_n751), .B1(new_n659), .B2(new_n857), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n763), .A2(new_n858), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n848), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n767), .A2(new_n771), .A3(new_n773), .A4(new_n774), .ZN(new_n866));
  INV_X1    g680(.A(new_n408), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n377), .A2(new_n867), .A3(new_n695), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT113), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n737), .A2(new_n869), .A3(new_n771), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n866), .B(new_n870), .C1(new_n698), .C2(new_n775), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n777), .A2(KEYINPUT107), .A3(new_n781), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n784), .B1(new_n783), .B2(new_n780), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n871), .B1(new_n874), .B2(new_n776), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n465), .A2(new_n679), .A3(new_n695), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT114), .B1(new_n619), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT114), .ZN(new_n878));
  INV_X1    g692(.A(new_n876), .ZN(new_n879));
  NOR4_X1   g693(.A1(new_n304), .A2(new_n878), .A3(new_n423), .A4(new_n879), .ZN(new_n880));
  OAI221_X1 g694(.A(new_n726), .B1(new_n877), .B2(new_n880), .C1(new_n759), .C2(new_n762), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n706), .A2(new_n712), .B1(new_n766), .B2(new_n767), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT52), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .A4(new_n740), .ZN(new_n884));
  XOR2_X1   g698(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n885));
  AOI21_X1  g699(.A(KEYINPUT102), .B1(new_n705), .B2(new_n614), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n710), .A2(new_n707), .A3(new_n711), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n740), .B(new_n768), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n760), .B(KEYINPUT105), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n726), .B1(new_n877), .B2(new_n880), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n885), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n865), .A2(new_n875), .A3(new_n884), .A4(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT52), .B1(new_n888), .B2(new_n891), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n884), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n685), .A2(new_n744), .A3(new_n747), .A4(new_n752), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n859), .A2(new_n861), .A3(new_n653), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n614), .A2(KEYINPUT105), .A3(new_n730), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n760), .A2(new_n761), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n757), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n900), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n615), .A2(new_n641), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT111), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n615), .A2(new_n641), .A3(new_n845), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n866), .A2(new_n870), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(new_n788), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n905), .A2(new_n786), .A3(new_n909), .A4(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n894), .B1(new_n899), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n896), .A2(new_n897), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT116), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n892), .A2(new_n884), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n915), .B(new_n894), .C1(new_n916), .C2(new_n912), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n915), .B1(new_n893), .B2(new_n894), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n899), .A2(new_n912), .A3(new_n894), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n844), .B(new_n914), .C1(new_n921), .C2(new_n897), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n894), .B1(new_n916), .B2(new_n912), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n899), .A2(new_n912), .ZN(new_n924));
  AOI22_X1  g738(.A1(new_n923), .A2(KEYINPUT116), .B1(new_n924), .B2(KEYINPUT53), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n897), .B1(new_n925), .B2(new_n917), .ZN(new_n926));
  INV_X1    g740(.A(new_n913), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n927), .A2(new_n895), .A3(KEYINPUT54), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT117), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n830), .A2(KEYINPUT51), .A3(new_n833), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n843), .A2(new_n922), .A3(new_n929), .A4(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(G952), .B2(G953), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n831), .A2(KEYINPUT49), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n470), .A2(new_n556), .A3(new_n652), .ZN(new_n934));
  NOR4_X1   g748(.A1(new_n933), .A2(new_n726), .A3(new_n793), .A4(new_n934), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n935), .B(new_n720), .C1(KEYINPUT49), .C2(new_n831), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n932), .A2(new_n936), .ZN(G75));
  NAND2_X1  g751(.A1(new_n896), .A2(new_n913), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n939), .A2(new_n188), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT56), .B1(new_n940), .B2(G210), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n574), .A2(new_n584), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(new_n582), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT55), .ZN(new_n944));
  OAI22_X1  g758(.A1(new_n941), .A2(new_n944), .B1(G952), .B2(new_n251), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n941), .B2(new_n944), .ZN(G51));
  NOR2_X1   g760(.A1(new_n251), .A2(G952), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n938), .A2(KEYINPUT54), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n914), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n804), .B(KEYINPUT57), .Z(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n298), .ZN(new_n952));
  OR3_X1    g766(.A1(new_n939), .A2(new_n188), .A3(new_n803), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n947), .B1(new_n952), .B2(new_n953), .ZN(G54));
  NAND3_X1  g768(.A1(new_n940), .A2(KEYINPUT58), .A3(G475), .ZN(new_n955));
  INV_X1    g769(.A(new_n372), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n957), .A2(new_n958), .A3(new_n947), .ZN(G60));
  XNOR2_X1  g773(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n960));
  NAND2_X1  g774(.A1(G478), .A2(G902), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n637), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n947), .B1(new_n949), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n962), .B1(new_n929), .B2(new_n922), .ZN(new_n965));
  INV_X1    g779(.A(new_n637), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(KEYINPUT119), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT119), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n969), .B(new_n964), .C1(new_n965), .C2(new_n966), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n968), .A2(new_n970), .ZN(G63));
  XOR2_X1   g785(.A(KEYINPUT120), .B(KEYINPUT60), .Z(new_n972));
  NAND2_X1  g786(.A1(G217), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n938), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n947), .B1(new_n975), .B2(new_n466), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n671), .A2(new_n672), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n976), .B1(new_n977), .B2(new_n975), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g793(.A(new_n414), .B1(G224), .B2(new_n251), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT121), .Z(new_n981));
  INV_X1    g795(.A(new_n865), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n981), .B1(new_n982), .B2(new_n251), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n942), .B1(G898), .B2(new_n251), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n983), .B(new_n984), .Z(G69));
  XOR2_X1   g799(.A(new_n497), .B(new_n366), .Z(new_n986));
  OR2_X1    g800(.A1(new_n810), .A2(new_n788), .ZN(new_n987));
  INV_X1    g801(.A(new_n888), .ZN(new_n988));
  OR3_X1    g802(.A1(new_n809), .A2(new_n889), .A3(new_n835), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n817), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n786), .ZN(new_n991));
  OR4_X1    g805(.A1(KEYINPUT125), .A2(new_n987), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n987), .A2(new_n991), .ZN(new_n993));
  OAI21_X1  g807(.A(KEYINPUT125), .B1(new_n993), .B2(new_n990), .ZN(new_n994));
  AOI21_X1  g808(.A(G953), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n986), .B1(new_n995), .B2(new_n690), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n732), .A2(new_n988), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(KEYINPUT62), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT122), .ZN(new_n999));
  OR2_X1    g813(.A1(new_n997), .A2(KEYINPUT62), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n839), .B1(new_n377), .B2(new_n408), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n555), .B1(new_n1001), .B2(KEYINPUT123), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n771), .A2(new_n619), .A3(new_n715), .ZN(new_n1003));
  AOI211_X1 g817(.A(new_n1002), .B(new_n1003), .C1(KEYINPUT123), .C2(new_n1001), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n810), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n999), .A2(new_n817), .A3(new_n1000), .A4(new_n1005), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n1006), .A2(new_n251), .ZN(new_n1007));
  OR2_X1    g821(.A1(new_n1007), .A2(new_n986), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n251), .B1(G227), .B2(G900), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1009), .B(KEYINPUT124), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n996), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1010), .B1(new_n996), .B2(new_n1008), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1011), .A2(new_n1012), .ZN(G72));
  NAND2_X1  g827(.A1(new_n499), .A2(new_n530), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n992), .A2(new_n994), .A3(new_n865), .ZN(new_n1015));
  XOR2_X1   g829(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1016));
  NAND2_X1  g830(.A1(G472), .A2(G902), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1014), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1018), .B1(new_n1006), .B2(new_n982), .ZN(new_n1020));
  AND2_X1   g834(.A1(new_n1020), .A2(new_n721), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n722), .A2(new_n1014), .A3(new_n1018), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT127), .Z(new_n1023));
  NOR2_X1   g837(.A1(new_n921), .A2(new_n1023), .ZN(new_n1024));
  NOR4_X1   g838(.A1(new_n1019), .A2(new_n1021), .A3(new_n947), .A4(new_n1024), .ZN(G57));
endmodule


