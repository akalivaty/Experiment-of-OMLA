//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n797, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929;
  INV_X1    g000(.A(G50gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G43gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT86), .ZN(new_n204));
  AOI21_X1  g003(.A(KEYINPUT15), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G43gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G50gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G29gat), .ZN(new_n210));
  INV_X1    g009(.A(G36gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT14), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT14), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(G29gat), .A2(G36gat), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n212), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n203), .B(new_n207), .C1(new_n204), .C2(KEYINPUT15), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n209), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n203), .A2(new_n207), .A3(KEYINPUT15), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT85), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n212), .A2(new_n214), .A3(new_n215), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n220), .B1(new_n219), .B2(new_n221), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n218), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(KEYINPUT87), .B(KEYINPUT17), .Z(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G15gat), .B(G22gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n228), .A2(G1gat), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n227), .A2(G1gat), .ZN(new_n231));
  OAI21_X1  g030(.A(G8gat), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n227), .A2(new_n229), .ZN(new_n233));
  INV_X1    g032(.A(G8gat), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n233), .B(new_n234), .C1(G1gat), .C2(new_n227), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  OAI211_X1 g036(.A(KEYINPUT17), .B(new_n218), .C1(new_n222), .C2(new_n223), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n226), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n224), .A2(new_n236), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT88), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G229gat), .A2(G233gat), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n226), .A2(new_n241), .A3(new_n237), .A4(new_n238), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT18), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n224), .B(new_n236), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n244), .B(KEYINPUT13), .Z(new_n250));
  AND2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n246), .A2(KEYINPUT89), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT89), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n243), .A2(new_n254), .A3(new_n244), .A4(new_n245), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n253), .A2(new_n247), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G169gat), .B(G197gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G113gat), .B(G141gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT12), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT90), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n256), .A2(new_n265), .ZN(new_n266));
  NOR3_X1   g065(.A1(new_n248), .A2(new_n251), .A3(new_n263), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n253), .A2(KEYINPUT90), .A3(new_n247), .A4(new_n255), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT91), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT91), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n266), .A2(new_n271), .A3(new_n267), .A4(new_n268), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n264), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT92), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G57gat), .ZN(new_n277));
  INV_X1    g076(.A(G64gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G57gat), .A2(G64gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n276), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(G71gat), .B(G78gat), .Z(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n280), .A2(KEYINPUT93), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n278), .B1(new_n277), .B2(KEYINPUT93), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n276), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT94), .B(KEYINPUT21), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT21), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n237), .B1(new_n288), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G183gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n294), .A2(G183gat), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n292), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n297), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n299), .A2(new_n295), .A3(new_n291), .ZN(new_n300));
  XNOR2_X1  g099(.A(G127gat), .B(G155gat), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n301), .B(KEYINPUT20), .Z(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  AND3_X1   g102(.A1(new_n298), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n303), .B1(new_n298), .B2(new_n300), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(G211gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(G231gat), .A2(G233gat), .ZN(new_n308));
  XOR2_X1   g107(.A(new_n307), .B(new_n308), .Z(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  OR3_X1    g109(.A1(new_n304), .A2(new_n305), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n304), .B2(new_n305), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(G99gat), .B(G106gat), .Z(new_n314));
  NAND2_X1  g113(.A1(G85gat), .A2(G92gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(KEYINPUT7), .ZN(new_n316));
  NAND2_X1  g115(.A1(G99gat), .A2(G106gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT8), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT96), .ZN(new_n319));
  OR2_X1    g118(.A1(G85gat), .A2(G92gat), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n319), .B1(new_n318), .B2(new_n320), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n316), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT97), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT97), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n325), .B(new_n316), .C1(new_n321), .C2(new_n322), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n314), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n324), .A2(new_n314), .A3(new_n326), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(KEYINPUT98), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT98), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n324), .A2(new_n314), .A3(new_n326), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n331), .B1(new_n332), .B2(new_n327), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n330), .A2(new_n333), .A3(new_n238), .A4(new_n226), .ZN(new_n334));
  NAND3_X1  g133(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n328), .A2(new_n224), .A3(new_n329), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G134gat), .B(G162gat), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n338), .B(KEYINPUT99), .Z(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G190gat), .B(G218gat), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n341), .B(new_n342), .Z(new_n343));
  INV_X1    g142(.A(new_n339), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n334), .A2(new_n344), .A3(new_n335), .A4(new_n336), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n340), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n343), .B1(new_n340), .B2(new_n345), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n313), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n328), .A2(new_n289), .A3(new_n329), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n288), .B1(new_n332), .B2(new_n327), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT10), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n328), .A2(KEYINPUT10), .A3(new_n289), .A4(new_n329), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G230gat), .ZN(new_n357));
  INV_X1    g156(.A(G233gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G120gat), .B(G148gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(G176gat), .B(G204gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  AND2_X1   g164(.A1(new_n351), .A2(new_n352), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n361), .B(new_n365), .C1(new_n366), .C2(new_n360), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT100), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n366), .A2(new_n360), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n359), .B1(new_n354), .B2(new_n355), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n364), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  OAI211_X1 g171(.A(KEYINPUT100), .B(new_n364), .C1(new_n369), .C2(new_n370), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n350), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT101), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT101), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n350), .A2(new_n377), .A3(new_n374), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT83), .ZN(new_n380));
  NAND2_X1  g179(.A1(G228gat), .A2(G233gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(G155gat), .A2(G162gat), .ZN(new_n382));
  INV_X1    g181(.A(G155gat), .ZN(new_n383));
  INV_X1    g182(.A(G162gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  XOR2_X1   g184(.A(KEYINPUT74), .B(KEYINPUT2), .Z(new_n386));
  XNOR2_X1  g185(.A(G141gat), .B(G148gat), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n382), .B(new_n385), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n387), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n382), .B1(new_n385), .B2(KEYINPUT2), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT22), .ZN(new_n393));
  INV_X1    g192(.A(G211gat), .ZN(new_n394));
  INV_X1    g193(.A(G218gat), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT72), .ZN(new_n397));
  XNOR2_X1  g196(.A(G197gat), .B(G204gat), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT72), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n399), .B(new_n393), .C1(new_n394), .C2(new_n395), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n397), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G211gat), .B(G218gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n403), .A2(KEYINPUT29), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n392), .B1(new_n404), .B2(KEYINPUT3), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n392), .A2(KEYINPUT3), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n403), .B1(new_n406), .B2(KEYINPUT29), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(G22gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n408), .A2(G22gat), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n381), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OR2_X1    g211(.A1(new_n408), .A2(G22gat), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n413), .A2(G228gat), .A3(G233gat), .A4(new_n409), .ZN(new_n414));
  XNOR2_X1  g213(.A(G78gat), .B(G106gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT31), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT76), .B(G50gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n412), .A2(new_n414), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT79), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT79), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n412), .A2(new_n414), .A3(new_n421), .A4(new_n418), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n412), .A2(new_n414), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n418), .B(KEYINPUT77), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT78), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n424), .A2(KEYINPUT78), .A3(new_n425), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n423), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT25), .ZN(new_n429));
  INV_X1    g228(.A(G169gat), .ZN(new_n430));
  INV_X1    g229(.A(G176gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(G169gat), .A2(G176gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT23), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT23), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n436), .B1(G169gat), .B2(G176gat), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT24), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n439), .A2(G183gat), .A3(G190gat), .ZN(new_n440));
  INV_X1    g239(.A(G183gat), .ZN(new_n441));
  INV_X1    g240(.A(G190gat), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT24), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(G183gat), .A2(G190gat), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n440), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n429), .B1(new_n438), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT64), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n429), .B1(new_n432), .B2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n434), .B(KEYINPUT65), .ZN(new_n449));
  OAI221_X1 g248(.A(new_n448), .B1(new_n445), .B2(KEYINPUT66), .C1(new_n436), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(KEYINPUT66), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n451), .B(new_n437), .C1(new_n447), .C2(new_n432), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n446), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT27), .B(G183gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n442), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT67), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n456), .A2(KEYINPUT28), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n455), .B(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n433), .B(new_n459), .C1(new_n449), .C2(KEYINPUT26), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n458), .B(new_n460), .C1(new_n441), .C2(new_n442), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n453), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(G113gat), .B(G120gat), .Z(new_n463));
  INV_X1    g262(.A(KEYINPUT1), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G127gat), .B(G134gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT69), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n463), .A2(new_n464), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT68), .B(G134gat), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n471), .A2(G127gat), .ZN(new_n472));
  INV_X1    g271(.A(G134gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n473), .A2(G127gat), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n470), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n465), .A2(KEYINPUT69), .A3(new_n466), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n469), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n477), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n469), .A2(new_n475), .A3(new_n476), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n479), .A2(new_n453), .A3(new_n461), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(G227gat), .A2(G233gat), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT33), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT70), .B(G71gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(G99gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(G15gat), .B(G43gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n481), .A2(KEYINPUT34), .A3(new_n483), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT34), .B1(new_n481), .B2(new_n483), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n484), .A2(KEYINPUT32), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n495), .B1(new_n493), .B2(new_n494), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n491), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n498), .ZN(new_n500));
  INV_X1    g299(.A(new_n491), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(new_n496), .A3(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT6), .ZN(new_n504));
  INV_X1    g303(.A(new_n392), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n477), .B(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G225gat), .A2(G233gat), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n479), .A2(new_n505), .ZN(new_n509));
  INV_X1    g308(.A(new_n406), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n392), .A2(KEYINPUT3), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n477), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n509), .A2(KEYINPUT4), .A3(new_n512), .ZN(new_n513));
  OR3_X1    g312(.A1(new_n477), .A2(KEYINPUT4), .A3(new_n392), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n507), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT4), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n508), .A2(new_n518), .A3(KEYINPUT5), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT5), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n515), .A2(new_n520), .A3(new_n507), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G57gat), .B(G85gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT75), .B(KEYINPUT0), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G1gat), .B(G29gat), .ZN(new_n526));
  XOR2_X1   g325(.A(new_n525), .B(new_n526), .Z(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n504), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n522), .A2(new_n528), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT81), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n522), .A2(KEYINPUT81), .A3(new_n528), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n529), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n530), .A2(new_n504), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n428), .B(new_n503), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(G226gat), .A2(G233gat), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n462), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(KEYINPUT29), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n539), .B1(new_n453), .B2(new_n461), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n538), .A2(new_n403), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G8gat), .B(G36gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(G64gat), .B(G92gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n403), .B1(new_n538), .B2(new_n540), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n542), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT73), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT30), .ZN(new_n551));
  INV_X1    g350(.A(new_n547), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n545), .B1(new_n552), .B2(new_n541), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n548), .A2(new_n549), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n551), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n556), .A2(KEYINPUT35), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n380), .B1(new_n536), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n529), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n530), .ZN(new_n561));
  INV_X1    g360(.A(new_n535), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n556), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n428), .A2(new_n503), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT35), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n532), .A2(new_n533), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n560), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(new_n562), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n424), .A2(new_n425), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT78), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n424), .A2(KEYINPUT78), .A3(new_n425), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n573), .A2(new_n574), .B1(new_n420), .B2(new_n422), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n499), .A2(new_n502), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n570), .A2(new_n577), .A3(KEYINPUT83), .A4(new_n557), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n559), .A2(new_n567), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n576), .A2(KEYINPUT71), .A3(KEYINPUT36), .ZN(new_n580));
  NAND2_X1  g379(.A1(KEYINPUT71), .A2(KEYINPUT36), .ZN(new_n581));
  OR2_X1    g380(.A1(KEYINPUT71), .A2(KEYINPUT36), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n499), .A2(new_n502), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n565), .A2(new_n575), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT82), .B(KEYINPUT38), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n548), .A2(new_n586), .ZN(new_n587));
  OR3_X1    g386(.A1(new_n552), .A2(KEYINPUT37), .A3(new_n541), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT37), .B1(new_n552), .B2(new_n541), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(new_n545), .A3(new_n589), .ZN(new_n590));
  MUX2_X1   g389(.A(new_n586), .B(new_n587), .S(new_n590), .Z(new_n591));
  NOR2_X1   g390(.A1(new_n570), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n513), .A2(new_n516), .A3(new_n514), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n593), .A2(KEYINPUT80), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(KEYINPUT80), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n506), .A2(new_n507), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n594), .A2(KEYINPUT39), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n594), .A2(new_n595), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n527), .B(new_n597), .C1(new_n598), .C2(KEYINPUT39), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT40), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n568), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n556), .B1(new_n599), .B2(new_n600), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n428), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n584), .B(new_n585), .C1(new_n592), .C2(new_n604), .ZN(new_n605));
  AOI211_X1 g404(.A(new_n273), .B(new_n379), .C1(new_n579), .C2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n563), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(G1gat), .ZN(G1324gat));
  INV_X1    g408(.A(new_n606), .ZN(new_n610));
  OAI21_X1  g409(.A(G8gat), .B1(new_n610), .B2(new_n564), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT42), .ZN(new_n612));
  NAND2_X1  g411(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n228), .A2(new_n234), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n606), .A2(new_n556), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n615), .A2(KEYINPUT102), .A3(new_n612), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT102), .B1(new_n615), .B2(new_n612), .ZN(new_n618));
  OAI221_X1 g417(.A(new_n611), .B1(new_n612), .B2(new_n615), .C1(new_n617), .C2(new_n618), .ZN(G1325gat));
  INV_X1    g418(.A(new_n584), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n606), .A2(G15gat), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n503), .ZN(new_n622));
  INV_X1    g421(.A(G15gat), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n622), .A2(KEYINPUT103), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT103), .B1(new_n622), .B2(new_n623), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT104), .ZN(G1326gat));
  NAND2_X1  g426(.A1(new_n606), .A2(new_n575), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT43), .B(G22gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(G1327gat));
  INV_X1    g429(.A(new_n374), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n631), .A2(KEYINPUT105), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(KEYINPUT105), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n313), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT107), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(new_n347), .B2(new_n348), .ZN(new_n639));
  INV_X1    g438(.A(new_n348), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n640), .A2(KEYINPUT107), .A3(new_n346), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(KEYINPUT44), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT106), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n579), .A2(new_n644), .A3(new_n605), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n644), .B1(new_n579), .B2(new_n605), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n579), .A2(new_n605), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n349), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT44), .ZN(new_n650));
  AOI211_X1 g449(.A(new_n273), .B(new_n637), .C1(new_n647), .C2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n210), .B1(new_n651), .B2(new_n607), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n273), .B1(new_n579), .B2(new_n605), .ZN(new_n653));
  INV_X1    g452(.A(new_n349), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n635), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n653), .A2(new_n607), .A3(new_n374), .A4(new_n655), .ZN(new_n656));
  OR3_X1    g455(.A1(new_n656), .A2(KEYINPUT45), .A3(G29gat), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT45), .B1(new_n656), .B2(G29gat), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT108), .B1(new_n652), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n647), .A2(new_n650), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n270), .A2(new_n272), .ZN(new_n663));
  INV_X1    g462(.A(new_n264), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n662), .A2(new_n665), .A3(new_n636), .ZN(new_n666));
  OAI21_X1  g465(.A(G29gat), .B1(new_n666), .B2(new_n563), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(new_n668), .A3(new_n659), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n661), .A2(new_n669), .ZN(G1328gat));
  INV_X1    g469(.A(KEYINPUT109), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n211), .B1(new_n651), .B2(new_n556), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n648), .A2(new_n665), .A3(new_n374), .A4(new_n655), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n673), .A2(G36gat), .A3(new_n564), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT46), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n671), .B1(new_n672), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(G36gat), .B1(new_n666), .B2(new_n564), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n674), .B(KEYINPUT46), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n678), .A2(KEYINPUT109), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n677), .A2(new_n680), .ZN(G1329gat));
  INV_X1    g480(.A(KEYINPUT47), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n662), .A2(new_n665), .A3(new_n620), .A4(new_n636), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(G43gat), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n673), .A2(G43gat), .A3(new_n576), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n682), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  AOI211_X1 g486(.A(KEYINPUT47), .B(new_n685), .C1(new_n683), .C2(G43gat), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(G1330gat));
  OAI21_X1  g488(.A(new_n202), .B1(new_n673), .B2(new_n428), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n575), .A2(G50gat), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n690), .B1(new_n666), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g492(.A1(new_n634), .A2(new_n350), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n273), .B(new_n694), .C1(new_n645), .C2(new_n646), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n563), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(new_n277), .ZN(G1332gat));
  NOR2_X1   g496(.A1(new_n695), .A2(new_n564), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT49), .B(G64gat), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n700), .B1(new_n698), .B2(new_n701), .ZN(G1333gat));
  INV_X1    g501(.A(KEYINPUT50), .ZN(new_n703));
  OAI21_X1  g502(.A(G71gat), .B1(new_n695), .B2(new_n584), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n648), .A2(KEYINPUT106), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n579), .A2(new_n605), .A3(new_n644), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n665), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(G71gat), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n707), .A2(new_n708), .A3(new_n503), .A4(new_n694), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT110), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n704), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n710), .B1(new_n704), .B2(new_n709), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n703), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n704), .A2(new_n709), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT110), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n716), .A2(KEYINPUT50), .A3(new_n711), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n714), .A2(new_n717), .ZN(G1334gat));
  NOR2_X1   g517(.A1(new_n695), .A2(new_n428), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(G78gat), .Z(G1335gat));
  INV_X1    g519(.A(KEYINPUT111), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n665), .A2(new_n635), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n662), .A2(new_n631), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n723), .B2(new_n563), .ZN(new_n724));
  INV_X1    g523(.A(new_n722), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n647), .B2(new_n650), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n726), .A2(KEYINPUT111), .A3(new_n607), .A4(new_n631), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n724), .A2(G85gat), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n648), .A2(new_n349), .A3(new_n722), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT51), .ZN(new_n730));
  OR2_X1    g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT112), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n730), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n729), .A2(KEYINPUT112), .A3(new_n730), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n734), .A2(new_n631), .A3(new_n735), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n563), .A2(G85gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n728), .B1(new_n736), .B2(new_n737), .ZN(G1336gat));
  NAND3_X1  g537(.A1(new_n726), .A2(new_n556), .A3(new_n631), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G92gat), .ZN(new_n740));
  INV_X1    g539(.A(new_n634), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n741), .A2(G92gat), .A3(new_n564), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n734), .A2(new_n735), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT52), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n740), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n731), .A2(new_n733), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n739), .A2(G92gat), .B1(new_n746), .B2(new_n742), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n747), .B2(new_n744), .ZN(G1337gat));
  OAI21_X1  g547(.A(G99gat), .B1(new_n723), .B2(new_n584), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n576), .A2(G99gat), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n736), .B2(new_n750), .ZN(G1338gat));
  NAND3_X1  g550(.A1(new_n726), .A2(new_n575), .A3(new_n631), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G106gat), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n741), .A2(G106gat), .A3(new_n428), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n734), .A2(new_n735), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n753), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  AOI22_X1  g556(.A1(new_n752), .A2(G106gat), .B1(new_n746), .B2(new_n754), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n758), .B2(new_n756), .ZN(G1339gat));
  NOR2_X1   g558(.A1(new_n375), .A2(new_n665), .ZN(new_n760));
  INV_X1    g559(.A(new_n262), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n244), .B1(new_n243), .B2(new_n245), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n249), .A2(new_n250), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n663), .A2(new_n631), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT113), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n354), .A2(new_n355), .A3(new_n359), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n361), .A2(KEYINPUT54), .A3(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT54), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n365), .B1(new_n370), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n768), .A2(KEYINPUT55), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n367), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT55), .B1(new_n768), .B2(new_n770), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n766), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n356), .A2(new_n769), .A3(new_n360), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n767), .A2(KEYINPUT54), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n364), .B(new_n775), .C1(new_n776), .C2(new_n370), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n779), .A2(new_n771), .A3(KEYINPUT113), .A4(new_n367), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n774), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n765), .B1(new_n781), .B2(new_n273), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n642), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n663), .A2(new_n764), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(new_n642), .ZN(new_n785));
  INV_X1    g584(.A(new_n781), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n760), .B1(new_n788), .B2(new_n313), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n566), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n563), .A2(new_n556), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n665), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(G113gat), .ZN(G1340gat));
  OAI21_X1  g594(.A(G120gat), .B1(new_n792), .B2(new_n741), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n792), .A2(G120gat), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n797), .B2(new_n374), .ZN(G1341gat));
  NAND2_X1  g597(.A1(new_n793), .A2(new_n635), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g599(.A1(new_n564), .A2(new_n349), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT114), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n790), .A2(new_n471), .A3(new_n607), .A4(new_n802), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n803), .B(KEYINPUT56), .Z(new_n804));
  OAI21_X1  g603(.A(G134gat), .B1(new_n792), .B2(new_n654), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(G1343gat));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n807));
  INV_X1    g606(.A(new_n642), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n665), .A2(new_n774), .A3(new_n780), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(new_n809), .B2(new_n765), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n781), .A2(new_n784), .A3(new_n642), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n313), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n760), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n428), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n807), .B1(new_n814), .B2(KEYINPUT57), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n777), .A2(KEYINPUT116), .A3(new_n778), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT116), .B1(new_n777), .B2(new_n778), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n273), .A2(new_n818), .A3(new_n772), .ZN(new_n819));
  INV_X1    g618(.A(new_n765), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n654), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n635), .B1(new_n821), .B2(new_n787), .ZN(new_n822));
  OAI211_X1 g621(.A(KEYINPUT57), .B(new_n575), .C1(new_n822), .C2(new_n760), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824));
  OAI211_X1 g623(.A(KEYINPUT115), .B(new_n824), .C1(new_n789), .C2(new_n428), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n815), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n584), .A2(new_n791), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n665), .A3(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(G141gat), .ZN(new_n830));
  OR2_X1    g629(.A1(new_n273), .A2(G141gat), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n814), .A2(new_n584), .A3(new_n791), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n831), .A2(new_n832), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT118), .ZN(new_n839));
  OAI21_X1  g638(.A(KEYINPUT58), .B1(new_n830), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n829), .A2(G141gat), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n842), .B1(new_n835), .B2(new_n837), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n782), .A2(new_n642), .B1(new_n785), .B2(new_n786), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n813), .B1(new_n845), .B2(new_n635), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n846), .A2(new_n575), .A3(new_n584), .A4(new_n791), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n848), .A2(KEYINPUT119), .A3(new_n836), .A4(new_n834), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n843), .A2(new_n844), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n841), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n841), .A2(new_n850), .A3(KEYINPUT120), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n840), .A2(new_n853), .A3(new_n854), .ZN(G1344gat));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n826), .A2(new_n828), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n856), .B(G148gat), .C1(new_n857), .C2(new_n374), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n827), .A2(KEYINPUT121), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n584), .A2(new_n860), .A3(new_n791), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n374), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n428), .A2(KEYINPUT57), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n654), .A2(new_n772), .A3(new_n773), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n663), .A3(new_n764), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n635), .B1(new_n821), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n379), .A2(new_n665), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n863), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n862), .B(new_n868), .C1(new_n814), .C2(new_n824), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT122), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n846), .A2(new_n575), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT57), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n872), .A2(new_n873), .A3(new_n868), .A4(new_n862), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n870), .A2(new_n874), .A3(G148gat), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n875), .A2(new_n876), .A3(KEYINPUT59), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n876), .B1(new_n875), .B2(KEYINPUT59), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n858), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OR3_X1    g678(.A1(new_n847), .A2(G148gat), .A3(new_n374), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1345gat));
  NOR3_X1   g680(.A1(new_n857), .A2(new_n383), .A3(new_n313), .ZN(new_n882));
  AOI21_X1  g681(.A(G155gat), .B1(new_n848), .B2(new_n635), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(G1346gat));
  OAI21_X1  g683(.A(G162gat), .B1(new_n857), .B2(new_n642), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n871), .A2(new_n620), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n384), .A3(new_n802), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n885), .B1(new_n563), .B2(new_n887), .ZN(G1347gat));
  NOR2_X1   g687(.A1(new_n607), .A2(new_n564), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT124), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n790), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(G169gat), .B1(new_n892), .B2(new_n273), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n790), .A2(new_n889), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n430), .A3(new_n665), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n893), .A2(new_n896), .ZN(G1348gat));
  OAI21_X1  g696(.A(new_n431), .B1(new_n894), .B2(new_n374), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT125), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n892), .A2(new_n431), .A3(new_n741), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(G1349gat));
  OAI21_X1  g700(.A(G183gat), .B1(new_n892), .B2(new_n313), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n895), .A2(new_n454), .A3(new_n635), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(KEYINPUT126), .A3(new_n903), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g704(.A(new_n442), .B1(new_n891), .B2(new_n349), .ZN(new_n906));
  XOR2_X1   g705(.A(new_n906), .B(KEYINPUT61), .Z(new_n907));
  NAND3_X1  g706(.A1(new_n895), .A2(new_n442), .A3(new_n808), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1351gat));
  NAND4_X1  g708(.A1(new_n872), .A2(new_n584), .A3(new_n868), .A4(new_n890), .ZN(new_n910));
  OAI21_X1  g709(.A(G197gat), .B1(new_n910), .B2(new_n273), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n886), .A2(new_n889), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n273), .A2(G197gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(G1352gat));
  NOR2_X1   g713(.A1(new_n910), .A2(new_n741), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n915), .A2(KEYINPUT127), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(KEYINPUT127), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n916), .A2(G204gat), .A3(new_n917), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n912), .A2(G204gat), .A3(new_n374), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT62), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1353gat));
  OR2_X1    g720(.A1(new_n910), .A2(new_n313), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT63), .B1(new_n922), .B2(G211gat), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n635), .A2(new_n394), .ZN(new_n926));
  OAI22_X1  g725(.A1(new_n924), .A2(new_n925), .B1(new_n912), .B2(new_n926), .ZN(G1354gat));
  OAI21_X1  g726(.A(G218gat), .B1(new_n910), .B2(new_n654), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n808), .A2(new_n395), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n912), .B2(new_n929), .ZN(G1355gat));
endmodule


