//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(G146), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT64), .A3(G143), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n193), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n197));
  XOR2_X1   g011(.A(KEYINPUT0), .B(G128), .Z(new_n198));
  AND3_X1   g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n197), .B1(new_n196), .B2(new_n198), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n194), .A2(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(new_n193), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT0), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NOR3_X1   g018(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NOR3_X1   g019(.A1(new_n199), .A2(new_n200), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT3), .B1(new_n207), .B2(G107), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G104), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n208), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(KEYINPUT79), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT4), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n208), .A2(new_n211), .A3(new_n214), .A4(new_n212), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n213), .A2(KEYINPUT4), .A3(new_n215), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n206), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT10), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n224));
  AND4_X1   g038(.A1(new_n224), .A2(new_n201), .A3(new_n193), .A4(G128), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT1), .B1(new_n191), .B2(G146), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT80), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n201), .A2(KEYINPUT80), .A3(KEYINPUT1), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(G128), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n225), .B1(new_n230), .B2(new_n202), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n210), .A2(G104), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n207), .A2(G107), .ZN(new_n233));
  OAI21_X1  g047(.A(G101), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n219), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n223), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n225), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n226), .A2(G128), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n196), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT81), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n219), .A2(new_n234), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n241), .B1(new_n219), .B2(new_n234), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n240), .B(KEYINPUT10), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n222), .A2(new_n236), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT11), .ZN(new_n246));
  INV_X1    g060(.A(G134), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n246), .B1(new_n247), .B2(G137), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(G137), .ZN(new_n249));
  INV_X1    g063(.A(G137), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(KEYINPUT11), .A3(G134), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G131), .ZN(new_n253));
  INV_X1    g067(.A(G131), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n248), .A2(new_n251), .A3(new_n254), .A4(new_n249), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n245), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n256), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n222), .A2(new_n258), .A3(new_n236), .A4(new_n244), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g074(.A(G110), .B(G140), .Z(new_n261));
  INV_X1    g075(.A(G227), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(G953), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n261), .B(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT83), .B1(new_n260), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n264), .B1(new_n257), .B2(new_n259), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT83), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n259), .A2(new_n264), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT12), .ZN(new_n271));
  INV_X1    g085(.A(new_n243), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n225), .B1(new_n196), .B2(new_n238), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n219), .A2(new_n234), .A3(new_n241), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n235), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n224), .B1(G143), .B2(new_n194), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n204), .B1(new_n277), .B2(KEYINPUT80), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n278), .A2(new_n228), .B1(new_n201), .B2(new_n193), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n276), .B1(new_n279), .B2(new_n225), .ZN(new_n280));
  AOI211_X1 g094(.A(new_n271), .B(new_n258), .C1(new_n275), .C2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n275), .A2(new_n280), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT12), .B1(new_n282), .B2(new_n256), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n270), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n265), .A2(new_n268), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G902), .ZN(new_n286));
  INV_X1    g100(.A(G469), .ZN(new_n287));
  OR2_X1    g101(.A1(new_n287), .A2(KEYINPUT82), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(KEYINPUT82), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n285), .A2(new_n286), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n259), .B1(new_n283), .B2(new_n281), .ZN(new_n291));
  XOR2_X1   g105(.A(new_n264), .B(KEYINPUT78), .Z(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n270), .A2(new_n257), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G469), .B1(new_n296), .B2(G902), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n189), .B1(new_n290), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(G475), .A2(G902), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n299), .B(KEYINPUT94), .ZN(new_n300));
  XOR2_X1   g114(.A(G113), .B(G122), .Z(new_n301));
  XNOR2_X1  g115(.A(new_n301), .B(KEYINPUT92), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(G104), .ZN(new_n303));
  INV_X1    g117(.A(G140), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G125), .ZN(new_n305));
  INV_X1    g119(.A(G125), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G140), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT90), .B1(new_n308), .B2(KEYINPUT19), .ZN(new_n309));
  NOR3_X1   g123(.A1(new_n306), .A2(KEYINPUT74), .A3(G140), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n305), .A2(new_n307), .A3(KEYINPUT74), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT19), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n309), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(G125), .B(G140), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n310), .B1(new_n316), .B2(KEYINPUT74), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(KEYINPUT90), .A3(KEYINPUT19), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n318), .A3(new_n194), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n313), .A2(KEYINPUT16), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT75), .B1(new_n305), .B2(KEYINPUT16), .ZN(new_n321));
  OR3_X1    g135(.A1(new_n305), .A2(KEYINPUT75), .A3(KEYINPUT16), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n320), .A2(G146), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT91), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT91), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n319), .A2(new_n326), .A3(new_n323), .ZN(new_n327));
  NOR2_X1   g141(.A1(G237), .A2(G953), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(G143), .A3(G214), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(G143), .B1(new_n328), .B2(G214), .ZN(new_n331));
  OAI21_X1  g145(.A(G131), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n331), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(new_n254), .A3(new_n329), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n325), .A2(new_n327), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n316), .A2(new_n194), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n337), .B1(new_n313), .B2(new_n194), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n330), .A2(new_n331), .ZN(new_n339));
  AND4_X1   g153(.A1(KEYINPUT89), .A2(new_n339), .A3(KEYINPUT18), .A4(G131), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n339), .A2(KEYINPUT89), .B1(KEYINPUT18), .B2(G131), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n338), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n303), .B1(new_n336), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT17), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n332), .A2(new_n334), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT93), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT16), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n321), .B(new_n322), .C1(new_n317), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n194), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n350), .B(new_n323), .C1(new_n344), .C2(new_n332), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n342), .B(new_n303), .C1(new_n347), .C2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n300), .B1(new_n343), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT20), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n327), .A2(new_n335), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n326), .B1(new_n319), .B2(new_n323), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n342), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n303), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n352), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT20), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n300), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n355), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n342), .B1(new_n347), .B2(new_n351), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n365), .A2(new_n359), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n286), .B1(new_n366), .B2(new_n353), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G475), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT96), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT95), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n191), .A2(G128), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n204), .A2(G143), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n371), .A2(new_n372), .A3(new_n247), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n247), .B1(new_n371), .B2(new_n372), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n370), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n371), .A2(new_n372), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G134), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n371), .A2(new_n372), .A3(new_n247), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(KEYINPUT95), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G116), .B(G122), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n210), .ZN(new_n381));
  INV_X1    g195(.A(G122), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G116), .ZN(new_n383));
  INV_X1    g197(.A(G116), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G122), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT14), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n387), .B(G107), .C1(new_n386), .C2(new_n385), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n375), .A2(new_n379), .A3(new_n381), .A4(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n380), .B(new_n210), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT13), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n391), .B(G134), .C1(KEYINPUT13), .C2(new_n371), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n392), .A3(new_n378), .ZN(new_n393));
  INV_X1    g207(.A(G217), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n187), .A2(new_n394), .A3(G953), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n389), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n395), .B1(new_n389), .B2(new_n393), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n369), .B1(new_n398), .B2(G902), .ZN(new_n399));
  INV_X1    g213(.A(G478), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(KEYINPUT15), .ZN(new_n401));
  OAI211_X1 g215(.A(KEYINPUT96), .B(new_n286), .C1(new_n396), .C2(new_n397), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  OR3_X1    g217(.A1(new_n398), .A2(G902), .A3(new_n401), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n364), .A2(new_n368), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G214), .B1(G237), .B2(G902), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G953), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n411), .A2(G952), .ZN(new_n412));
  NAND2_X1  g226(.A1(G234), .A2(G237), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  XOR2_X1   g228(.A(new_n414), .B(KEYINPUT97), .Z(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT21), .B(G898), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n413), .A2(G902), .A3(G953), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n416), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(G210), .B1(G237), .B2(G902), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(KEYINPUT88), .ZN(new_n422));
  INV_X1    g236(.A(G224), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(G953), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n196), .A2(new_n198), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT65), .ZN(new_n426));
  INV_X1    g240(.A(new_n205), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n196), .A2(new_n198), .A3(new_n197), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(KEYINPUT84), .A3(G125), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n237), .A2(new_n239), .A3(new_n306), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n429), .A2(G125), .B1(KEYINPUT84), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n424), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(KEYINPUT84), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n435), .B1(new_n206), .B2(new_n306), .ZN(new_n436));
  INV_X1    g250(.A(new_n424), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(new_n437), .A3(new_n430), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT2), .B(G113), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(G116), .B(G119), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n442), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n221), .A2(new_n445), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n384), .A2(KEYINPUT5), .A3(G119), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n442), .B2(KEYINPUT5), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n448), .A2(G113), .B1(new_n442), .B2(new_n441), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n449), .B1(new_n242), .B2(new_n243), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G110), .B(G122), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n446), .A2(new_n452), .A3(new_n450), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(KEYINPUT6), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT6), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n451), .A2(new_n457), .A3(new_n453), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n439), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n286), .ZN(new_n460));
  XOR2_X1   g274(.A(KEYINPUT86), .B(KEYINPUT7), .Z(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n436), .A2(new_n430), .B1(new_n437), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(KEYINPUT87), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n436), .A2(KEYINPUT7), .A3(new_n437), .A4(new_n430), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT85), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n449), .B2(new_n276), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n442), .A2(KEYINPUT5), .ZN(new_n468));
  INV_X1    g282(.A(new_n447), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(G113), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n444), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(KEYINPUT85), .A3(new_n235), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n467), .A2(new_n472), .A3(new_n450), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n452), .B(KEYINPUT8), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n465), .A2(new_n455), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT87), .ZN(new_n477));
  AOI221_X4 g291(.A(new_n477), .B1(new_n437), .B2(new_n462), .C1(new_n436), .C2(new_n430), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n464), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n422), .B1(new_n460), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n461), .B1(new_n431), .B2(new_n433), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n434), .A2(new_n481), .A3(new_n477), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n465), .A2(new_n455), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n463), .A2(KEYINPUT87), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n482), .A2(new_n483), .A3(new_n475), .A4(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n422), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n485), .A2(new_n459), .A3(new_n286), .A4(new_n486), .ZN(new_n487));
  AOI211_X1 g301(.A(new_n410), .B(new_n420), .C1(new_n480), .C2(new_n487), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n298), .A2(new_n408), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n255), .A2(KEYINPUT66), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n250), .A2(G134), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n254), .B1(new_n249), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(KEYINPUT66), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n240), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n256), .A2(new_n426), .A3(new_n427), .A4(new_n428), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT68), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n199), .A2(new_n200), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n501), .A2(KEYINPUT68), .A3(new_n256), .A4(new_n427), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n497), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n445), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n504), .B1(new_n498), .B2(new_n496), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT70), .ZN(new_n507));
  OR2_X1    g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n507), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n505), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT28), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT28), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n498), .A2(new_n496), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n512), .B1(new_n513), .B2(new_n445), .ZN(new_n514));
  XOR2_X1   g328(.A(KEYINPUT26), .B(G101), .Z(new_n515));
  NAND2_X1  g329(.A1(new_n328), .A2(G210), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n517), .B(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n511), .A2(new_n514), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT68), .B1(new_n206), .B2(new_n256), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n498), .A2(new_n499), .ZN(new_n522));
  OAI211_X1 g336(.A(KEYINPUT30), .B(new_n496), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT30), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n513), .A2(KEYINPUT67), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT67), .B1(new_n513), .B2(new_n524), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n523), .B(new_n445), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n505), .ZN(new_n528));
  INV_X1    g342(.A(new_n519), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT29), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n520), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n505), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT71), .B1(new_n503), .B2(new_n504), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n496), .B1(new_n521), .B2(new_n522), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n445), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT71), .A3(new_n505), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n535), .A2(new_n538), .A3(KEYINPUT28), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n539), .A2(KEYINPUT29), .A3(new_n514), .A4(new_n519), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n532), .A2(new_n540), .A3(new_n286), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(G472), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n527), .A2(new_n505), .A3(new_n519), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT31), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n503), .A2(new_n504), .B1(new_n507), .B2(new_n506), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n512), .B1(new_n545), .B2(new_n508), .ZN(new_n546));
  INV_X1    g360(.A(new_n514), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n529), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT31), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n527), .A2(new_n549), .A3(new_n505), .A4(new_n519), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n544), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT32), .ZN(new_n552));
  NOR2_X1   g366(.A1(G472), .A2(G902), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n552), .B1(new_n551), .B2(new_n553), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n542), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT23), .B1(new_n204), .B2(G119), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT73), .B1(new_n204), .B2(G119), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n557), .A2(new_n558), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OR2_X1    g375(.A1(KEYINPUT24), .A2(G110), .ZN(new_n562));
  NAND2_X1  g376(.A1(KEYINPUT24), .A2(G110), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT72), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n562), .A2(KEYINPUT72), .A3(new_n563), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(G119), .B(G128), .ZN(new_n569));
  OAI22_X1  g383(.A1(new_n561), .A2(G110), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n570), .A2(new_n323), .A3(new_n337), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n350), .A2(new_n323), .ZN(new_n572));
  OAI21_X1  g386(.A(G110), .B1(new_n559), .B2(new_n560), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n566), .A2(new_n569), .A3(new_n567), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT76), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT76), .ZN(new_n578));
  AOI211_X1 g392(.A(new_n578), .B(new_n575), .C1(new_n350), .C2(new_n323), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n571), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n411), .A2(G221), .A3(G234), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT22), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(G137), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n571), .B(new_n583), .C1(new_n577), .C2(new_n579), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n286), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT25), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n394), .B1(G234), .B2(new_n286), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT25), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n585), .A2(new_n590), .A3(new_n286), .A4(new_n586), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n588), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n585), .A2(new_n586), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT77), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n589), .A2(G902), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n585), .A2(KEYINPUT77), .A3(new_n586), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n592), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n489), .A2(new_n556), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G101), .ZN(G3));
  NAND2_X1  g416(.A1(new_n551), .A2(new_n286), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(G472), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n551), .A2(new_n553), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n604), .A2(new_n600), .A3(new_n605), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n298), .A2(new_n488), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n396), .A2(new_n397), .A3(KEYINPUT33), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n389), .A2(new_n393), .ZN(new_n611));
  INV_X1    g425(.A(new_n395), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n389), .A2(new_n393), .A3(new_n395), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n610), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI211_X1 g429(.A(G478), .B(new_n286), .C1(new_n609), .C2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT98), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT33), .B1(new_n396), .B2(new_n397), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n613), .A2(new_n610), .A3(new_n614), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n622), .A2(KEYINPUT98), .A3(G478), .A4(new_n286), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n618), .A2(new_n619), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT99), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT99), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n618), .A2(new_n619), .A3(new_n626), .A4(new_n623), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n364), .A2(new_n368), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n608), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT34), .B(G104), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n355), .A2(new_n634), .A3(new_n363), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n634), .B1(new_n355), .B2(new_n363), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n368), .B(new_n405), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n608), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT35), .B(G107), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  INV_X1    g454(.A(G472), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n551), .B2(new_n286), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n551), .B2(new_n553), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n584), .A2(KEYINPUT36), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n580), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n580), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(new_n596), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n592), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n489), .A2(new_n643), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT101), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT37), .B(G110), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G12));
  INV_X1    g467(.A(G900), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n416), .B1(new_n654), .B2(new_n419), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n637), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n290), .A2(new_n297), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n410), .B1(new_n480), .B2(new_n487), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n657), .A2(new_n188), .A3(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n556), .A2(new_n656), .A3(new_n659), .A4(new_n649), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT102), .B(G128), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G30));
  INV_X1    g476(.A(new_n535), .ZN(new_n663));
  INV_X1    g477(.A(new_n538), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n529), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n528), .A2(new_n519), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n665), .A2(new_n666), .A3(new_n286), .ZN(new_n667));
  OAI22_X1  g481(.A1(new_n554), .A2(new_n555), .B1(new_n641), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n480), .A2(new_n487), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT103), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT38), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n671), .A2(KEYINPUT103), .ZN(new_n675));
  OR3_X1    g489(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n674), .B1(new_n673), .B2(new_n675), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n649), .A2(new_n410), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n406), .B1(new_n364), .B2(new_n368), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n655), .B(KEYINPUT39), .Z(new_n683));
  NAND2_X1  g497(.A1(new_n298), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT105), .B(KEYINPUT40), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(new_n686));
  OR4_X1    g500(.A1(new_n670), .A2(new_n680), .A3(new_n682), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G143), .ZN(G45));
  INV_X1    g502(.A(new_n655), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n628), .A2(new_n629), .A3(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n556), .A2(new_n659), .A3(new_n649), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G146), .ZN(G48));
  NAND2_X1  g507(.A1(new_n605), .A2(KEYINPUT32), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n599), .B1(new_n696), .B2(new_n542), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n266), .A2(new_n267), .ZN(new_n698));
  AOI211_X1 g512(.A(KEYINPUT83), .B(new_n264), .C1(new_n257), .C2(new_n259), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n283), .A2(new_n281), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n269), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n698), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(G469), .B1(new_n702), .B2(G902), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n290), .A3(new_n188), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(KEYINPUT106), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n703), .A2(new_n290), .A3(new_n706), .A4(new_n188), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n630), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n697), .A2(new_n708), .A3(new_n488), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  INV_X1    g526(.A(new_n637), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n697), .A2(new_n708), .A3(new_n488), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  AND2_X1   g529(.A1(new_n488), .A2(new_n408), .ZN(new_n716));
  INV_X1    g530(.A(new_n704), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n556), .A2(new_n716), .A3(new_n649), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n720), .B1(new_n603), .B2(G472), .ZN(new_n721));
  AOI211_X1 g535(.A(KEYINPUT107), .B(new_n641), .C1(new_n551), .C2(new_n286), .ZN(new_n722));
  INV_X1    g536(.A(new_n553), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n544), .A2(new_n550), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n539), .A2(new_n514), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n529), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n723), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n721), .A2(new_n722), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n682), .B1(new_n705), .B2(new_n707), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(new_n729), .A3(new_n600), .A4(new_n488), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  NOR2_X1   g545(.A1(new_n721), .A2(new_n722), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n658), .A2(new_n188), .A3(new_n703), .A4(new_n290), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n690), .ZN(new_n734));
  INV_X1    g548(.A(new_n727), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n732), .A2(new_n734), .A3(new_n649), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  NOR2_X1   g551(.A1(new_n671), .A2(new_n410), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n298), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n697), .A2(new_n691), .A3(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT42), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n744), .B1(new_n554), .B2(new_n555), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n694), .A2(KEYINPUT108), .A3(new_n695), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n746), .A3(new_n542), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n747), .A2(KEYINPUT42), .A3(new_n600), .A4(new_n298), .ZN(new_n748));
  INV_X1    g562(.A(new_n738), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n690), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n743), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT109), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n254), .ZN(G33));
  NAND4_X1  g568(.A1(new_n740), .A2(new_n556), .A3(new_n656), .A4(new_n600), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  NAND3_X1  g570(.A1(new_n296), .A2(KEYINPUT110), .A3(KEYINPUT45), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n287), .B1(new_n295), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n760), .B1(new_n295), .B2(new_n758), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n757), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(G469), .A2(G902), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT46), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n762), .A2(KEYINPUT46), .A3(new_n763), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n290), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n188), .A3(new_n683), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n364), .A2(new_n368), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n628), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT43), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n643), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n774), .A3(new_n649), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT44), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n769), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(KEYINPUT111), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n775), .A2(new_n780), .A3(new_n776), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n738), .B(new_n777), .C1(new_n779), .C2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G137), .ZN(G39));
  NAND3_X1  g597(.A1(new_n696), .A2(new_n599), .A3(new_n542), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n768), .A2(KEYINPUT47), .A3(new_n188), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT47), .B1(new_n768), .B2(new_n188), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n750), .B(new_n785), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(KEYINPUT49), .ZN(new_n791));
  NOR4_X1   g605(.A1(new_n678), .A2(new_n599), .A3(new_n771), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n189), .A2(new_n410), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n703), .A2(new_n290), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n790), .A2(KEYINPUT49), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n794), .B(new_n795), .Z(new_n796));
  NAND4_X1  g610(.A1(new_n792), .A2(new_n670), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  AOI211_X1 g611(.A(new_n787), .B(new_n786), .C1(new_n189), .C2(new_n794), .ZN(new_n798));
  AND4_X1   g612(.A1(new_n600), .A2(new_n773), .A3(new_n416), .A4(new_n728), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n738), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n678), .A2(new_n409), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n799), .A2(new_n717), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n749), .A2(new_n415), .A3(new_n704), .ZN(new_n806));
  AND4_X1   g620(.A1(new_n649), .A2(new_n773), .A3(new_n728), .A4(new_n806), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n670), .A2(new_n600), .A3(new_n806), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n628), .A2(new_n629), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n801), .A2(new_n805), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n801), .A2(new_n805), .A3(KEYINPUT51), .A4(new_n810), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n813), .A2(new_n412), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n799), .A2(new_n658), .A3(new_n717), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n736), .A2(new_n660), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT116), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n655), .B(KEYINPUT114), .Z(new_n819));
  NAND3_X1  g633(.A1(new_n592), .A2(new_n648), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n592), .A2(KEYINPUT115), .A3(new_n648), .A4(new_n819), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n681), .A2(new_n658), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n668), .A2(new_n824), .A3(new_n825), .A4(new_n298), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n817), .A2(new_n818), .A3(new_n692), .A4(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n736), .A2(new_n660), .A3(new_n826), .A4(new_n692), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT116), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n827), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n829), .A2(new_n828), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n834));
  INV_X1    g648(.A(new_n649), .ZN(new_n835));
  INV_X1    g649(.A(new_n636), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n355), .A2(new_n634), .A3(new_n363), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n836), .A2(new_n837), .B1(G475), .B2(new_n367), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n405), .A2(new_n655), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n556), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n604), .A2(KEYINPUT107), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n642), .A2(new_n720), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n841), .A2(new_n691), .A3(new_n735), .A4(new_n842), .ZN(new_n843));
  AOI211_X1 g657(.A(new_n835), .B(new_n739), .C1(new_n840), .C2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n630), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n407), .B1(new_n770), .B2(new_n628), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n846), .B1(new_n847), .B2(new_n845), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n607), .A3(new_n606), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n755), .A3(new_n601), .A4(new_n650), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n844), .A2(new_n850), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n710), .A2(new_n714), .A3(new_n730), .A4(new_n718), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n851), .A2(new_n852), .A3(new_n752), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n833), .A2(new_n834), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n851), .A2(new_n852), .A3(new_n752), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n829), .A2(KEYINPUT116), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n829), .A2(KEYINPUT116), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT52), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n855), .B1(new_n858), .B2(new_n831), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n854), .B(KEYINPUT54), .C1(new_n834), .C2(new_n859), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n856), .A2(new_n857), .A3(KEYINPUT52), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n828), .B1(new_n827), .B2(new_n830), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n853), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n834), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n865));
  INV_X1    g679(.A(new_n851), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n710), .A2(new_n714), .A3(new_n730), .A4(new_n718), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n747), .A2(new_n600), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n868), .A2(KEYINPUT42), .A3(new_n298), .A4(new_n750), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n867), .B1(new_n743), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT117), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n866), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n852), .A2(new_n752), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n834), .B1(new_n873), .B2(KEYINPUT117), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n872), .A2(new_n874), .A3(new_n833), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n864), .A2(new_n865), .A3(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n815), .A2(new_n816), .A3(new_n860), .A4(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n808), .A2(new_n709), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n868), .A2(new_n773), .A3(new_n806), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT48), .Z(new_n880));
  NOR3_X1   g694(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(G952), .A2(G953), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n797), .B1(new_n881), .B2(new_n882), .ZN(G75));
  NAND2_X1  g697(.A1(new_n864), .A2(new_n875), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(G902), .A3(new_n422), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT119), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n456), .A2(new_n458), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT118), .Z(new_n888));
  XOR2_X1   g702(.A(new_n439), .B(KEYINPUT55), .Z(new_n889));
  XNOR2_X1  g703(.A(new_n888), .B(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT56), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n886), .A2(new_n890), .B1(new_n891), .B2(new_n885), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n893));
  AND4_X1   g707(.A1(new_n893), .A2(new_n885), .A3(new_n891), .A4(new_n890), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n411), .A2(G952), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(G51));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n872), .A2(new_n833), .A3(new_n874), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n858), .A2(new_n831), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT53), .B1(new_n899), .B2(new_n853), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(new_n286), .ZN(new_n902));
  INV_X1    g716(.A(new_n762), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n897), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR4_X1   g718(.A1(new_n901), .A2(KEYINPUT121), .A3(new_n286), .A4(new_n762), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT54), .B1(new_n898), .B2(new_n900), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n907), .A2(new_n908), .A3(new_n876), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n901), .A2(KEYINPUT120), .A3(new_n865), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n763), .B(KEYINPUT57), .Z(new_n911));
  NAND3_X1  g725(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n285), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n895), .B1(new_n906), .B2(new_n913), .ZN(G54));
  NAND3_X1  g728(.A1(new_n902), .A2(KEYINPUT58), .A3(G475), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n915), .A2(new_n360), .A3(new_n352), .ZN(new_n916));
  INV_X1    g730(.A(new_n895), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n902), .A2(KEYINPUT58), .A3(G475), .A4(new_n361), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(G60));
  INV_X1    g733(.A(new_n622), .ZN(new_n920));
  NAND2_X1  g734(.A1(G478), .A2(G902), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT59), .Z(new_n922));
  NOR2_X1   g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n909), .A2(new_n910), .A3(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT122), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n876), .A2(new_n860), .ZN(new_n927));
  INV_X1    g741(.A(new_n922), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n895), .B1(new_n929), .B2(new_n920), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT122), .A4(new_n923), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n926), .A2(new_n930), .A3(new_n931), .ZN(G63));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n646), .A2(new_n647), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT60), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n935), .B(new_n938), .C1(new_n898), .C2(new_n900), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n917), .ZN(new_n940));
  AOI22_X1  g754(.A1(new_n884), .A2(new_n938), .B1(new_n597), .B2(new_n595), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n940), .A2(new_n941), .A3(KEYINPUT123), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n937), .B1(new_n864), .B2(new_n875), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n895), .B1(new_n944), .B2(new_n935), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n938), .B1(new_n898), .B2(new_n900), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n595), .A2(new_n597), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n943), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n933), .B1(new_n942), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(KEYINPUT123), .B1(new_n940), .B2(new_n941), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n945), .A2(new_n943), .A3(new_n948), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n951), .A2(new_n952), .A3(KEYINPUT61), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n950), .A2(new_n953), .ZN(G66));
  OAI21_X1  g768(.A(G953), .B1(new_n417), .B2(new_n423), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n849), .A2(new_n601), .A3(new_n650), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n852), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n955), .B1(new_n958), .B2(G953), .ZN(new_n959));
  INV_X1    g773(.A(new_n888), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(G898), .B2(new_n411), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n959), .B(new_n961), .ZN(G69));
  NAND2_X1  g776(.A1(new_n817), .A2(new_n692), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n963), .A2(KEYINPUT125), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(KEYINPUT125), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n964), .A2(new_n687), .A3(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n782), .A2(new_n788), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n697), .A2(new_n683), .A3(new_n848), .A4(new_n740), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n411), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n315), .A2(new_n318), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT124), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(G953), .B1(new_n262), .B2(new_n654), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(KEYINPUT126), .ZN(new_n979));
  OR2_X1    g793(.A1(new_n978), .A2(KEYINPUT126), .ZN(new_n980));
  NAND2_X1  g794(.A1(G900), .A2(G953), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n868), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n983), .A2(new_n769), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n825), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n782), .A2(new_n755), .A3(new_n788), .A4(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n964), .A2(new_n752), .A3(new_n965), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n982), .B1(new_n988), .B2(new_n411), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n977), .A2(new_n979), .A3(new_n980), .A4(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n976), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(new_n971), .B2(new_n411), .ZN(new_n993));
  OAI211_X1 g807(.A(KEYINPUT126), .B(new_n978), .C1(new_n993), .C2(new_n989), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n991), .A2(new_n994), .ZN(G72));
  OR2_X1    g809(.A1(new_n971), .A2(new_n957), .ZN(new_n996));
  NAND2_X1  g810(.A1(G472), .A2(G902), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT63), .Z(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT127), .Z(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n666), .B1(new_n996), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n999), .B1(new_n988), .B2(new_n958), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n1002), .A2(new_n519), .A3(new_n528), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n854), .B(new_n998), .C1(new_n834), .C2(new_n859), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n530), .A2(new_n543), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n917), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n1001), .A2(new_n1003), .A3(new_n1006), .ZN(G57));
endmodule


