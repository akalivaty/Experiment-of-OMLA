

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739;

  XNOR2_X1 U370 ( .A(n380), .B(n524), .ZN(n727) );
  INV_X1 U371 ( .A(G953), .ZN(n730) );
  XNOR2_X2 U372 ( .A(KEYINPUT91), .B(KEYINPUT18), .ZN(n402) );
  XNOR2_X2 U373 ( .A(G137), .B(KEYINPUT71), .ZN(n378) );
  XNOR2_X2 U374 ( .A(n557), .B(KEYINPUT33), .ZN(n663) );
  NOR2_X2 U375 ( .A1(n567), .A2(n556), .ZN(n557) );
  NOR2_X2 U376 ( .A1(n364), .A2(n624), .ZN(n488) );
  XNOR2_X2 U377 ( .A(n537), .B(n536), .ZN(n598) );
  XNOR2_X2 U378 ( .A(n513), .B(KEYINPUT22), .ZN(n552) );
  NAND2_X2 U379 ( .A1(n427), .A2(n512), .ZN(n513) );
  AND2_X1 U380 ( .A1(n467), .A2(n633), .ZN(n563) );
  XNOR2_X1 U381 ( .A(n607), .B(n357), .ZN(n608) );
  AND2_X1 U382 ( .A1(n391), .A2(n390), .ZN(n387) );
  NOR2_X1 U383 ( .A1(n432), .A2(n434), .ZN(n368) );
  INV_X1 U384 ( .A(n427), .ZN(n558) );
  NAND2_X1 U385 ( .A1(n608), .A2(n490), .ZN(n492) );
  XNOR2_X1 U386 ( .A(n428), .B(KEYINPUT38), .ZN(n682) );
  XNOR2_X1 U387 ( .A(n369), .B(n348), .ZN(n554) );
  NOR2_X1 U388 ( .A1(G902), .A2(n703), .ZN(n537) );
  XNOR2_X1 U389 ( .A(n379), .B(n522), .ZN(n626) );
  XNOR2_X1 U390 ( .A(n506), .B(n466), .ZN(n726) );
  XNOR2_X1 U391 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U392 ( .A(n399), .B(G125), .ZN(n506) );
  XNOR2_X1 U393 ( .A(n404), .B(G122), .ZN(n508) );
  XNOR2_X1 U394 ( .A(KEYINPUT83), .B(KEYINPUT17), .ZN(n401) );
  XNOR2_X1 U395 ( .A(n523), .B(n441), .ZN(n675) );
  INV_X1 U396 ( .A(G472), .ZN(n441) );
  NAND2_X1 U397 ( .A1(n367), .A2(n354), .ZN(n729) );
  XNOR2_X1 U398 ( .A(n368), .B(n363), .ZN(n367) );
  INV_X1 U399 ( .A(n655), .ZN(n366) );
  XNOR2_X1 U400 ( .A(n611), .B(n425), .ZN(n424) );
  INV_X1 U401 ( .A(KEYINPUT47), .ZN(n425) );
  XOR2_X1 U402 ( .A(KEYINPUT70), .B(G131), .Z(n514) );
  INV_X1 U403 ( .A(G146), .ZN(n399) );
  XNOR2_X1 U404 ( .A(n508), .B(n507), .ZN(n465) );
  XNOR2_X1 U405 ( .A(n475), .B(KEYINPUT76), .ZN(n525) );
  INV_X1 U406 ( .A(G107), .ZN(n475) );
  XNOR2_X1 U407 ( .A(n409), .B(n347), .ZN(n569) );
  OR2_X1 U408 ( .A1(n704), .A2(G902), .ZN(n409) );
  NAND2_X1 U409 ( .A1(n596), .A2(n594), .ZN(n669) );
  XNOR2_X1 U410 ( .A(n443), .B(n442), .ZN(n521) );
  XNOR2_X1 U411 ( .A(G116), .B(KEYINPUT3), .ZN(n442) );
  XNOR2_X1 U412 ( .A(n444), .B(G101), .ZN(n443) );
  XNOR2_X1 U413 ( .A(KEYINPUT74), .B(G113), .ZN(n444) );
  XNOR2_X1 U414 ( .A(n405), .B(G110), .ZN(n365) );
  INV_X1 U415 ( .A(G119), .ZN(n405) );
  NAND2_X1 U416 ( .A1(n388), .A2(n625), .ZN(n446) );
  NAND2_X1 U417 ( .A1(n413), .A2(n412), .ZN(n620) );
  NOR2_X1 U418 ( .A1(n729), .A2(n660), .ZN(n412) );
  INV_X1 U419 ( .A(n411), .ZN(n428) );
  XNOR2_X1 U420 ( .A(n371), .B(KEYINPUT28), .ZN(n599) );
  NOR2_X1 U421 ( .A1(n605), .A2(n597), .ZN(n371) );
  NAND2_X1 U422 ( .A1(n373), .A2(n372), .ZN(n433) );
  XNOR2_X1 U423 ( .A(n456), .B(KEYINPUT87), .ZN(n455) );
  INV_X1 U424 ( .A(KEYINPUT68), .ZN(n383) );
  XNOR2_X1 U425 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n498) );
  XNOR2_X1 U426 ( .A(G143), .B(KEYINPUT11), .ZN(n462) );
  XNOR2_X1 U427 ( .A(n514), .B(n355), .ZN(n463) );
  INV_X1 U428 ( .A(G104), .ZN(n404) );
  XNOR2_X1 U429 ( .A(G128), .B(G137), .ZN(n539) );
  XNOR2_X1 U430 ( .A(n419), .B(n544), .ZN(n414) );
  XNOR2_X1 U431 ( .A(n365), .B(n420), .ZN(n419) );
  INV_X1 U432 ( .A(KEYINPUT23), .ZN(n420) );
  XNOR2_X1 U433 ( .A(G140), .B(KEYINPUT10), .ZN(n466) );
  XNOR2_X1 U434 ( .A(KEYINPUT85), .B(n658), .ZN(n662) );
  NOR2_X1 U435 ( .A1(n686), .A2(n684), .ZN(n600) );
  XNOR2_X1 U436 ( .A(n437), .B(n436), .ZN(n602) );
  INV_X1 U437 ( .A(KEYINPUT39), .ZN(n436) );
  NAND2_X1 U438 ( .A1(n411), .A2(n681), .ZN(n607) );
  AND2_X1 U439 ( .A1(n606), .A2(n458), .ZN(n457) );
  INV_X1 U440 ( .A(n605), .ZN(n458) );
  NAND2_X1 U441 ( .A1(n454), .A2(n559), .ZN(n453) );
  NAND2_X1 U442 ( .A1(n558), .A2(KEYINPUT34), .ZN(n451) );
  INV_X1 U443 ( .A(n558), .ZN(n454) );
  OR2_X1 U444 ( .A1(n710), .A2(G902), .ZN(n369) );
  INV_X1 U445 ( .A(KEYINPUT25), .ZN(n547) );
  XNOR2_X1 U446 ( .A(n570), .B(n459), .ZN(n604) );
  INV_X1 U447 ( .A(KEYINPUT102), .ZN(n459) );
  NOR2_X1 U448 ( .A1(n564), .A2(n669), .ZN(n593) );
  XNOR2_X1 U449 ( .A(n520), .B(n521), .ZN(n522) );
  XNOR2_X1 U450 ( .A(n727), .B(n533), .ZN(n703) );
  XNOR2_X1 U451 ( .A(G101), .B(G140), .ZN(n532) );
  AND2_X1 U452 ( .A1(n446), .A2(G469), .ZN(n393) );
  NAND2_X1 U453 ( .A1(n659), .A2(n438), .ZN(n439) );
  AND2_X1 U454 ( .A1(n446), .A2(G210), .ZN(n438) );
  XNOR2_X1 U455 ( .A(n400), .B(G128), .ZN(n493) );
  NOR2_X1 U456 ( .A1(G953), .A2(G237), .ZN(n518) );
  XNOR2_X1 U457 ( .A(n493), .B(n449), .ZN(n515) );
  INV_X1 U458 ( .A(G134), .ZN(n449) );
  XNOR2_X1 U459 ( .A(n525), .B(n474), .ZN(n479) );
  XNOR2_X1 U460 ( .A(KEYINPUT82), .B(KEYINPUT92), .ZN(n474) );
  NAND2_X1 U461 ( .A1(G234), .A2(G237), .ZN(n483) );
  OR2_X1 U462 ( .A1(n455), .A2(n435), .ZN(n434) );
  XNOR2_X1 U463 ( .A(n433), .B(KEYINPUT46), .ZN(n432) );
  INV_X1 U464 ( .A(KEYINPUT48), .ZN(n614) );
  NAND2_X1 U465 ( .A1(n554), .A2(n418), .ZN(n605) );
  NOR2_X1 U466 ( .A1(n664), .A2(n595), .ZN(n418) );
  XNOR2_X1 U467 ( .A(n598), .B(n538), .ZN(n668) );
  INV_X1 U468 ( .A(KEYINPUT1), .ZN(n538) );
  XNOR2_X1 U469 ( .A(G146), .B(G119), .ZN(n516) );
  XOR2_X1 U470 ( .A(KEYINPUT97), .B(KEYINPUT5), .Z(n517) );
  XNOR2_X1 U471 ( .A(n408), .B(n515), .ZN(n380) );
  XNOR2_X1 U472 ( .A(n448), .B(n514), .ZN(n408) );
  XNOR2_X1 U473 ( .A(n378), .B(KEYINPUT4), .ZN(n448) );
  XNOR2_X1 U474 ( .A(G116), .B(G107), .ZN(n494) );
  XOR2_X1 U475 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n495) );
  XNOR2_X1 U476 ( .A(n463), .B(n461), .ZN(n460) );
  XNOR2_X1 U477 ( .A(n726), .B(n465), .ZN(n464) );
  XNOR2_X1 U478 ( .A(n462), .B(G113), .ZN(n461) );
  XNOR2_X1 U479 ( .A(G146), .B(G104), .ZN(n526) );
  XNOR2_X1 U480 ( .A(n528), .B(n527), .ZN(n529) );
  INV_X1 U481 ( .A(G110), .ZN(n527) );
  AND2_X1 U482 ( .A1(n592), .A2(n593), .ZN(n612) );
  XNOR2_X1 U483 ( .A(n440), .B(KEYINPUT30), .ZN(n591) );
  NAND2_X1 U484 ( .A1(n675), .A2(n681), .ZN(n440) );
  XNOR2_X1 U485 ( .A(n569), .B(KEYINPUT99), .ZN(n571) );
  XNOR2_X1 U486 ( .A(n377), .B(n521), .ZN(n715) );
  XOR2_X1 U487 ( .A(KEYINPUT77), .B(KEYINPUT16), .Z(n478) );
  XNOR2_X1 U488 ( .A(n370), .B(n545), .ZN(n710) );
  XNOR2_X1 U489 ( .A(n414), .B(n543), .ZN(n370) );
  AND2_X1 U490 ( .A1(n659), .A2(n446), .ZN(n395) );
  AND2_X1 U491 ( .A1(n446), .A2(G475), .ZN(n445) );
  NAND2_X1 U492 ( .A1(n661), .A2(n431), .ZN(n430) );
  NOR2_X1 U493 ( .A1(n662), .A2(n353), .ZN(n431) );
  NAND2_X1 U494 ( .A1(n619), .A2(n428), .ZN(n656) );
  XNOR2_X1 U495 ( .A(n601), .B(n374), .ZN(n373) );
  INV_X1 U496 ( .A(KEYINPUT42), .ZN(n374) );
  NOR2_X1 U497 ( .A1(n602), .A2(n604), .ZN(n603) );
  NAND2_X1 U498 ( .A1(n417), .A2(n616), .ZN(n456) );
  XNOR2_X1 U499 ( .A(n410), .B(KEYINPUT36), .ZN(n417) );
  NOR2_X1 U500 ( .A1(n615), .A2(n607), .ZN(n410) );
  INV_X1 U501 ( .A(KEYINPUT35), .ZN(n560) );
  NOR2_X1 U502 ( .A1(n663), .A2(n453), .ZN(n452) );
  XNOR2_X1 U503 ( .A(n568), .B(KEYINPUT31), .ZN(n407) );
  NOR2_X1 U504 ( .A1(n610), .A2(n609), .ZN(n641) );
  INV_X1 U505 ( .A(n593), .ZN(n426) );
  NAND2_X1 U506 ( .A1(n472), .A2(n390), .ZN(n471) );
  XNOR2_X1 U507 ( .A(n473), .B(n359), .ZN(n472) );
  NAND2_X1 U508 ( .A1(n469), .A2(n390), .ZN(n468) );
  XNOR2_X1 U509 ( .A(n470), .B(n360), .ZN(n469) );
  INV_X1 U510 ( .A(KEYINPUT56), .ZN(n385) );
  NAND2_X1 U511 ( .A1(n389), .A2(n390), .ZN(n386) );
  XNOR2_X1 U512 ( .A(n439), .B(n362), .ZN(n389) );
  XNOR2_X1 U513 ( .A(n382), .B(n381), .ZN(G75) );
  INV_X1 U514 ( .A(KEYINPUT53), .ZN(n381) );
  NAND2_X1 U515 ( .A1(n430), .A2(n429), .ZN(n382) );
  AND2_X1 U516 ( .A1(n701), .A2(n730), .ZN(n429) );
  XOR2_X1 U517 ( .A(KEYINPUT13), .B(G475), .Z(n347) );
  XOR2_X1 U518 ( .A(n548), .B(n547), .Z(n348) );
  AND2_X1 U519 ( .A1(G224), .A2(n730), .ZN(n349) );
  NAND2_X1 U520 ( .A1(G210), .A2(n489), .ZN(n350) );
  AND2_X1 U521 ( .A1(n572), .A2(n569), .ZN(n351) );
  AND2_X1 U522 ( .A1(n451), .A2(n351), .ZN(n352) );
  AND2_X1 U523 ( .A1(n729), .A2(n660), .ZN(n353) );
  INV_X1 U524 ( .A(n554), .ZN(n594) );
  AND2_X1 U525 ( .A1(n656), .A2(n366), .ZN(n354) );
  AND2_X1 U526 ( .A1(G214), .A2(n518), .ZN(n355) );
  AND2_X1 U527 ( .A1(n351), .A2(n411), .ZN(n356) );
  BUF_X1 U528 ( .A(n668), .Z(n423) );
  XNOR2_X1 U529 ( .A(KEYINPUT19), .B(KEYINPUT66), .ZN(n357) );
  XNOR2_X1 U530 ( .A(n491), .B(KEYINPUT90), .ZN(n358) );
  XNOR2_X1 U531 ( .A(n604), .B(KEYINPUT106), .ZN(n645) );
  XOR2_X1 U532 ( .A(n626), .B(KEYINPUT62), .Z(n359) );
  XOR2_X1 U533 ( .A(n703), .B(n702), .Z(n360) );
  XNOR2_X1 U534 ( .A(n704), .B(n476), .ZN(n361) );
  XOR2_X1 U535 ( .A(n482), .B(n481), .Z(n362) );
  XOR2_X1 U536 ( .A(n614), .B(KEYINPUT72), .Z(n363) );
  NOR2_X1 U537 ( .A1(G952), .A2(n730), .ZN(n714) );
  INV_X1 U538 ( .A(n714), .ZN(n390) );
  XNOR2_X1 U539 ( .A(n364), .B(KEYINPUT84), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n375), .B(n715), .ZN(n364) );
  XNOR2_X1 U541 ( .A(n563), .B(KEYINPUT89), .ZN(n580) );
  XNOR2_X1 U542 ( .A(n365), .B(n508), .ZN(n403) );
  INV_X1 U543 ( .A(n739), .ZN(n372) );
  XNOR2_X1 U544 ( .A(n373), .B(G137), .ZN(G39) );
  XNOR2_X1 U545 ( .A(n376), .B(n480), .ZN(n375) );
  XNOR2_X1 U546 ( .A(n396), .B(n398), .ZN(n376) );
  XNOR2_X1 U547 ( .A(n403), .B(n478), .ZN(n377) );
  INV_X1 U548 ( .A(n380), .ZN(n379) );
  XNOR2_X1 U549 ( .A(n384), .B(n383), .ZN(n581) );
  NOR2_X1 U550 ( .A1(n737), .A2(KEYINPUT44), .ZN(n384) );
  XNOR2_X1 U551 ( .A(n386), .B(n385), .ZN(G51) );
  XNOR2_X1 U552 ( .A(n387), .B(n705), .ZN(G60) );
  NOR2_X1 U553 ( .A1(n668), .A2(n669), .ZN(n555) );
  NAND2_X1 U554 ( .A1(n623), .A2(n624), .ZN(n388) );
  XNOR2_X1 U555 ( .A(n447), .B(n361), .ZN(n391) );
  NAND2_X1 U556 ( .A1(n392), .A2(n685), .ZN(n575) );
  NAND2_X1 U557 ( .A1(n406), .A2(n629), .ZN(n392) );
  NOR2_X1 U558 ( .A1(n680), .A2(n610), .ZN(n421) );
  AND2_X1 U559 ( .A1(n446), .A2(G472), .ZN(n394) );
  NAND2_X1 U560 ( .A1(n659), .A2(n393), .ZN(n470) );
  NAND2_X1 U561 ( .A1(n659), .A2(n394), .ZN(n473) );
  NAND2_X1 U562 ( .A1(n395), .A2(G478), .ZN(n707) );
  NAND2_X1 U563 ( .A1(n395), .A2(G217), .ZN(n711) );
  XNOR2_X1 U564 ( .A(n397), .B(n493), .ZN(n396) );
  XNOR2_X1 U565 ( .A(n401), .B(n402), .ZN(n397) );
  XNOR2_X1 U566 ( .A(n349), .B(n506), .ZN(n398) );
  INV_X1 U567 ( .A(G143), .ZN(n400) );
  INV_X1 U568 ( .A(n407), .ZN(n406) );
  AND2_X1 U569 ( .A1(n407), .A2(n642), .ZN(n647) );
  AND2_X1 U570 ( .A1(n407), .A2(n634), .ZN(n651) );
  NOR2_X1 U571 ( .A1(n571), .A2(n572), .ZN(n570) );
  NAND2_X1 U572 ( .A1(n642), .A2(n457), .ZN(n615) );
  XNOR2_X2 U573 ( .A(n488), .B(n350), .ZN(n411) );
  NOR2_X1 U574 ( .A1(n657), .A2(n729), .ZN(n623) );
  INV_X1 U575 ( .A(n657), .ZN(n413) );
  NAND2_X1 U576 ( .A1(n415), .A2(n554), .ZN(n633) );
  XNOR2_X1 U577 ( .A(n553), .B(KEYINPUT64), .ZN(n415) );
  NAND2_X1 U578 ( .A1(n416), .A2(KEYINPUT44), .ZN(n578) );
  NAND2_X1 U579 ( .A1(n563), .A2(n562), .ZN(n416) );
  XNOR2_X1 U580 ( .A(n464), .B(n460), .ZN(n704) );
  XNOR2_X1 U581 ( .A(n421), .B(KEYINPUT108), .ZN(n601) );
  NOR2_X1 U582 ( .A1(n422), .A2(n452), .ZN(n561) );
  NAND2_X1 U583 ( .A1(n450), .A2(n352), .ZN(n422) );
  NAND2_X1 U584 ( .A1(n424), .A2(n640), .ZN(n613) );
  XNOR2_X2 U585 ( .A(n492), .B(n358), .ZN(n427) );
  NOR2_X1 U586 ( .A1(n558), .A2(n426), .ZN(n565) );
  NAND2_X1 U587 ( .A1(n677), .A2(n454), .ZN(n568) );
  XNOR2_X1 U588 ( .A(n613), .B(KEYINPUT78), .ZN(n435) );
  NAND2_X1 U589 ( .A1(n612), .A2(n682), .ZN(n437) );
  XNOR2_X2 U590 ( .A(n620), .B(KEYINPUT80), .ZN(n659) );
  INV_X1 U591 ( .A(n675), .ZN(n597) );
  NAND2_X1 U592 ( .A1(n445), .A2(n659), .ZN(n447) );
  NAND2_X1 U593 ( .A1(n663), .A2(KEYINPUT34), .ZN(n450) );
  INV_X1 U594 ( .A(n456), .ZN(n652) );
  XNOR2_X1 U595 ( .A(n467), .B(G119), .ZN(G21) );
  XNOR2_X2 U596 ( .A(n550), .B(KEYINPUT32), .ZN(n467) );
  XNOR2_X1 U597 ( .A(n468), .B(KEYINPUT121), .ZN(G54) );
  XNOR2_X1 U598 ( .A(n471), .B(KEYINPUT63), .ZN(G57) );
  INV_X1 U599 ( .A(n645), .ZN(n642) );
  XNOR2_X2 U600 ( .A(n584), .B(KEYINPUT45), .ZN(n657) );
  NOR2_X2 U601 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U602 ( .A(KEYINPUT59), .B(KEYINPUT65), .Z(n476) );
  AND2_X1 U603 ( .A1(n518), .A2(G210), .ZN(n477) );
  XNOR2_X1 U604 ( .A(n519), .B(n477), .ZN(n520) );
  XNOR2_X1 U605 ( .A(n530), .B(n529), .ZN(n531) );
  BUF_X1 U606 ( .A(n737), .Z(n738) );
  XOR2_X1 U607 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n482) );
  XNOR2_X1 U608 ( .A(KEYINPUT4), .B(n479), .ZN(n480) );
  XNOR2_X1 U609 ( .A(n483), .B(KEYINPUT14), .ZN(n485) );
  NAND2_X1 U610 ( .A1(G952), .A2(n485), .ZN(n697) );
  NOR2_X1 U611 ( .A1(G953), .A2(n697), .ZN(n484) );
  XNOR2_X1 U612 ( .A(KEYINPUT93), .B(n484), .ZN(n585) );
  NAND2_X1 U613 ( .A1(G902), .A2(n485), .ZN(n586) );
  INV_X1 U614 ( .A(n586), .ZN(n486) );
  NOR2_X1 U615 ( .A1(G898), .A2(n730), .ZN(n717) );
  NAND2_X1 U616 ( .A1(n486), .A2(n717), .ZN(n487) );
  NAND2_X1 U617 ( .A1(n585), .A2(n487), .ZN(n490) );
  XNOR2_X1 U618 ( .A(G902), .B(KEYINPUT15), .ZN(n621) );
  INV_X1 U619 ( .A(n621), .ZN(n624) );
  OR2_X1 U620 ( .A1(G237), .A2(G902), .ZN(n489) );
  NAND2_X1 U621 ( .A1(G214), .A2(n489), .ZN(n681) );
  XNOR2_X1 U622 ( .A(KEYINPUT0), .B(KEYINPUT67), .ZN(n491) );
  XNOR2_X1 U623 ( .A(KEYINPUT101), .B(G478), .ZN(n505) );
  INV_X1 U624 ( .A(n515), .ZN(n497) );
  XNOR2_X1 U625 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U626 ( .A(n497), .B(n496), .Z(n503) );
  XOR2_X1 U627 ( .A(G122), .B(KEYINPUT100), .Z(n501) );
  NAND2_X1 U628 ( .A1(n730), .A2(G234), .ZN(n499) );
  XNOR2_X1 U629 ( .A(n498), .B(n499), .ZN(n542) );
  NAND2_X1 U630 ( .A1(G217), .A2(n542), .ZN(n500) );
  XNOR2_X1 U631 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U632 ( .A(n503), .B(n502), .ZN(n706) );
  NOR2_X1 U633 ( .A1(G902), .A2(n706), .ZN(n504) );
  XNOR2_X1 U634 ( .A(n505), .B(n504), .ZN(n572) );
  XOR2_X1 U635 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n507) );
  NOR2_X1 U636 ( .A1(n572), .A2(n569), .ZN(n509) );
  XNOR2_X1 U637 ( .A(KEYINPUT103), .B(n509), .ZN(n684) );
  NAND2_X1 U638 ( .A1(G234), .A2(n621), .ZN(n510) );
  XNOR2_X1 U639 ( .A(KEYINPUT20), .B(n510), .ZN(n546) );
  NAND2_X1 U640 ( .A1(n546), .A2(G221), .ZN(n511) );
  XNOR2_X1 U641 ( .A(KEYINPUT21), .B(n511), .ZN(n664) );
  NOR2_X1 U642 ( .A1(n684), .A2(n664), .ZN(n512) );
  XNOR2_X1 U643 ( .A(n517), .B(n516), .ZN(n519) );
  NOR2_X1 U644 ( .A1(n626), .A2(G902), .ZN(n523) );
  XOR2_X1 U645 ( .A(KEYINPUT6), .B(n675), .Z(n606) );
  NOR2_X2 U646 ( .A1(n552), .A2(n606), .ZN(n574) );
  INV_X1 U647 ( .A(KEYINPUT94), .ZN(n524) );
  XNOR2_X1 U648 ( .A(n526), .B(n525), .ZN(n530) );
  NAND2_X1 U649 ( .A1(G227), .A2(n730), .ZN(n528) );
  XNOR2_X1 U650 ( .A(n532), .B(n531), .ZN(n533) );
  INV_X1 U651 ( .A(G469), .ZN(n535) );
  INV_X1 U652 ( .A(KEYINPUT73), .ZN(n534) );
  INV_X1 U653 ( .A(n423), .ZN(n616) );
  XOR2_X1 U654 ( .A(KEYINPUT75), .B(KEYINPUT24), .Z(n540) );
  XNOR2_X1 U655 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U656 ( .A(n541), .B(n726), .ZN(n545) );
  NAND2_X1 U657 ( .A1(G221), .A2(n542), .ZN(n543) );
  XOR2_X1 U658 ( .A(KEYINPUT81), .B(KEYINPUT95), .Z(n544) );
  NAND2_X1 U659 ( .A1(G217), .A2(n546), .ZN(n548) );
  XNOR2_X1 U660 ( .A(KEYINPUT104), .B(n554), .ZN(n665) );
  AND2_X1 U661 ( .A1(n616), .A2(n665), .ZN(n549) );
  NAND2_X1 U662 ( .A1(n574), .A2(n549), .ZN(n550) );
  NAND2_X1 U663 ( .A1(n423), .A2(n597), .ZN(n551) );
  NOR2_X1 U664 ( .A1(n552), .A2(n551), .ZN(n553) );
  INV_X1 U665 ( .A(KEYINPUT34), .ZN(n559) );
  INV_X1 U666 ( .A(n664), .ZN(n596) );
  XNOR2_X1 U667 ( .A(n555), .B(KEYINPUT79), .ZN(n567) );
  INV_X1 U668 ( .A(n606), .ZN(n556) );
  XNOR2_X1 U669 ( .A(n561), .B(n560), .ZN(n737) );
  INV_X1 U670 ( .A(n737), .ZN(n562) );
  INV_X1 U671 ( .A(n598), .ZN(n564) );
  XNOR2_X1 U672 ( .A(n565), .B(KEYINPUT96), .ZN(n566) );
  NAND2_X1 U673 ( .A1(n566), .A2(n597), .ZN(n629) );
  NOR2_X1 U674 ( .A1(n597), .A2(n567), .ZN(n677) );
  NAND2_X1 U675 ( .A1(n572), .A2(n571), .ZN(n649) );
  NAND2_X1 U676 ( .A1(n604), .A2(n649), .ZN(n685) );
  NOR2_X1 U677 ( .A1(n616), .A2(n665), .ZN(n573) );
  NAND2_X1 U678 ( .A1(n574), .A2(n573), .ZN(n627) );
  NAND2_X1 U679 ( .A1(n575), .A2(n627), .ZN(n576) );
  XNOR2_X1 U680 ( .A(KEYINPUT105), .B(n576), .ZN(n577) );
  NAND2_X1 U681 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U682 ( .A(n579), .B(KEYINPUT88), .ZN(n583) );
  NOR2_X1 U683 ( .A1(n581), .A2(n580), .ZN(n582) );
  INV_X1 U684 ( .A(n585), .ZN(n590) );
  NOR2_X1 U685 ( .A1(G900), .A2(n586), .ZN(n587) );
  NAND2_X1 U686 ( .A1(G953), .A2(n587), .ZN(n588) );
  XNOR2_X1 U687 ( .A(KEYINPUT107), .B(n588), .ZN(n589) );
  NOR2_X1 U688 ( .A1(n590), .A2(n589), .ZN(n595) );
  NOR2_X1 U689 ( .A1(n595), .A2(n591), .ZN(n592) );
  NOR2_X1 U690 ( .A1(n649), .A2(n602), .ZN(n655) );
  NAND2_X1 U691 ( .A1(n599), .A2(n598), .ZN(n610) );
  NAND2_X1 U692 ( .A1(n682), .A2(n681), .ZN(n686) );
  XNOR2_X1 U693 ( .A(n600), .B(KEYINPUT41), .ZN(n680) );
  XNOR2_X1 U694 ( .A(KEYINPUT40), .B(n603), .ZN(n739) );
  INV_X1 U695 ( .A(n608), .ZN(n609) );
  NAND2_X1 U696 ( .A1(n641), .A2(n685), .ZN(n611) );
  NAND2_X1 U697 ( .A1(n612), .A2(n356), .ZN(n640) );
  NOR2_X1 U698 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U699 ( .A1(n617), .A2(n681), .ZN(n618) );
  XNOR2_X1 U700 ( .A(KEYINPUT43), .B(n618), .ZN(n619) );
  XOR2_X1 U701 ( .A(n621), .B(KEYINPUT86), .Z(n622) );
  NAND2_X1 U702 ( .A1(n622), .A2(KEYINPUT2), .ZN(n625) );
  XNOR2_X1 U703 ( .A(G101), .B(n627), .ZN(G3) );
  NOR2_X1 U704 ( .A1(n645), .A2(n629), .ZN(n628) );
  XOR2_X1 U705 ( .A(G104), .B(n628), .Z(G6) );
  NOR2_X1 U706 ( .A1(n649), .A2(n629), .ZN(n631) );
  XNOR2_X1 U707 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n630) );
  XNOR2_X1 U708 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U709 ( .A(G107), .B(n632), .ZN(G9) );
  XNOR2_X1 U710 ( .A(n633), .B(G110), .ZN(G12) );
  XNOR2_X1 U711 ( .A(G128), .B(KEYINPUT110), .ZN(n638) );
  XOR2_X1 U712 ( .A(KEYINPUT29), .B(KEYINPUT111), .Z(n636) );
  INV_X1 U713 ( .A(n649), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n641), .A2(n634), .ZN(n635) );
  XNOR2_X1 U715 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U716 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U717 ( .A(KEYINPUT109), .B(n639), .ZN(G30) );
  XNOR2_X1 U718 ( .A(G143), .B(n640), .ZN(G45) );
  NAND2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U720 ( .A(n643), .B(KEYINPUT112), .ZN(n644) );
  XNOR2_X1 U721 ( .A(G146), .B(n644), .ZN(G48) );
  XNOR2_X1 U722 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n646) );
  XNOR2_X1 U723 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U724 ( .A(G113), .B(n648), .ZN(G15) );
  XNOR2_X1 U725 ( .A(G116), .B(KEYINPUT115), .ZN(n650) );
  XNOR2_X1 U726 ( .A(n651), .B(n650), .ZN(G18) );
  XNOR2_X1 U727 ( .A(n652), .B(KEYINPUT116), .ZN(n653) );
  XNOR2_X1 U728 ( .A(n653), .B(KEYINPUT37), .ZN(n654) );
  XNOR2_X1 U729 ( .A(G125), .B(n654), .ZN(G27) );
  XOR2_X1 U730 ( .A(G134), .B(n655), .Z(G36) );
  XNOR2_X1 U731 ( .A(G140), .B(n656), .ZN(G42) );
  INV_X1 U732 ( .A(KEYINPUT2), .ZN(n660) );
  NAND2_X1 U733 ( .A1(n657), .A2(n660), .ZN(n658) );
  BUF_X1 U734 ( .A(n659), .Z(n661) );
  BUF_X1 U735 ( .A(n663), .Z(n690) );
  NOR2_X1 U736 ( .A1(n680), .A2(n690), .ZN(n700) );
  NAND2_X1 U737 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U738 ( .A(n666), .B(KEYINPUT49), .ZN(n667) );
  XNOR2_X1 U739 ( .A(KEYINPUT117), .B(n667), .ZN(n673) );
  NAND2_X1 U740 ( .A1(n669), .A2(n423), .ZN(n670) );
  XNOR2_X1 U741 ( .A(n670), .B(KEYINPUT118), .ZN(n671) );
  XNOR2_X1 U742 ( .A(KEYINPUT50), .B(n671), .ZN(n672) );
  NAND2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U746 ( .A(KEYINPUT51), .B(n678), .Z(n679) );
  NOR2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n694) );
  NOR2_X1 U748 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n689) );
  INV_X1 U750 ( .A(n685), .ZN(n687) );
  NOR2_X1 U751 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U752 ( .A1(n689), .A2(n688), .ZN(n691) );
  NOR2_X1 U753 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U754 ( .A(KEYINPUT119), .B(n692), .Z(n693) );
  NOR2_X1 U755 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U756 ( .A(KEYINPUT120), .B(n695), .Z(n696) );
  XOR2_X1 U757 ( .A(KEYINPUT52), .B(n696), .Z(n698) );
  NOR2_X1 U758 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U759 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U760 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n702) );
  XNOR2_X1 U761 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n705) );
  XOR2_X1 U762 ( .A(n706), .B(KEYINPUT123), .Z(n708) );
  XNOR2_X1 U763 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U764 ( .A1(n714), .A2(n709), .ZN(G63) );
  XNOR2_X1 U765 ( .A(n710), .B(KEYINPUT124), .ZN(n712) );
  XNOR2_X1 U766 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U767 ( .A1(n714), .A2(n713), .ZN(G66) );
  XNOR2_X1 U768 ( .A(G107), .B(KEYINPUT126), .ZN(n716) );
  XNOR2_X1 U769 ( .A(n716), .B(n715), .ZN(n718) );
  NOR2_X1 U770 ( .A1(n718), .A2(n717), .ZN(n725) );
  XOR2_X1 U771 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n720) );
  NAND2_X1 U772 ( .A1(G224), .A2(G953), .ZN(n719) );
  XNOR2_X1 U773 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U774 ( .A1(n721), .A2(G898), .ZN(n723) );
  OR2_X1 U775 ( .A1(n657), .A2(G953), .ZN(n722) );
  NAND2_X1 U776 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U777 ( .A(n725), .B(n724), .ZN(G69) );
  XOR2_X1 U778 ( .A(n727), .B(n726), .Z(n732) );
  XOR2_X1 U779 ( .A(KEYINPUT127), .B(n732), .Z(n728) );
  XNOR2_X1 U780 ( .A(n729), .B(n728), .ZN(n731) );
  NAND2_X1 U781 ( .A1(n731), .A2(n730), .ZN(n736) );
  XNOR2_X1 U782 ( .A(G227), .B(n732), .ZN(n733) );
  NAND2_X1 U783 ( .A1(n733), .A2(G900), .ZN(n734) );
  NAND2_X1 U784 ( .A1(n734), .A2(G953), .ZN(n735) );
  NAND2_X1 U785 ( .A1(n736), .A2(n735), .ZN(G72) );
  XOR2_X1 U786 ( .A(n738), .B(G122), .Z(G24) );
  XOR2_X1 U787 ( .A(G131), .B(n739), .Z(G33) );
endmodule

