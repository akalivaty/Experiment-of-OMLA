//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n202));
  AOI22_X1  g001(.A1(new_n202), .A2(KEYINPUT88), .B1(G43gat), .B2(G50gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT88), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT15), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  OR2_X1    g005(.A1(KEYINPUT89), .A2(G50gat), .ZN(new_n207));
  INV_X1    g006(.A(G43gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(KEYINPUT89), .A2(G50gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT15), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT14), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(G29gat), .B2(G36gat), .ZN(new_n216));
  OR3_X1    g015(.A1(new_n215), .A2(G29gat), .A3(G36gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(G29gat), .A2(G36gat), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n214), .A2(new_n216), .A3(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n217), .A2(new_n216), .A3(new_n218), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(new_n213), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G15gat), .B(G22gat), .ZN(new_n224));
  INV_X1    g023(.A(G1gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT16), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(G1gat), .B2(new_n224), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(G8gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n223), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n229), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n220), .A2(new_n222), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n235), .B(KEYINPUT13), .Z(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT90), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n220), .A2(new_n238), .A3(KEYINPUT17), .A4(new_n222), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n206), .A2(new_n210), .B1(KEYINPUT15), .B2(new_n212), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n238), .B(new_n222), .C1(new_n240), .C2(new_n221), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT17), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n229), .B1(new_n239), .B2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n231), .A2(new_n232), .ZN(new_n245));
  INV_X1    g044(.A(new_n235), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n237), .B1(new_n247), .B2(KEYINPUT18), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n239), .A2(new_n243), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n231), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(new_n235), .A3(new_n230), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT18), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G113gat), .B(G141gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(G197gat), .ZN(new_n255));
  XOR2_X1   g054(.A(KEYINPUT11), .B(G169gat), .Z(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT12), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NOR3_X1   g058(.A1(new_n248), .A2(new_n253), .A3(new_n259), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n251), .A2(new_n252), .B1(new_n234), .B2(new_n236), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n247), .A2(KEYINPUT18), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n258), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n265));
  INV_X1    g064(.A(G120gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G113gat), .ZN(new_n267));
  INV_X1    g066(.A(G113gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G120gat), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT1), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G127gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G134gat), .ZN(new_n272));
  INV_X1    g071(.A(G134gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(G127gat), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT69), .B1(new_n271), .B2(G134gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n272), .A2(new_n274), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n277), .B1(new_n278), .B2(KEYINPUT69), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n276), .B1(new_n279), .B2(new_n270), .ZN(new_n280));
  AND2_X1   g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G141gat), .B(G148gat), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n283), .B1(new_n284), .B2(KEYINPUT2), .ZN(new_n285));
  INV_X1    g084(.A(G148gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(G141gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT74), .B(G148gat), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(G141gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT2), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n281), .B1(new_n290), .B2(new_n282), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n285), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT75), .B1(new_n280), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n286), .A2(KEYINPUT74), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT74), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G148gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n296), .A3(G141gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n287), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n290), .ZN(new_n300));
  INV_X1    g099(.A(G155gat), .ZN(new_n301));
  INV_X1    g100(.A(G162gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G141gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n304), .A2(G148gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n290), .B1(new_n287), .B2(new_n305), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n299), .A2(new_n303), .B1(new_n306), .B2(new_n283), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT69), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n309), .B1(new_n272), .B2(new_n274), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n267), .A2(new_n269), .ZN(new_n311));
  OAI22_X1  g110(.A1(new_n277), .A2(new_n310), .B1(new_n311), .B2(KEYINPUT1), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n307), .A2(new_n308), .A3(new_n312), .A4(new_n276), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n293), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT76), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT4), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT3), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n307), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n292), .A2(KEYINPUT3), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(new_n320), .A3(new_n280), .ZN(new_n321));
  NAND2_X1  g120(.A1(G225gat), .A2(G233gat), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT4), .B1(new_n293), .B2(new_n313), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n280), .A2(new_n292), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT76), .B1(new_n325), .B2(new_n316), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n317), .B(new_n323), .C1(new_n324), .C2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT77), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n280), .A2(new_n292), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n293), .A2(new_n313), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n322), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n328), .B1(new_n332), .B2(KEYINPUT5), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT5), .ZN(new_n334));
  AOI211_X1 g133(.A(KEYINPUT77), .B(new_n334), .C1(new_n330), .C2(new_n331), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n327), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G1gat), .B(G29gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(KEYINPUT0), .ZN(new_n338));
  XNOR2_X1  g137(.A(G57gat), .B(G85gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n321), .ZN(new_n341));
  NOR3_X1   g140(.A1(new_n341), .A2(KEYINPUT5), .A3(new_n331), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n325), .A2(KEYINPUT4), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n343), .B1(KEYINPUT4), .B2(new_n314), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n340), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n336), .A2(KEYINPUT78), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n340), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n342), .A2(new_n344), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n347), .B1(new_n336), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n265), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT78), .B1(new_n336), .B2(new_n345), .ZN(new_n351));
  INV_X1    g150(.A(new_n265), .ZN(new_n352));
  INV_X1    g151(.A(new_n348), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n332), .A2(KEYINPUT5), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT77), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n332), .A2(new_n328), .A3(KEYINPUT5), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n353), .B1(new_n357), .B2(new_n327), .ZN(new_n358));
  OAI22_X1  g157(.A1(new_n351), .A2(new_n352), .B1(new_n358), .B2(new_n347), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n350), .A2(new_n359), .ZN(new_n360));
  AND2_X1   g159(.A1(G211gat), .A2(G218gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(G211gat), .A2(G218gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(G197gat), .A2(G204gat), .ZN(new_n364));
  AND2_X1   g163(.A1(G197gat), .A2(G204gat), .ZN(new_n365));
  OAI22_X1  g164(.A1(new_n364), .A2(new_n365), .B1(new_n361), .B2(KEYINPUT22), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n363), .B1(new_n367), .B2(KEYINPUT70), .ZN(new_n368));
  INV_X1    g167(.A(new_n363), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT70), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT25), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT24), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n374), .A2(G183gat), .A3(G190gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(G183gat), .B(G190gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(new_n374), .ZN(new_n377));
  INV_X1    g176(.A(G169gat), .ZN(new_n378));
  INV_X1    g177(.A(G176gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT23), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT23), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(G169gat), .B2(G176gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(G169gat), .A2(G176gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n380), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n373), .B1(new_n377), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT64), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g186(.A(KEYINPUT64), .B(new_n373), .C1(new_n377), .C2(new_n384), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT25), .B1(new_n383), .B2(KEYINPUT65), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n383), .A2(KEYINPUT65), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n380), .A2(new_n390), .A3(new_n382), .ZN(new_n391));
  OR3_X1    g190(.A1(new_n377), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n387), .A2(new_n388), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(G183gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT27), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT27), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(G183gat), .ZN(new_n397));
  INV_X1    g196(.A(G190gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n395), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT66), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n399), .A2(new_n400), .A3(KEYINPUT28), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT28), .B1(new_n399), .B2(new_n400), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT67), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT26), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT26), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n406), .A2(new_n378), .A3(new_n379), .A4(KEYINPUT67), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n383), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G183gat), .A2(G190gat), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n408), .A2(KEYINPUT68), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT68), .B1(new_n408), .B2(new_n409), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n403), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G226gat), .A2(G233gat), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n393), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT29), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n417), .B1(new_n393), .B2(new_n412), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n372), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n393), .A2(new_n412), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n416), .ZN(new_n421));
  INV_X1    g220(.A(new_n372), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n393), .A2(new_n412), .A3(new_n413), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G8gat), .B(G36gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(G64gat), .B(G92gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  NAND3_X1  g226(.A1(new_n419), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT72), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n419), .A2(new_n424), .A3(KEYINPUT72), .A4(new_n427), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n419), .A2(new_n424), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT86), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n434), .B(KEYINPUT37), .C1(KEYINPUT86), .C2(new_n419), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT37), .ZN(new_n436));
  AOI211_X1 g235(.A(KEYINPUT38), .B(new_n427), .C1(new_n433), .C2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n432), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT87), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n436), .B1(new_n419), .B2(new_n424), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n439), .B1(new_n440), .B2(new_n427), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n433), .A2(new_n436), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n440), .A2(new_n439), .A3(new_n427), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT38), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n360), .A2(new_n438), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n322), .B1(new_n344), .B2(new_n321), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT39), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n340), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT39), .B1(new_n330), .B2(new_n331), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT84), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT84), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n452), .B(KEYINPUT39), .C1(new_n330), .C2(new_n331), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n316), .B1(new_n293), .B2(new_n313), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n454), .A2(new_n341), .A3(new_n343), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n451), .B(new_n453), .C1(new_n455), .C2(new_n322), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n449), .A2(KEYINPUT40), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT40), .B1(new_n449), .B2(new_n456), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n457), .A2(new_n458), .A3(new_n349), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT73), .B(KEYINPUT30), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n430), .A2(new_n431), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT30), .ZN(new_n462));
  OR3_X1    g261(.A1(new_n428), .A2(KEYINPUT71), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n427), .B1(new_n419), .B2(new_n424), .ZN(new_n464));
  OAI22_X1  g263(.A1(new_n464), .A2(KEYINPUT71), .B1(new_n428), .B2(new_n462), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n461), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n459), .A2(KEYINPUT85), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT85), .B1(new_n459), .B2(new_n466), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n446), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  XOR2_X1   g268(.A(G78gat), .B(G106gat), .Z(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(KEYINPUT81), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(G22gat), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT31), .B(G50gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(G228gat), .A2(G233gat), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT83), .B1(new_n422), .B2(new_n415), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n368), .A2(KEYINPUT83), .A3(new_n415), .A4(new_n371), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n318), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n292), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n422), .B1(new_n415), .B2(new_n319), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n475), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT29), .B1(new_n369), .B2(new_n366), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(new_n369), .B2(new_n366), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT82), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT3), .B1(new_n484), .B2(new_n485), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n307), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n475), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n488), .A2(new_n480), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n474), .B1(new_n482), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NOR3_X1   g291(.A1(new_n482), .A2(new_n490), .A3(new_n474), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n473), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n493), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(new_n491), .A3(new_n472), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n469), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT80), .B1(new_n360), .B2(new_n466), .ZN(new_n500));
  INV_X1    g299(.A(new_n466), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT80), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n501), .A2(new_n502), .A3(new_n359), .A4(new_n350), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n497), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(G15gat), .B(G43gat), .Z(new_n508));
  XNOR2_X1  g307(.A(G71gat), .B(G99gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n393), .A2(new_n412), .A3(new_n280), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n280), .B1(new_n393), .B2(new_n412), .ZN(new_n512));
  INV_X1    g311(.A(G227gat), .ZN(new_n513));
  INV_X1    g312(.A(G233gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n511), .A2(new_n512), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n510), .B1(new_n517), .B2(KEYINPUT33), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n511), .A2(new_n512), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT34), .B1(new_n519), .B2(new_n515), .ZN(new_n520));
  INV_X1    g319(.A(new_n280), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n420), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n393), .A2(new_n412), .A3(new_n280), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT34), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n525), .A3(new_n516), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n518), .A2(new_n520), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n510), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n522), .A2(new_n515), .A3(new_n523), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT33), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n525), .B1(new_n524), .B2(new_n516), .ZN(new_n532));
  AOI211_X1 g331(.A(KEYINPUT34), .B(new_n515), .C1(new_n522), .C2(new_n523), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n529), .A2(KEYINPUT32), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n527), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n536), .B1(new_n527), .B2(new_n534), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT36), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n527), .A2(new_n534), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n535), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT36), .B1(new_n543), .B2(new_n537), .ZN(new_n544));
  OAI22_X1  g343(.A1(new_n499), .A2(new_n507), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n497), .A2(new_n537), .A3(new_n543), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT35), .ZN(new_n548));
  INV_X1    g347(.A(new_n360), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n501), .A4(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n546), .B1(new_n500), .B2(new_n503), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n550), .B1(new_n551), .B2(new_n548), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n264), .B1(new_n545), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  OR2_X1    g353(.A1(G57gat), .A2(G64gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(G57gat), .A2(G64gat), .ZN(new_n556));
  AND2_X1   g355(.A1(G71gat), .A2(G78gat), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n555), .B(new_n556), .C1(new_n557), .C2(KEYINPUT9), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n557), .A2(KEYINPUT91), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(G71gat), .A2(G78gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n558), .B(new_n559), .C1(new_n557), .C2(new_n561), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n229), .B1(KEYINPUT21), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n565), .ZN(new_n567));
  NAND2_X1  g366(.A1(G231gat), .A2(G233gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT92), .B(KEYINPUT21), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n568), .B1(new_n567), .B2(new_n569), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n271), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n572), .A2(new_n271), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n566), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n575), .ZN(new_n577));
  INV_X1    g376(.A(new_n566), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(new_n578), .A3(new_n573), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(new_n301), .ZN(new_n582));
  XNOR2_X1  g381(.A(G183gat), .B(G211gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n582), .B(new_n583), .Z(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n576), .A2(new_n579), .A3(new_n584), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n591));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G190gat), .B(G218gat), .Z(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G85gat), .A2(G92gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT7), .ZN(new_n598));
  NOR2_X1   g397(.A1(G85gat), .A2(G92gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(G99gat), .A2(G106gat), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n599), .B1(KEYINPUT8), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(G99gat), .B(G106gat), .Z(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n605), .A2(new_n598), .A3(new_n601), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(KEYINPUT93), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT93), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n602), .A2(new_n608), .A3(new_n603), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n249), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n609), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n223), .A2(new_n612), .B1(KEYINPUT41), .B2(new_n590), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n596), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n612), .B1(new_n239), .B2(new_n243), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n616), .B1(new_n610), .B2(new_n232), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n615), .A2(new_n617), .A3(new_n595), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n594), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n611), .A2(new_n596), .A3(new_n613), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n595), .B1(new_n615), .B2(new_n617), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n620), .A2(new_n621), .A3(new_n593), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(KEYINPUT94), .B1(new_n589), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT94), .ZN(new_n625));
  INV_X1    g424(.A(new_n623), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n588), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(G230gat), .A2(G233gat), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT10), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n565), .B1(new_n607), .B2(new_n609), .ZN(new_n631));
  AOI22_X1  g430(.A1(new_n604), .A2(new_n606), .B1(new_n563), .B2(new_n564), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n612), .A2(KEYINPUT10), .A3(new_n565), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n629), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OR3_X1    g435(.A1(new_n631), .A2(new_n628), .A3(new_n632), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G120gat), .B(G148gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT95), .ZN(new_n640));
  XNOR2_X1  g439(.A(G176gat), .B(G204gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n640), .B(new_n641), .Z(new_n642));
  NAND2_X1  g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n642), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n636), .A2(new_n637), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n624), .A2(new_n627), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n360), .B(KEYINPUT96), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n554), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(new_n225), .ZN(G1324gat));
  NOR2_X1   g451(.A1(new_n554), .A2(new_n648), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n466), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT16), .B(G8gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT97), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT42), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n659), .B1(new_n654), .B2(G8gat), .ZN(new_n660));
  NOR2_X1   g459(.A1(KEYINPUT98), .A2(KEYINPUT42), .ZN(new_n661));
  MUX2_X1   g460(.A(KEYINPUT98), .B(new_n661), .S(new_n657), .Z(new_n662));
  AOI22_X1  g461(.A1(new_n658), .A2(new_n660), .B1(new_n655), .B2(new_n662), .ZN(G1325gat));
  INV_X1    g462(.A(new_n653), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT99), .B1(new_n541), .B2(new_n544), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n540), .B1(new_n538), .B2(new_n539), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n543), .A2(KEYINPUT36), .A3(new_n537), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT99), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(G15gat), .B1(new_n664), .B2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n538), .A2(new_n539), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n674), .A2(G15gat), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n672), .B1(new_n664), .B2(new_n675), .ZN(G1326gat));
  NAND2_X1  g475(.A1(new_n653), .A2(new_n505), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT43), .B(G22gat), .Z(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n678), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n653), .A2(new_n505), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n682), .B(new_n684), .ZN(G1327gat));
  NOR2_X1   g484(.A1(new_n588), .A2(new_n646), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n553), .A2(new_n623), .A3(new_n686), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n687), .A2(G29gat), .A3(new_n650), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT45), .Z(new_n689));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n670), .B1(new_n498), .B2(new_n506), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n552), .A2(KEYINPUT103), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n550), .B(new_n693), .C1(new_n551), .C2(new_n548), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n691), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n690), .B1(new_n695), .B2(new_n626), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n545), .A2(new_n552), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n626), .A2(new_n690), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n259), .B1(new_n248), .B2(new_n253), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n261), .A2(new_n258), .A3(new_n262), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n701), .A2(new_n702), .A3(KEYINPUT102), .ZN(new_n703));
  AOI21_X1  g502(.A(KEYINPUT102), .B1(new_n701), .B2(new_n702), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n686), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n700), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(G29gat), .B1(new_n709), .B2(new_n650), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n689), .A2(new_n710), .ZN(G1328gat));
  NOR3_X1   g510(.A1(new_n687), .A2(G36gat), .A3(new_n501), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT46), .ZN(new_n713));
  OAI21_X1  g512(.A(G36gat), .B1(new_n709), .B2(new_n501), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(G1329gat));
  NOR3_X1   g514(.A1(new_n687), .A2(G43gat), .A3(new_n674), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n670), .A3(new_n708), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n716), .B1(new_n717), .B2(G43gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g518(.A1(new_n207), .A2(new_n209), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n505), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n687), .A2(new_n497), .ZN(new_n722));
  OAI22_X1  g521(.A1(new_n709), .A2(new_n721), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g523(.A1(new_n692), .A2(new_n694), .ZN(new_n725));
  INV_X1    g524(.A(new_n691), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AND4_X1   g526(.A1(new_n624), .A2(new_n706), .A3(new_n627), .A4(new_n646), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n649), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g531(.A1(new_n729), .A2(new_n501), .ZN(new_n733));
  NOR2_X1   g532(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n734));
  AND2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n733), .B2(new_n734), .ZN(G1333gat));
  OR3_X1    g536(.A1(new_n729), .A2(G71gat), .A3(new_n674), .ZN(new_n738));
  OAI21_X1  g537(.A(G71gat), .B1(new_n729), .B2(new_n671), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g540(.A1(new_n730), .A2(new_n505), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g542(.A1(new_n705), .A2(new_n588), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(new_n647), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n696), .A2(new_n649), .A3(new_n699), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G85gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n727), .A2(new_n623), .A3(new_n744), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT51), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n695), .A2(new_n626), .A3(new_n745), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(G85gat), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n649), .A2(new_n755), .A3(new_n646), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n748), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1336gat));
  NOR2_X1   g558(.A1(KEYINPUT105), .A2(KEYINPUT51), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n749), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n760), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n751), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n501), .A2(G92gat), .A3(new_n647), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n696), .A2(new_n466), .A3(new_n699), .A4(new_n746), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G92gat), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT52), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n626), .B1(new_n725), .B2(new_n726), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n752), .B1(new_n771), .B2(new_n744), .ZN(new_n772));
  NOR4_X1   g571(.A1(new_n695), .A2(KEYINPUT51), .A3(new_n626), .A4(new_n745), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT52), .B1(new_n774), .B2(new_n765), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT106), .B1(new_n775), .B2(new_n768), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n750), .A2(new_n753), .A3(new_n765), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  AND4_X1   g577(.A1(KEYINPUT106), .A2(new_n777), .A3(new_n768), .A4(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n770), .B1(new_n776), .B2(new_n779), .ZN(G1337gat));
  NAND3_X1  g579(.A1(new_n700), .A2(new_n670), .A3(new_n746), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G99gat), .ZN(new_n782));
  OR3_X1    g581(.A1(new_n674), .A2(G99gat), .A3(new_n647), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n754), .B2(new_n783), .ZN(G1338gat));
  NOR3_X1   g583(.A1(new_n497), .A2(G106gat), .A3(new_n647), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n750), .A2(new_n753), .A3(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n696), .A2(new_n505), .A3(new_n699), .A4(new_n746), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G106gat), .ZN(new_n788));
  XNOR2_X1  g587(.A(KEYINPUT107), .B(KEYINPUT53), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n786), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n762), .B1(new_n771), .B2(new_n744), .ZN(new_n792));
  NOR4_X1   g591(.A1(new_n695), .A2(new_n626), .A3(new_n745), .A4(new_n760), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n785), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n791), .B1(new_n794), .B2(new_n788), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT108), .B1(new_n790), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT108), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n786), .A2(new_n788), .A3(new_n789), .ZN(new_n798));
  AOI22_X1  g597(.A1(new_n764), .A2(new_n785), .B1(G106gat), .B2(new_n787), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n797), .B(new_n798), .C1(new_n799), .C2(new_n791), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n796), .A2(new_n800), .ZN(G1339gat));
  NAND4_X1  g600(.A1(new_n624), .A2(new_n706), .A3(new_n627), .A4(new_n647), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n633), .A2(new_n629), .A3(new_n634), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n636), .A2(KEYINPUT54), .A3(new_n804), .ZN(new_n805));
  XOR2_X1   g604(.A(KEYINPUT109), .B(KEYINPUT54), .Z(new_n806));
  AOI21_X1  g605(.A(new_n644), .B1(new_n635), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n805), .A2(KEYINPUT55), .A3(new_n807), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(new_n645), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n235), .B1(new_n250), .B2(new_n230), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n234), .A2(new_n236), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n257), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n623), .A2(new_n702), .A3(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n812), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n702), .A2(new_n815), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n705), .A2(new_n819), .B1(new_n646), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n818), .B1(new_n821), .B2(new_n623), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n588), .B1(new_n822), .B2(KEYINPUT110), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT110), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n824), .B(new_n818), .C1(new_n821), .C2(new_n623), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n803), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(new_n650), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n828), .A3(new_n547), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT102), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(new_n260), .B2(new_n263), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n701), .A2(new_n702), .A3(KEYINPUT102), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n811), .A2(new_n645), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n831), .A2(new_n832), .A3(new_n810), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n646), .A2(new_n702), .A3(new_n815), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n623), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT110), .B1(new_n836), .B2(new_n817), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n825), .A2(new_n837), .A3(new_n589), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n802), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(new_n547), .A3(new_n649), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT113), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n829), .A2(new_n501), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(new_n268), .A3(new_n705), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n650), .A2(new_n466), .A3(new_n674), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n839), .A2(new_n497), .A3(new_n845), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT111), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n701), .A2(new_n702), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n850), .A2(KEYINPUT112), .A3(G113gat), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT112), .B1(new_n850), .B2(G113gat), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n844), .B1(new_n851), .B2(new_n852), .ZN(G1340gat));
  NOR3_X1   g652(.A1(new_n847), .A2(new_n266), .A3(new_n647), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n843), .A2(new_n646), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n855), .B2(new_n266), .ZN(G1341gat));
  OAI21_X1  g655(.A(G127gat), .B1(new_n847), .B2(new_n589), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n588), .A2(new_n271), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(new_n842), .B2(new_n858), .ZN(G1342gat));
  OAI21_X1  g658(.A(G134gat), .B1(new_n847), .B2(new_n626), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT114), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n862), .B(G134gat), .C1(new_n847), .C2(new_n626), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n623), .A2(new_n273), .ZN(new_n865));
  OR3_X1    g664(.A1(new_n842), .A2(KEYINPUT56), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT56), .B1(new_n842), .B2(new_n865), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n867), .A2(KEYINPUT115), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n867), .A2(KEYINPUT115), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n864), .B(new_n866), .C1(new_n868), .C2(new_n869), .ZN(G1343gat));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n871), .B(new_n872), .C1(new_n826), .C2(new_n497), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n497), .B1(new_n838), .B2(new_n802), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT116), .B1(new_n874), .B2(KEYINPUT57), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n835), .B1(new_n812), .B2(new_n264), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n817), .B1(new_n877), .B2(new_n626), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n876), .B1(new_n878), .B2(new_n588), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n833), .A2(new_n849), .A3(new_n810), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n623), .B1(new_n880), .B2(new_n835), .ZN(new_n881));
  OAI211_X1 g680(.A(KEYINPUT117), .B(new_n589), .C1(new_n881), .C2(new_n817), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n879), .A2(new_n802), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n497), .A2(new_n872), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n883), .A2(KEYINPUT118), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT118), .B1(new_n883), .B2(new_n884), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n873), .A2(new_n875), .A3(new_n887), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n650), .A2(new_n670), .A3(new_n466), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n849), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(G141gat), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT58), .ZN(new_n892));
  AND4_X1   g691(.A1(new_n505), .A2(new_n827), .A3(new_n501), .A4(new_n671), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n304), .A3(new_n849), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n891), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n888), .A2(new_n705), .A3(new_n889), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(G141gat), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n897), .A2(new_n894), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n895), .B1(new_n898), .B2(new_n892), .ZN(G1344gat));
  NAND3_X1  g698(.A1(new_n893), .A2(new_n288), .A3(new_n646), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n888), .A2(new_n646), .A3(new_n889), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n288), .A2(KEYINPUT59), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n589), .B1(new_n881), .B2(new_n817), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n904), .B1(new_n648), .B2(new_n849), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n497), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n904), .B(KEYINPUT119), .C1(new_n648), .C2(new_n849), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT57), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n884), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n910), .B1(new_n838), .B2(new_n802), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n646), .B(new_n889), .C1(new_n909), .C2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(G148gat), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n913), .A2(KEYINPUT59), .ZN(new_n914));
  OAI211_X1 g713(.A(KEYINPUT120), .B(new_n900), .C1(new_n903), .C2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n916));
  AOI22_X1  g715(.A1(new_n901), .A2(new_n902), .B1(KEYINPUT59), .B2(new_n913), .ZN(new_n917));
  INV_X1    g716(.A(new_n900), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n915), .A2(new_n919), .ZN(G1345gat));
  AOI21_X1  g719(.A(G155gat), .B1(new_n893), .B2(new_n588), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n888), .A2(new_n889), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n588), .A2(G155gat), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT121), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n921), .B1(new_n922), .B2(new_n924), .ZN(G1346gat));
  AOI21_X1  g724(.A(G162gat), .B1(new_n893), .B2(new_n623), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n626), .A2(new_n302), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n926), .B1(new_n922), .B2(new_n927), .ZN(G1347gat));
  NOR2_X1   g727(.A1(new_n826), .A2(new_n649), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n546), .A2(new_n501), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT122), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(G169gat), .B1(new_n933), .B2(new_n705), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n839), .A2(new_n497), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n650), .A2(new_n466), .A3(new_n673), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n264), .A2(new_n378), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(G1348gat));
  NAND3_X1  g738(.A1(new_n933), .A2(new_n379), .A3(new_n646), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n935), .A2(new_n647), .A3(new_n936), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n379), .B2(new_n941), .ZN(G1349gat));
  INV_X1    g741(.A(KEYINPUT124), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n395), .A2(new_n397), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n588), .A2(new_n944), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n935), .A2(new_n589), .A3(new_n936), .ZN(new_n946));
  OAI221_X1 g745(.A(new_n943), .B1(new_n932), .B2(new_n945), .C1(new_n394), .C2(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n932), .A2(new_n945), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n394), .B1(new_n937), .B2(new_n588), .ZN(new_n949));
  OAI21_X1  g748(.A(KEYINPUT124), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AND4_X1   g749(.A1(KEYINPUT123), .A2(new_n947), .A3(new_n950), .A4(KEYINPUT60), .ZN(new_n951));
  AOI22_X1  g750(.A1(new_n947), .A2(new_n950), .B1(KEYINPUT123), .B2(KEYINPUT60), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(G1350gat));
  AOI21_X1  g752(.A(new_n398), .B1(new_n937), .B2(new_n623), .ZN(new_n954));
  XOR2_X1   g753(.A(new_n954), .B(KEYINPUT61), .Z(new_n955));
  NAND3_X1  g754(.A1(new_n933), .A2(new_n398), .A3(new_n623), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1351gat));
  OR2_X1    g756(.A1(new_n909), .A2(new_n911), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n670), .A2(new_n501), .A3(new_n649), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(KEYINPUT126), .B1(new_n960), .B2(new_n264), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(G197gat), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n960), .A2(KEYINPUT126), .A3(new_n264), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n670), .A2(new_n497), .A3(new_n501), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT125), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n929), .A2(new_n965), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n706), .A2(G197gat), .ZN(new_n967));
  OAI22_X1  g766(.A1(new_n962), .A2(new_n963), .B1(new_n966), .B2(new_n967), .ZN(G1352gat));
  INV_X1    g767(.A(new_n960), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n969), .A2(KEYINPUT127), .A3(new_n646), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n971), .B1(new_n960), .B2(new_n647), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n970), .A2(G204gat), .A3(new_n972), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n966), .A2(G204gat), .A3(new_n647), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT62), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n975), .ZN(G1353gat));
  OR3_X1    g775(.A1(new_n966), .A2(G211gat), .A3(new_n589), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n969), .A2(new_n588), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n978), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT63), .B1(new_n978), .B2(G211gat), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(G1354gat));
  OAI21_X1  g780(.A(G218gat), .B1(new_n960), .B2(new_n626), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n626), .A2(G218gat), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n982), .B1(new_n966), .B2(new_n983), .ZN(G1355gat));
endmodule


