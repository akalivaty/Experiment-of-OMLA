

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U557 ( .A1(n703), .A2(n604), .ZN(n641) );
  XOR2_X1 U558 ( .A(n622), .B(KEYINPUT26), .Z(n521) );
  AND2_X1 U559 ( .A1(n641), .A2(G1996), .ZN(n622) );
  NOR2_X1 U560 ( .A1(n982), .A2(n624), .ZN(n638) );
  INV_X1 U561 ( .A(n704), .ZN(n604) );
  XNOR2_X1 U562 ( .A(n603), .B(KEYINPUT64), .ZN(n703) );
  NOR2_X1 U563 ( .A1(G651), .A2(n565), .ZN(n783) );
  NOR2_X1 U564 ( .A1(n548), .A2(n547), .ZN(G160) );
  XOR2_X1 U565 ( .A(G543), .B(KEYINPUT0), .Z(n565) );
  INV_X1 U566 ( .A(G651), .ZN(n529) );
  NOR2_X1 U567 ( .A1(n565), .A2(n529), .ZN(n782) );
  NAND2_X1 U568 ( .A1(n782), .A2(G76), .ZN(n522) );
  XNOR2_X1 U569 ( .A(KEYINPUT77), .B(n522), .ZN(n525) );
  NOR2_X1 U570 ( .A1(G543), .A2(G651), .ZN(n778) );
  NAND2_X1 U571 ( .A1(n778), .A2(G89), .ZN(n523) );
  XOR2_X1 U572 ( .A(n523), .B(KEYINPUT4), .Z(n524) );
  NOR2_X1 U573 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U574 ( .A(KEYINPUT78), .B(n526), .Z(n527) );
  XNOR2_X1 U575 ( .A(KEYINPUT5), .B(n527), .ZN(n535) );
  NAND2_X1 U576 ( .A1(n783), .A2(G51), .ZN(n528) );
  XOR2_X1 U577 ( .A(KEYINPUT79), .B(n528), .Z(n532) );
  NOR2_X1 U578 ( .A1(G543), .A2(n529), .ZN(n530) );
  XOR2_X1 U579 ( .A(KEYINPUT1), .B(n530), .Z(n779) );
  NAND2_X1 U580 ( .A1(n779), .A2(G63), .ZN(n531) );
  NAND2_X1 U581 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U582 ( .A(KEYINPUT6), .B(n533), .Z(n534) );
  NAND2_X1 U583 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U584 ( .A(n536), .B(KEYINPUT7), .ZN(n537) );
  XNOR2_X1 U585 ( .A(KEYINPUT80), .B(n537), .ZN(G168) );
  XOR2_X1 U586 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  AND2_X1 U587 ( .A1(G2105), .A2(G2104), .ZN(n871) );
  NAND2_X1 U588 ( .A1(n871), .A2(G113), .ZN(n540) );
  INV_X1 U589 ( .A(G2104), .ZN(n541) );
  AND2_X1 U590 ( .A1(n541), .A2(G2105), .ZN(n870) );
  NAND2_X1 U591 ( .A1(G125), .A2(n870), .ZN(n538) );
  XOR2_X1 U592 ( .A(KEYINPUT65), .B(n538), .Z(n539) );
  NAND2_X1 U593 ( .A1(n540), .A2(n539), .ZN(n548) );
  NOR2_X4 U594 ( .A1(G2105), .A2(n541), .ZN(n864) );
  NAND2_X1 U595 ( .A1(G101), .A2(n864), .ZN(n542) );
  XOR2_X1 U596 ( .A(KEYINPUT66), .B(n542), .Z(n543) );
  XNOR2_X1 U597 ( .A(n543), .B(KEYINPUT23), .ZN(n546) );
  NOR2_X1 U598 ( .A1(G2105), .A2(G2104), .ZN(n544) );
  XOR2_X2 U599 ( .A(KEYINPUT17), .B(n544), .Z(n865) );
  NAND2_X1 U600 ( .A1(G137), .A2(n865), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U602 ( .A1(G48), .A2(n783), .ZN(n549) );
  XNOR2_X1 U603 ( .A(n549), .B(KEYINPUT86), .ZN(n556) );
  NAND2_X1 U604 ( .A1(G86), .A2(n778), .ZN(n551) );
  NAND2_X1 U605 ( .A1(G61), .A2(n779), .ZN(n550) );
  NAND2_X1 U606 ( .A1(n551), .A2(n550), .ZN(n554) );
  NAND2_X1 U607 ( .A1(n782), .A2(G73), .ZN(n552) );
  XOR2_X1 U608 ( .A(KEYINPUT2), .B(n552), .Z(n553) );
  NOR2_X1 U609 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U610 ( .A1(n556), .A2(n555), .ZN(G305) );
  NAND2_X1 U611 ( .A1(G138), .A2(n865), .ZN(n558) );
  NAND2_X1 U612 ( .A1(G102), .A2(n864), .ZN(n557) );
  NAND2_X1 U613 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U614 ( .A1(G126), .A2(n870), .ZN(n560) );
  NAND2_X1 U615 ( .A1(G114), .A2(n871), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U617 ( .A1(n562), .A2(n561), .ZN(G164) );
  NAND2_X1 U618 ( .A1(G74), .A2(G651), .ZN(n563) );
  XOR2_X1 U619 ( .A(KEYINPUT84), .B(n563), .Z(n564) );
  NOR2_X1 U620 ( .A1(n779), .A2(n564), .ZN(n567) );
  NAND2_X1 U621 ( .A1(n565), .A2(G87), .ZN(n566) );
  NAND2_X1 U622 ( .A1(n567), .A2(n566), .ZN(n570) );
  NAND2_X1 U623 ( .A1(G49), .A2(n783), .ZN(n568) );
  XNOR2_X1 U624 ( .A(KEYINPUT83), .B(n568), .ZN(n569) );
  NOR2_X1 U625 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U626 ( .A(KEYINPUT85), .B(n571), .ZN(G288) );
  NAND2_X1 U627 ( .A1(G64), .A2(n779), .ZN(n572) );
  XNOR2_X1 U628 ( .A(n572), .B(KEYINPUT69), .ZN(n579) );
  NAND2_X1 U629 ( .A1(G77), .A2(n782), .ZN(n574) );
  NAND2_X1 U630 ( .A1(G90), .A2(n778), .ZN(n573) );
  NAND2_X1 U631 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U632 ( .A(n575), .B(KEYINPUT9), .ZN(n577) );
  NAND2_X1 U633 ( .A1(G52), .A2(n783), .ZN(n576) );
  NAND2_X1 U634 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U635 ( .A1(n579), .A2(n578), .ZN(G171) );
  NAND2_X1 U636 ( .A1(G78), .A2(n782), .ZN(n581) );
  NAND2_X1 U637 ( .A1(G91), .A2(n778), .ZN(n580) );
  NAND2_X1 U638 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U639 ( .A1(n779), .A2(G65), .ZN(n582) );
  XOR2_X1 U640 ( .A(KEYINPUT70), .B(n582), .Z(n583) );
  NOR2_X1 U641 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U642 ( .A1(n783), .A2(G53), .ZN(n585) );
  NAND2_X1 U643 ( .A1(n586), .A2(n585), .ZN(G299) );
  NAND2_X1 U644 ( .A1(G75), .A2(n782), .ZN(n588) );
  NAND2_X1 U645 ( .A1(G88), .A2(n778), .ZN(n587) );
  NAND2_X1 U646 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U647 ( .A1(G62), .A2(n779), .ZN(n589) );
  XNOR2_X1 U648 ( .A(KEYINPUT87), .B(n589), .ZN(n590) );
  NOR2_X1 U649 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U650 ( .A1(n783), .A2(G50), .ZN(n592) );
  NAND2_X1 U651 ( .A1(n593), .A2(n592), .ZN(G303) );
  NAND2_X1 U652 ( .A1(G60), .A2(n779), .ZN(n594) );
  XNOR2_X1 U653 ( .A(n594), .B(KEYINPUT68), .ZN(n596) );
  NAND2_X1 U654 ( .A1(n782), .A2(G72), .ZN(n595) );
  NAND2_X1 U655 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U656 ( .A1(G85), .A2(n778), .ZN(n597) );
  XNOR2_X1 U657 ( .A(KEYINPUT67), .B(n597), .ZN(n598) );
  NOR2_X1 U658 ( .A1(n599), .A2(n598), .ZN(n601) );
  NAND2_X1 U659 ( .A1(n783), .A2(G47), .ZN(n600) );
  NAND2_X1 U660 ( .A1(n601), .A2(n600), .ZN(G290) );
  XNOR2_X1 U661 ( .A(KEYINPUT106), .B(G1981), .ZN(n602) );
  XNOR2_X1 U662 ( .A(n602), .B(G305), .ZN(n689) );
  NOR2_X1 U663 ( .A1(G1384), .A2(G164), .ZN(n603) );
  NAND2_X1 U664 ( .A1(G160), .A2(G40), .ZN(n704) );
  INV_X1 U665 ( .A(n641), .ZN(n664) );
  NAND2_X1 U666 ( .A1(G8), .A2(n664), .ZN(n700) );
  NOR2_X1 U667 ( .A1(G1976), .A2(G288), .ZN(n691) );
  XNOR2_X1 U668 ( .A(KEYINPUT105), .B(n691), .ZN(n605) );
  NOR2_X1 U669 ( .A1(n700), .A2(n605), .ZN(n606) );
  NOR2_X1 U670 ( .A1(n689), .A2(n606), .ZN(n607) );
  NAND2_X1 U671 ( .A1(n607), .A2(KEYINPUT33), .ZN(n686) );
  OR2_X1 U672 ( .A1(n641), .A2(G1961), .ZN(n610) );
  XNOR2_X1 U673 ( .A(G2078), .B(KEYINPUT100), .ZN(n608) );
  XNOR2_X1 U674 ( .A(n608), .B(KEYINPUT25), .ZN(n947) );
  NAND2_X1 U675 ( .A1(n641), .A2(n947), .ZN(n609) );
  NAND2_X1 U676 ( .A1(n610), .A2(n609), .ZN(n658) );
  NAND2_X1 U677 ( .A1(n658), .A2(G171), .ZN(n653) );
  NAND2_X1 U678 ( .A1(n779), .A2(G56), .ZN(n611) );
  XNOR2_X1 U679 ( .A(KEYINPUT14), .B(n611), .ZN(n617) );
  NAND2_X1 U680 ( .A1(n778), .A2(G81), .ZN(n612) );
  XNOR2_X1 U681 ( .A(n612), .B(KEYINPUT12), .ZN(n614) );
  NAND2_X1 U682 ( .A1(G68), .A2(n782), .ZN(n613) );
  NAND2_X1 U683 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U684 ( .A(KEYINPUT13), .B(n615), .ZN(n616) );
  NAND2_X1 U685 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U686 ( .A(n618), .B(KEYINPUT73), .ZN(n620) );
  NAND2_X1 U687 ( .A1(n783), .A2(G43), .ZN(n619) );
  NAND2_X1 U688 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U689 ( .A(KEYINPUT74), .B(n621), .ZN(n982) );
  NAND2_X1 U690 ( .A1(n664), .A2(G1341), .ZN(n623) );
  NAND2_X1 U691 ( .A1(n521), .A2(n623), .ZN(n624) );
  NAND2_X1 U692 ( .A1(G92), .A2(n778), .ZN(n626) );
  NAND2_X1 U693 ( .A1(G66), .A2(n779), .ZN(n625) );
  NAND2_X1 U694 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U695 ( .A1(G79), .A2(n782), .ZN(n628) );
  NAND2_X1 U696 ( .A1(G54), .A2(n783), .ZN(n627) );
  NAND2_X1 U697 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U698 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U699 ( .A(KEYINPUT15), .B(n631), .Z(n893) );
  NAND2_X1 U700 ( .A1(n638), .A2(n893), .ZN(n636) );
  INV_X1 U701 ( .A(G2067), .ZN(n944) );
  NOR2_X1 U702 ( .A1(n664), .A2(n944), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n632), .B(KEYINPUT101), .ZN(n634) );
  NAND2_X1 U704 ( .A1(n664), .A2(G1348), .ZN(n633) );
  NAND2_X1 U705 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U706 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U707 ( .A(n637), .B(KEYINPUT102), .ZN(n640) );
  OR2_X1 U708 ( .A1(n638), .A2(n893), .ZN(n639) );
  NAND2_X1 U709 ( .A1(n640), .A2(n639), .ZN(n646) );
  INV_X1 U710 ( .A(G299), .ZN(n975) );
  NAND2_X1 U711 ( .A1(n641), .A2(G2072), .ZN(n642) );
  XNOR2_X1 U712 ( .A(n642), .B(KEYINPUT27), .ZN(n644) );
  AND2_X1 U713 ( .A1(G1956), .A2(n664), .ZN(n643) );
  NOR2_X1 U714 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U715 ( .A1(n975), .A2(n647), .ZN(n645) );
  NAND2_X1 U716 ( .A1(n646), .A2(n645), .ZN(n650) );
  NOR2_X1 U717 ( .A1(n975), .A2(n647), .ZN(n648) );
  XOR2_X1 U718 ( .A(n648), .B(KEYINPUT28), .Z(n649) );
  NAND2_X1 U719 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U720 ( .A(n651), .B(KEYINPUT29), .Z(n652) );
  NAND2_X1 U721 ( .A1(n653), .A2(n652), .ZN(n663) );
  NOR2_X1 U722 ( .A1(G1966), .A2(n700), .ZN(n677) );
  NOR2_X1 U723 ( .A1(n664), .A2(G2084), .ZN(n654) );
  XNOR2_X1 U724 ( .A(n654), .B(KEYINPUT99), .ZN(n673) );
  NAND2_X1 U725 ( .A1(G8), .A2(n673), .ZN(n655) );
  NOR2_X1 U726 ( .A1(n677), .A2(n655), .ZN(n656) );
  XOR2_X1 U727 ( .A(KEYINPUT30), .B(n656), .Z(n657) );
  NOR2_X1 U728 ( .A1(G168), .A2(n657), .ZN(n660) );
  NOR2_X1 U729 ( .A1(G171), .A2(n658), .ZN(n659) );
  NOR2_X1 U730 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U731 ( .A(KEYINPUT31), .B(n661), .Z(n662) );
  NAND2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n675) );
  NAND2_X1 U733 ( .A1(n675), .A2(G286), .ZN(n670) );
  NOR2_X1 U734 ( .A1(G1971), .A2(n700), .ZN(n666) );
  NOR2_X1 U735 ( .A1(G2090), .A2(n664), .ZN(n665) );
  NOR2_X1 U736 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U737 ( .A1(n667), .A2(G303), .ZN(n668) );
  XOR2_X1 U738 ( .A(KEYINPUT103), .B(n668), .Z(n669) );
  NAND2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U740 ( .A1(n671), .A2(G8), .ZN(n672) );
  XNOR2_X1 U741 ( .A(n672), .B(KEYINPUT32), .ZN(n681) );
  INV_X1 U742 ( .A(n673), .ZN(n674) );
  NAND2_X1 U743 ( .A1(G8), .A2(n674), .ZN(n679) );
  INV_X1 U744 ( .A(n675), .ZN(n676) );
  NOR2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U747 ( .A1(n681), .A2(n680), .ZN(n692) );
  NOR2_X1 U748 ( .A1(G2090), .A2(G303), .ZN(n682) );
  NAND2_X1 U749 ( .A1(G8), .A2(n682), .ZN(n683) );
  NAND2_X1 U750 ( .A1(n692), .A2(n683), .ZN(n684) );
  NAND2_X1 U751 ( .A1(n684), .A2(n700), .ZN(n685) );
  NAND2_X1 U752 ( .A1(n686), .A2(n685), .ZN(n702) );
  NOR2_X1 U753 ( .A1(G1981), .A2(G305), .ZN(n687) );
  XNOR2_X1 U754 ( .A(KEYINPUT24), .B(n687), .ZN(n698) );
  NAND2_X1 U755 ( .A1(G288), .A2(G1976), .ZN(n688) );
  XNOR2_X1 U756 ( .A(n688), .B(KEYINPUT104), .ZN(n976) );
  INV_X1 U757 ( .A(n689), .ZN(n965) );
  NAND2_X1 U758 ( .A1(n976), .A2(n965), .ZN(n696) );
  NOR2_X1 U759 ( .A1(G1971), .A2(G303), .ZN(n690) );
  NOR2_X1 U760 ( .A1(n691), .A2(n690), .ZN(n968) );
  NAND2_X1 U761 ( .A1(n692), .A2(n968), .ZN(n694) );
  NOR2_X1 U762 ( .A1(KEYINPUT105), .A2(KEYINPUT33), .ZN(n693) );
  NAND2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U764 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U765 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U766 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U767 ( .A1(n702), .A2(n701), .ZN(n738) );
  NOR2_X1 U768 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U769 ( .A(KEYINPUT94), .B(n705), .Z(n751) );
  NAND2_X1 U770 ( .A1(G129), .A2(n870), .ZN(n707) );
  NAND2_X1 U771 ( .A1(G117), .A2(n871), .ZN(n706) );
  NAND2_X1 U772 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U773 ( .A(KEYINPUT98), .B(n708), .ZN(n711) );
  NAND2_X1 U774 ( .A1(n864), .A2(G105), .ZN(n709) );
  XOR2_X1 U775 ( .A(KEYINPUT38), .B(n709), .Z(n710) );
  NOR2_X1 U776 ( .A1(n711), .A2(n710), .ZN(n713) );
  NAND2_X1 U777 ( .A1(n865), .A2(G141), .ZN(n712) );
  NAND2_X1 U778 ( .A1(n713), .A2(n712), .ZN(n882) );
  AND2_X1 U779 ( .A1(n882), .A2(G1996), .ZN(n723) );
  NAND2_X1 U780 ( .A1(G131), .A2(n865), .ZN(n720) );
  NAND2_X1 U781 ( .A1(G119), .A2(n870), .ZN(n715) );
  NAND2_X1 U782 ( .A1(G107), .A2(n871), .ZN(n714) );
  NAND2_X1 U783 ( .A1(n715), .A2(n714), .ZN(n718) );
  NAND2_X1 U784 ( .A1(n864), .A2(G95), .ZN(n716) );
  XOR2_X1 U785 ( .A(KEYINPUT96), .B(n716), .Z(n717) );
  NOR2_X1 U786 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U787 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U788 ( .A(n721), .B(KEYINPUT97), .ZN(n879) );
  INV_X1 U789 ( .A(G1991), .ZN(n940) );
  NOR2_X1 U790 ( .A1(n879), .A2(n940), .ZN(n722) );
  NOR2_X1 U791 ( .A1(n723), .A2(n722), .ZN(n929) );
  NOR2_X1 U792 ( .A1(n751), .A2(n929), .ZN(n743) );
  INV_X1 U793 ( .A(n743), .ZN(n736) );
  XOR2_X1 U794 ( .A(KEYINPUT37), .B(G2067), .Z(n739) );
  NAND2_X1 U795 ( .A1(G128), .A2(n870), .ZN(n725) );
  NAND2_X1 U796 ( .A1(G116), .A2(n871), .ZN(n724) );
  NAND2_X1 U797 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U798 ( .A(n726), .B(KEYINPUT35), .ZN(n731) );
  NAND2_X1 U799 ( .A1(G104), .A2(n864), .ZN(n728) );
  NAND2_X1 U800 ( .A1(G140), .A2(n865), .ZN(n727) );
  NAND2_X1 U801 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U802 ( .A(KEYINPUT34), .B(n729), .Z(n730) );
  NAND2_X1 U803 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U804 ( .A(n732), .B(KEYINPUT36), .ZN(n887) );
  NAND2_X1 U805 ( .A1(n739), .A2(n887), .ZN(n923) );
  NOR2_X1 U806 ( .A1(n751), .A2(n923), .ZN(n748) );
  XOR2_X1 U807 ( .A(G1986), .B(G290), .Z(n969) );
  NOR2_X1 U808 ( .A1(n969), .A2(n751), .ZN(n733) );
  XOR2_X1 U809 ( .A(KEYINPUT95), .B(n733), .Z(n734) );
  NOR2_X1 U810 ( .A1(n748), .A2(n734), .ZN(n735) );
  NAND2_X1 U811 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U812 ( .A1(n738), .A2(n737), .ZN(n753) );
  NOR2_X1 U813 ( .A1(n739), .A2(n887), .ZN(n935) );
  NOR2_X1 U814 ( .A1(G1996), .A2(n882), .ZN(n915) );
  NOR2_X1 U815 ( .A1(G1986), .A2(G290), .ZN(n741) );
  INV_X1 U816 ( .A(n879), .ZN(n740) );
  NOR2_X1 U817 ( .A1(G1991), .A2(n740), .ZN(n927) );
  NOR2_X1 U818 ( .A1(n741), .A2(n927), .ZN(n742) );
  NOR2_X1 U819 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U820 ( .A1(n915), .A2(n744), .ZN(n745) );
  XNOR2_X1 U821 ( .A(n745), .B(KEYINPUT107), .ZN(n746) );
  XNOR2_X1 U822 ( .A(KEYINPUT39), .B(n746), .ZN(n747) );
  NOR2_X1 U823 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U824 ( .A1(n935), .A2(n749), .ZN(n750) );
  NOR2_X1 U825 ( .A1(n751), .A2(n750), .ZN(n752) );
  OR2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U827 ( .A(n754), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U828 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U829 ( .A1(G111), .A2(n871), .ZN(n756) );
  NAND2_X1 U830 ( .A1(G135), .A2(n865), .ZN(n755) );
  NAND2_X1 U831 ( .A1(n756), .A2(n755), .ZN(n759) );
  NAND2_X1 U832 ( .A1(n870), .A2(G123), .ZN(n757) );
  XOR2_X1 U833 ( .A(KEYINPUT18), .B(n757), .Z(n758) );
  NOR2_X1 U834 ( .A1(n759), .A2(n758), .ZN(n761) );
  NAND2_X1 U835 ( .A1(n864), .A2(G99), .ZN(n760) );
  NAND2_X1 U836 ( .A1(n761), .A2(n760), .ZN(n924) );
  XNOR2_X1 U837 ( .A(G2096), .B(n924), .ZN(n762) );
  OR2_X1 U838 ( .A1(G2100), .A2(n762), .ZN(G156) );
  INV_X1 U839 ( .A(G57), .ZN(G237) );
  NAND2_X1 U840 ( .A1(G7), .A2(G661), .ZN(n763) );
  XNOR2_X1 U841 ( .A(n763), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U842 ( .A(G223), .ZN(n821) );
  NAND2_X1 U843 ( .A1(n821), .A2(G567), .ZN(n764) );
  XOR2_X1 U844 ( .A(KEYINPUT11), .B(n764), .Z(G234) );
  INV_X1 U845 ( .A(G860), .ZN(n771) );
  OR2_X1 U846 ( .A1(n771), .A2(n982), .ZN(n765) );
  XOR2_X1 U847 ( .A(KEYINPUT75), .B(n765), .Z(G153) );
  INV_X1 U848 ( .A(G171), .ZN(G301) );
  INV_X1 U849 ( .A(n893), .ZN(n970) );
  NOR2_X1 U850 ( .A1(G868), .A2(n970), .ZN(n767) );
  INV_X1 U851 ( .A(G868), .ZN(n800) );
  NOR2_X1 U852 ( .A1(n800), .A2(G301), .ZN(n766) );
  NOR2_X1 U853 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U854 ( .A(KEYINPUT76), .B(n768), .ZN(G284) );
  NAND2_X1 U855 ( .A1(G868), .A2(G286), .ZN(n770) );
  NAND2_X1 U856 ( .A1(G299), .A2(n800), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n770), .A2(n769), .ZN(G297) );
  NAND2_X1 U858 ( .A1(n771), .A2(G559), .ZN(n772) );
  NAND2_X1 U859 ( .A1(n772), .A2(n893), .ZN(n773) );
  XNOR2_X1 U860 ( .A(n773), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U861 ( .A1(n970), .A2(n800), .ZN(n774) );
  XNOR2_X1 U862 ( .A(n774), .B(KEYINPUT81), .ZN(n775) );
  NOR2_X1 U863 ( .A1(G559), .A2(n775), .ZN(n777) );
  NOR2_X1 U864 ( .A1(n982), .A2(G868), .ZN(n776) );
  NOR2_X1 U865 ( .A1(n777), .A2(n776), .ZN(G282) );
  NAND2_X1 U866 ( .A1(G93), .A2(n778), .ZN(n781) );
  NAND2_X1 U867 ( .A1(G67), .A2(n779), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n787) );
  NAND2_X1 U869 ( .A1(G80), .A2(n782), .ZN(n785) );
  NAND2_X1 U870 ( .A1(G55), .A2(n783), .ZN(n784) );
  NAND2_X1 U871 ( .A1(n785), .A2(n784), .ZN(n786) );
  OR2_X1 U872 ( .A1(n787), .A2(n786), .ZN(n801) );
  NAND2_X1 U873 ( .A1(G559), .A2(n893), .ZN(n788) );
  XNOR2_X1 U874 ( .A(n788), .B(KEYINPUT82), .ZN(n798) );
  XNOR2_X1 U875 ( .A(n982), .B(n798), .ZN(n789) );
  NOR2_X1 U876 ( .A1(G860), .A2(n789), .ZN(n790) );
  XOR2_X1 U877 ( .A(n801), .B(n790), .Z(G145) );
  INV_X1 U878 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U879 ( .A(KEYINPUT19), .B(n801), .ZN(n791) );
  XNOR2_X1 U880 ( .A(G288), .B(n791), .ZN(n792) );
  XNOR2_X1 U881 ( .A(n792), .B(G290), .ZN(n793) );
  XNOR2_X1 U882 ( .A(n793), .B(G305), .ZN(n794) );
  XOR2_X1 U883 ( .A(n794), .B(G166), .Z(n796) );
  XNOR2_X1 U884 ( .A(n982), .B(n975), .ZN(n795) );
  XNOR2_X1 U885 ( .A(n796), .B(n795), .ZN(n892) );
  XNOR2_X1 U886 ( .A(KEYINPUT88), .B(n892), .ZN(n797) );
  XNOR2_X1 U887 ( .A(n798), .B(n797), .ZN(n799) );
  NOR2_X1 U888 ( .A1(n800), .A2(n799), .ZN(n803) );
  NOR2_X1 U889 ( .A1(G868), .A2(n801), .ZN(n802) );
  NOR2_X1 U890 ( .A1(n803), .A2(n802), .ZN(G295) );
  NAND2_X1 U891 ( .A1(G2078), .A2(G2084), .ZN(n804) );
  XNOR2_X1 U892 ( .A(n804), .B(KEYINPUT89), .ZN(n805) );
  XNOR2_X1 U893 ( .A(n805), .B(KEYINPUT20), .ZN(n806) );
  NAND2_X1 U894 ( .A1(n806), .A2(G2090), .ZN(n809) );
  XOR2_X1 U895 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n807) );
  XNOR2_X1 U896 ( .A(KEYINPUT21), .B(n807), .ZN(n808) );
  XNOR2_X1 U897 ( .A(n809), .B(n808), .ZN(n810) );
  NAND2_X1 U898 ( .A1(n810), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U899 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U900 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  XNOR2_X1 U901 ( .A(KEYINPUT71), .B(G132), .ZN(G219) );
  NOR2_X1 U902 ( .A1(G220), .A2(G219), .ZN(n812) );
  XNOR2_X1 U903 ( .A(KEYINPUT92), .B(KEYINPUT22), .ZN(n811) );
  XNOR2_X1 U904 ( .A(n812), .B(n811), .ZN(n813) );
  NAND2_X1 U905 ( .A1(n813), .A2(G96), .ZN(n814) );
  NOR2_X1 U906 ( .A1(G218), .A2(n814), .ZN(n815) );
  XNOR2_X1 U907 ( .A(KEYINPUT93), .B(n815), .ZN(n825) );
  NAND2_X1 U908 ( .A1(n825), .A2(G2106), .ZN(n819) );
  NAND2_X1 U909 ( .A1(G69), .A2(G120), .ZN(n816) );
  NOR2_X1 U910 ( .A1(G237), .A2(n816), .ZN(n817) );
  NAND2_X1 U911 ( .A1(G108), .A2(n817), .ZN(n826) );
  NAND2_X1 U912 ( .A1(n826), .A2(G567), .ZN(n818) );
  NAND2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n827) );
  NAND2_X1 U914 ( .A1(G483), .A2(G661), .ZN(n820) );
  NOR2_X1 U915 ( .A1(n827), .A2(n820), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n824), .A2(G36), .ZN(G176) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n821), .ZN(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U919 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U921 ( .A1(n824), .A2(n823), .ZN(G188) );
  XNOR2_X1 U922 ( .A(G96), .B(KEYINPUT109), .ZN(G221) );
  INV_X1 U924 ( .A(G120), .ZN(G236) );
  INV_X1 U925 ( .A(G69), .ZN(G235) );
  NOR2_X1 U926 ( .A1(n826), .A2(n825), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  INV_X1 U928 ( .A(n827), .ZN(G319) );
  XOR2_X1 U929 ( .A(KEYINPUT111), .B(KEYINPUT110), .Z(n829) );
  XNOR2_X1 U930 ( .A(G2678), .B(KEYINPUT43), .ZN(n828) );
  XNOR2_X1 U931 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U932 ( .A(KEYINPUT42), .B(G2090), .Z(n831) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2072), .ZN(n830) );
  XNOR2_X1 U934 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U935 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U936 ( .A(G2096), .B(G2100), .ZN(n834) );
  XNOR2_X1 U937 ( .A(n835), .B(n834), .ZN(n837) );
  XOR2_X1 U938 ( .A(G2078), .B(G2084), .Z(n836) );
  XNOR2_X1 U939 ( .A(n837), .B(n836), .ZN(G227) );
  XOR2_X1 U940 ( .A(G1976), .B(G1971), .Z(n839) );
  XNOR2_X1 U941 ( .A(G1961), .B(G1956), .ZN(n838) );
  XNOR2_X1 U942 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U943 ( .A(n840), .B(KEYINPUT41), .Z(n842) );
  XNOR2_X1 U944 ( .A(G1966), .B(G1981), .ZN(n841) );
  XNOR2_X1 U945 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U946 ( .A(G2474), .B(G1991), .Z(n844) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1996), .ZN(n843) );
  XNOR2_X1 U948 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U949 ( .A(n846), .B(n845), .ZN(G229) );
  NAND2_X1 U950 ( .A1(G124), .A2(n870), .ZN(n847) );
  XNOR2_X1 U951 ( .A(n847), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U952 ( .A1(G100), .A2(n864), .ZN(n848) );
  XNOR2_X1 U953 ( .A(n848), .B(KEYINPUT112), .ZN(n849) );
  NAND2_X1 U954 ( .A1(n850), .A2(n849), .ZN(n854) );
  NAND2_X1 U955 ( .A1(G112), .A2(n871), .ZN(n852) );
  NAND2_X1 U956 ( .A1(G136), .A2(n865), .ZN(n851) );
  NAND2_X1 U957 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U958 ( .A1(n854), .A2(n853), .ZN(G162) );
  NAND2_X1 U959 ( .A1(G103), .A2(n864), .ZN(n856) );
  NAND2_X1 U960 ( .A1(G139), .A2(n865), .ZN(n855) );
  NAND2_X1 U961 ( .A1(n856), .A2(n855), .ZN(n862) );
  NAND2_X1 U962 ( .A1(G127), .A2(n870), .ZN(n858) );
  NAND2_X1 U963 ( .A1(G115), .A2(n871), .ZN(n857) );
  NAND2_X1 U964 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U965 ( .A(KEYINPUT115), .B(n859), .ZN(n860) );
  XNOR2_X1 U966 ( .A(KEYINPUT47), .B(n860), .ZN(n861) );
  NOR2_X1 U967 ( .A1(n862), .A2(n861), .ZN(n917) );
  XOR2_X1 U968 ( .A(G162), .B(n917), .Z(n863) );
  XNOR2_X1 U969 ( .A(n924), .B(n863), .ZN(n878) );
  NAND2_X1 U970 ( .A1(G106), .A2(n864), .ZN(n867) );
  NAND2_X1 U971 ( .A1(G142), .A2(n865), .ZN(n866) );
  NAND2_X1 U972 ( .A1(n867), .A2(n866), .ZN(n869) );
  XOR2_X1 U973 ( .A(KEYINPUT114), .B(KEYINPUT45), .Z(n868) );
  XNOR2_X1 U974 ( .A(n869), .B(n868), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G130), .A2(n870), .ZN(n873) );
  NAND2_X1 U976 ( .A1(G118), .A2(n871), .ZN(n872) );
  NAND2_X1 U977 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U978 ( .A(KEYINPUT113), .B(n874), .Z(n875) );
  NOR2_X1 U979 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U980 ( .A(n878), .B(n877), .Z(n881) );
  XNOR2_X1 U981 ( .A(G160), .B(n879), .ZN(n880) );
  XNOR2_X1 U982 ( .A(n881), .B(n880), .ZN(n886) );
  XOR2_X1 U983 ( .A(KEYINPUT116), .B(KEYINPUT46), .Z(n884) );
  XOR2_X1 U984 ( .A(n882), .B(KEYINPUT48), .Z(n883) );
  XNOR2_X1 U985 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U986 ( .A(n886), .B(n885), .Z(n889) );
  XNOR2_X1 U987 ( .A(G164), .B(n887), .ZN(n888) );
  XNOR2_X1 U988 ( .A(n889), .B(n888), .ZN(n890) );
  NOR2_X1 U989 ( .A1(G37), .A2(n890), .ZN(n891) );
  XOR2_X1 U990 ( .A(KEYINPUT117), .B(n891), .Z(G395) );
  XOR2_X1 U991 ( .A(KEYINPUT118), .B(n892), .Z(n895) );
  XNOR2_X1 U992 ( .A(G171), .B(n893), .ZN(n894) );
  XNOR2_X1 U993 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n896), .B(G286), .ZN(n897) );
  NOR2_X1 U995 ( .A1(G37), .A2(n897), .ZN(G397) );
  XOR2_X1 U996 ( .A(G2438), .B(G2435), .Z(n899) );
  XNOR2_X1 U997 ( .A(G2443), .B(KEYINPUT108), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U999 ( .A(n900), .B(G2454), .Z(n902) );
  XNOR2_X1 U1000 ( .A(G1341), .B(G1348), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n906) );
  XOR2_X1 U1002 ( .A(G2451), .B(G2427), .Z(n904) );
  XNOR2_X1 U1003 ( .A(G2430), .B(G2446), .ZN(n903) );
  XNOR2_X1 U1004 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1005 ( .A(n906), .B(n905), .Z(n907) );
  NAND2_X1 U1006 ( .A1(G14), .A2(n907), .ZN(n913) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n913), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n908) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1010 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1012 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  INV_X1 U1015 ( .A(n913), .ZN(G401) );
  XOR2_X1 U1016 ( .A(G2090), .B(G162), .Z(n914) );
  NOR2_X1 U1017 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1018 ( .A(KEYINPUT51), .B(n916), .Z(n933) );
  XNOR2_X1 U1019 ( .A(KEYINPUT119), .B(KEYINPUT50), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(G2072), .B(n917), .ZN(n919) );
  XNOR2_X1 U1021 ( .A(G164), .B(G2078), .ZN(n918) );
  NAND2_X1 U1022 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1023 ( .A(n921), .B(n920), .ZN(n922) );
  NAND2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n931) );
  XNOR2_X1 U1025 ( .A(G160), .B(G2084), .ZN(n925) );
  NAND2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1032 ( .A(KEYINPUT52), .B(n936), .Z(n937) );
  NOR2_X1 U1033 ( .A1(KEYINPUT55), .A2(n937), .ZN(n938) );
  XOR2_X1 U1034 ( .A(KEYINPUT120), .B(n938), .Z(n939) );
  NAND2_X1 U1035 ( .A1(G29), .A2(n939), .ZN(n1020) );
  XOR2_X1 U1036 ( .A(G2090), .B(G35), .Z(n957) );
  XNOR2_X1 U1037 ( .A(G25), .B(n940), .ZN(n941) );
  NAND2_X1 U1038 ( .A1(n941), .A2(G28), .ZN(n953) );
  XNOR2_X1 U1039 ( .A(KEYINPUT121), .B(G2072), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(n942), .B(G33), .ZN(n951) );
  INV_X1 U1041 ( .A(G1996), .ZN(n943) );
  XNOR2_X1 U1042 ( .A(n943), .B(G32), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(n944), .B(G26), .ZN(n945) );
  NAND2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n949) );
  XOR2_X1 U1045 ( .A(n947), .B(G27), .Z(n948) );
  NOR2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1049 ( .A(KEYINPUT122), .B(n954), .Z(n955) );
  XNOR2_X1 U1050 ( .A(n955), .B(KEYINPUT53), .ZN(n956) );
  NAND2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(G34), .B(G2084), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(KEYINPUT54), .B(n958), .ZN(n959) );
  NOR2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(n961), .B(KEYINPUT55), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(G29), .B(KEYINPUT123), .ZN(n962) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(G11), .A2(n964), .ZN(n1018) );
  XNOR2_X1 U1059 ( .A(G16), .B(KEYINPUT56), .ZN(n988) );
  XNOR2_X1 U1060 ( .A(G168), .B(G1966), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(n967), .B(KEYINPUT57), .ZN(n986) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(G1348), .B(n970), .ZN(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n981) );
  XNOR2_X1 U1066 ( .A(G171), .B(G1961), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(G1971), .A2(G303), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n979) );
  XNOR2_X1 U1069 ( .A(n975), .B(G1956), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n984) );
  XNOR2_X1 U1073 ( .A(G1341), .B(n982), .ZN(n983) );
  NOR2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n1016) );
  INV_X1 U1077 ( .A(G16), .ZN(n1014) );
  XOR2_X1 U1078 ( .A(G20), .B(G1956), .Z(n992) );
  XNOR2_X1 U1079 ( .A(G1341), .B(G19), .ZN(n990) );
  XNOR2_X1 U1080 ( .A(G6), .B(G1981), .ZN(n989) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n995) );
  XOR2_X1 U1083 ( .A(KEYINPUT59), .B(G1348), .Z(n993) );
  XNOR2_X1 U1084 ( .A(G4), .B(n993), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(KEYINPUT124), .B(n996), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(n997), .B(KEYINPUT60), .ZN(n1009) );
  XOR2_X1 U1088 ( .A(G1986), .B(KEYINPUT127), .Z(n998) );
  XNOR2_X1 U1089 ( .A(G24), .B(n998), .ZN(n1004) );
  XOR2_X1 U1090 ( .A(G1971), .B(G22), .Z(n999) );
  XNOR2_X1 U1091 ( .A(KEYINPUT125), .B(n999), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(G23), .B(G1976), .ZN(n1000) );
  NOR2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1094 ( .A(KEYINPUT126), .B(n1002), .Z(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1096 ( .A(KEYINPUT58), .B(n1005), .Z(n1007) );
  XNOR2_X1 U1097 ( .A(G1966), .B(G21), .ZN(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(G5), .B(G1961), .ZN(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1012), .ZN(n1013) );
  NAND2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1021), .Z(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

