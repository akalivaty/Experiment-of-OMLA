//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NAND2_X1  g0005(.A1(G116), .A2(G270), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n207));
  INV_X1    g0007(.A(KEYINPUT66), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(KEYINPUT66), .A2(G68), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n206), .B(new_n207), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(KEYINPUT67), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n214), .A2(KEYINPUT67), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n205), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT1), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT64), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G20), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G58), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(new_n209), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n205), .A2(G13), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n233), .B(G250), .C1(G257), .C2(G264), .ZN(new_n234));
  INV_X1    g0034(.A(KEYINPUT0), .ZN(new_n235));
  AOI22_X1  g0035(.A1(new_n228), .A2(new_n232), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g0036(.A(new_n236), .B1(new_n235), .B2(new_n234), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT65), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n221), .A2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT2), .B(G226), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G250), .B(G257), .Z(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G358));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT68), .ZN(new_n249));
  XOR2_X1   g0049(.A(G50), .B(G58), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G116), .Z(new_n252));
  XNOR2_X1  g0052(.A(G97), .B(G107), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G50), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n227), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n256), .A2(G20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n260), .B1(new_n265), .B2(new_n259), .ZN(new_n266));
  XOR2_X1   g0066(.A(KEYINPUT8), .B(G58), .Z(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n226), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G150), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  OAI22_X1  g0073(.A1(new_n271), .A2(new_n273), .B1(new_n201), .B2(new_n222), .ZN(new_n274));
  OR2_X1    g0074(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n266), .B1(new_n275), .B2(new_n262), .ZN(new_n276));
  OR2_X1    g0076(.A1(new_n276), .A2(KEYINPUT9), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(KEYINPUT9), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT10), .ZN(new_n280));
  INV_X1    g0080(.A(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n287), .A2(G223), .B1(G77), .B2(new_n285), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n285), .A2(G1698), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(KEYINPUT70), .A3(G222), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT70), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT3), .B(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n286), .ZN(new_n293));
  INV_X1    g0093(.A(G222), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n291), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n288), .A2(new_n290), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n227), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G41), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n256), .B(G274), .C1(G41), .C2(G45), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT69), .ZN(new_n303));
  INV_X1    g0103(.A(G41), .ZN(new_n304));
  INV_X1    g0104(.A(G45), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT69), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n306), .A2(new_n307), .A3(new_n256), .A4(G274), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n256), .A2(new_n306), .B1(new_n297), .B2(new_n298), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n310), .B1(G226), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n301), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G190), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n313), .A2(G200), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n279), .A2(new_n280), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n277), .A2(new_n317), .A3(new_n278), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT10), .B1(new_n319), .B2(new_n315), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n289), .A2(G232), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n287), .A2(G238), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n285), .A2(G107), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n300), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n310), .B1(G244), .B2(new_n311), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G169), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G179), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n326), .A2(new_n331), .A3(new_n327), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT64), .B(G20), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n267), .A2(new_n272), .B1(new_n333), .B2(G77), .ZN(new_n334));
  XOR2_X1   g0134(.A(KEYINPUT15), .B(G87), .Z(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n334), .B1(new_n269), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n262), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n262), .B1(new_n256), .B2(G20), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G77), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n338), .B(new_n340), .C1(G77), .C2(new_n257), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n330), .A2(new_n332), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n341), .B1(new_n328), .B2(G200), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n314), .B2(new_n328), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n276), .B1(new_n313), .B2(new_n329), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(G179), .B2(new_n313), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n321), .A2(new_n342), .A3(new_n344), .A4(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n292), .A2(G232), .A3(G1698), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G97), .ZN(new_n349));
  INV_X1    g0149(.A(G226), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n348), .B(new_n349), .C1(new_n293), .C2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n300), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n311), .A2(G238), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n355), .A2(new_n309), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n352), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n354), .B1(new_n352), .B2(new_n356), .ZN(new_n358));
  OAI21_X1  g0158(.A(G200), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n352), .A2(new_n354), .A3(new_n356), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n355), .A2(new_n309), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(new_n300), .B2(new_n351), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT13), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n360), .B(G190), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n269), .A2(new_n202), .ZN(new_n365));
  XOR2_X1   g0165(.A(KEYINPUT66), .B(G68), .Z(new_n366));
  OAI22_X1  g0166(.A1(new_n366), .A2(new_n222), .B1(new_n259), .B2(new_n273), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n262), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT11), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT11), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n370), .B(new_n262), .C1(new_n365), .C2(new_n367), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n212), .A2(new_n258), .A3(KEYINPUT12), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT12), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n257), .B2(G68), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n372), .B(new_n374), .C1(new_n265), .C2(new_n209), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT72), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n339), .A2(G68), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT72), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n377), .A2(new_n372), .A3(new_n378), .A4(new_n374), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n369), .A2(new_n371), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n359), .A2(new_n364), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT73), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n359), .A2(new_n364), .A3(KEYINPUT73), .A4(new_n380), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n380), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n360), .B(G179), .C1(new_n362), .C2(new_n363), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n352), .A2(new_n356), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n353), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n329), .B1(new_n389), .B2(new_n360), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT14), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n387), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n391), .B(G169), .C1(new_n357), .C2(new_n358), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n386), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n385), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n265), .A2(new_n267), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n268), .A2(new_n257), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT74), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT74), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT7), .B1(new_n292), .B2(G20), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n226), .A2(new_n285), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n406), .A3(G68), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n272), .A2(G159), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n210), .A2(G58), .A3(new_n211), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n230), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n408), .B1(new_n410), .B2(G20), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n407), .A2(new_n411), .A3(KEYINPUT16), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n262), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n285), .A2(new_n405), .A3(new_n222), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n223), .A2(new_n225), .B1(new_n282), .B2(new_n284), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n414), .B(new_n366), .C1(new_n415), .C2(new_n405), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT16), .B1(new_n416), .B2(new_n411), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n403), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n282), .A2(new_n284), .A3(G226), .A4(G1698), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n282), .A2(new_n284), .A3(G223), .A4(new_n286), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G87), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n300), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n311), .A2(G232), .B1(new_n303), .B2(new_n308), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n423), .A2(G190), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G200), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(new_n423), .B2(new_n424), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT17), .B1(new_n418), .B2(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n416), .A2(new_n411), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n262), .B(new_n412), .C1(new_n430), .C2(KEYINPUT16), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n425), .A2(new_n427), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT17), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n431), .A2(new_n432), .A3(new_n433), .A4(new_n403), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n423), .A2(new_n331), .A3(new_n424), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(G169), .B1(new_n423), .B2(new_n424), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT75), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT75), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n423), .A2(new_n424), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n440), .B(new_n436), .C1(new_n441), .C2(G169), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n443), .A2(KEYINPUT18), .A3(new_n418), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT18), .B1(new_n443), .B2(new_n418), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n435), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n347), .A2(new_n396), .A3(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n282), .A2(new_n284), .A3(G257), .A4(new_n286), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n282), .A2(new_n284), .A3(G264), .A4(G1698), .ZN(new_n449));
  INV_X1    g0249(.A(G303), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n448), .B(new_n449), .C1(new_n450), .C2(new_n292), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n300), .ZN(new_n452));
  AND2_X1   g0252(.A1(KEYINPUT5), .A2(G41), .ZN(new_n453));
  NOR2_X1   g0253(.A1(KEYINPUT5), .A2(G41), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n256), .A2(G45), .A3(G274), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g0257(.A(KEYINPUT5), .B(G41), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n305), .A2(G1), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n458), .A2(new_n459), .B1(new_n297), .B2(new_n298), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n457), .B1(new_n460), .B2(G270), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n329), .B1(new_n452), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n257), .A2(G116), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n256), .A2(G33), .ZN(new_n464));
  AND4_X1   g0264(.A1(new_n227), .A2(new_n257), .A3(new_n261), .A4(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n463), .B1(new_n465), .B2(G116), .ZN(new_n466));
  INV_X1    g0266(.A(G116), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n261), .A2(new_n227), .B1(G20), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n281), .A2(G97), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G283), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n468), .B(KEYINPUT20), .C1(new_n333), .C2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n224), .A2(G20), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n470), .B(new_n469), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT20), .B1(new_n476), .B2(new_n468), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n466), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT21), .B1(new_n462), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n452), .A2(new_n461), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G200), .ZN(new_n482));
  INV_X1    g0282(.A(new_n478), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n482), .B(new_n483), .C1(new_n314), .C2(new_n481), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n478), .A2(new_n481), .A3(KEYINPUT21), .A4(G169), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n256), .A2(G45), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n299), .B(G270), .C1(new_n455), .C2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n458), .A2(G274), .A3(new_n459), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n489), .B1(new_n300), .B2(new_n451), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(new_n478), .A3(G179), .ZN(new_n491));
  AND4_X1   g0291(.A1(new_n480), .A2(new_n484), .A3(new_n485), .A4(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n298), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n486), .B(G250), .C1(new_n493), .C2(new_n227), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n456), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n282), .A2(new_n284), .A3(G244), .A4(G1698), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n282), .A2(new_n284), .A3(G238), .A4(new_n286), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G116), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AOI211_X1 g0299(.A(G179), .B(new_n495), .C1(new_n499), .C2(new_n300), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n335), .A2(new_n257), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n226), .A2(G33), .A3(G97), .ZN(new_n502));
  AND2_X1   g0302(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n503));
  NOR2_X1   g0303(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n504));
  OR2_X1    g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  OR3_X1    g0306(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n503), .A2(new_n504), .A3(new_n349), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(new_n333), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n226), .A2(new_n292), .A3(G68), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n506), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n501), .B1(new_n511), .B2(new_n262), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n465), .A2(new_n335), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n500), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n495), .B1(new_n499), .B2(new_n300), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n329), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(G200), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n515), .A2(G190), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n465), .A2(G87), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n519), .A2(new_n512), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n299), .B(G257), .C1(new_n455), .C2(new_n486), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n457), .B1(new_n524), .B2(KEYINPUT78), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT78), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n460), .A2(new_n526), .A3(G257), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n282), .A2(new_n284), .A3(G244), .A4(new_n286), .ZN(new_n529));
  NOR2_X1   g0329(.A1(KEYINPUT76), .A2(KEYINPUT4), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n530), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n292), .A2(G244), .A3(new_n286), .A4(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n282), .A2(new_n284), .A3(G250), .A4(G1698), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n531), .A2(new_n533), .A3(new_n470), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n300), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n528), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n329), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT6), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n253), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(G107), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(KEYINPUT6), .A3(G97), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n543), .A2(new_n333), .B1(G77), .B2(new_n272), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n414), .B(G107), .C1(new_n415), .C2(new_n405), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n262), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n257), .A2(G97), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n465), .B2(G97), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT77), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n470), .B(new_n534), .C1(new_n529), .C2(new_n530), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n529), .A2(new_n530), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n551), .B(new_n300), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n551), .B1(new_n535), .B2(new_n300), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n528), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n538), .B(new_n550), .C1(G179), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(G200), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n547), .A2(new_n549), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n528), .A2(KEYINPUT79), .A3(G190), .A4(new_n536), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n536), .A2(G190), .A3(new_n527), .A4(new_n525), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT79), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n559), .A2(new_n560), .A3(new_n561), .A4(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n492), .A2(new_n523), .A3(new_n558), .A4(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n258), .A2(KEYINPUT25), .A3(new_n541), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT25), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n257), .B2(G107), .ZN(new_n569));
  AOI22_X1  g0369(.A1(G107), .A2(new_n465), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT23), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n223), .A2(new_n225), .A3(new_n571), .A4(new_n541), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n498), .A2(new_n571), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n222), .ZN(new_n574));
  NAND2_X1  g0374(.A1(KEYINPUT23), .A2(G107), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n226), .A2(new_n292), .A3(G87), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT22), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT22), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n226), .A2(new_n292), .A3(new_n579), .A4(G87), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n576), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n262), .B1(new_n581), .B2(KEYINPUT24), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT24), .ZN(new_n583));
  AOI211_X1 g0383(.A(new_n583), .B(new_n576), .C1(new_n578), .C2(new_n580), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n570), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n282), .A2(new_n284), .A3(G250), .A4(new_n286), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT81), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n292), .A2(KEYINPUT81), .A3(G250), .A4(new_n286), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G33), .A2(G294), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n292), .A2(G257), .A3(G1698), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n588), .A2(new_n589), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n300), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n460), .A2(G264), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n593), .A2(new_n331), .A3(new_n594), .A4(new_n488), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n488), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n329), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n585), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n578), .A2(new_n580), .ZN(new_n599));
  INV_X1    g0399(.A(new_n576), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n583), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n581), .A2(KEYINPUT24), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n262), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n596), .A2(G200), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n593), .A2(G190), .A3(new_n594), .A4(new_n488), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n570), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n598), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT82), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n598), .A2(new_n607), .A3(KEYINPUT82), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n566), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n447), .A2(new_n612), .ZN(G372));
  AND3_X1   g0413(.A1(new_n512), .A2(new_n520), .A3(new_n521), .ZN(new_n614));
  INV_X1    g0414(.A(new_n495), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n499), .A2(KEYINPUT83), .A3(new_n300), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT83), .B1(new_n499), .B2(new_n300), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G200), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n329), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n614), .A2(new_n619), .B1(new_n514), .B2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n565), .A2(new_n607), .A3(new_n621), .A4(new_n558), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n485), .A2(new_n491), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n623), .A2(new_n479), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT84), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n624), .A2(new_n598), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n625), .B1(new_n624), .B2(new_n598), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n622), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n538), .A2(new_n550), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n557), .A2(G179), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(new_n633), .A3(new_n621), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n518), .A2(new_n522), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT26), .B1(new_n635), .B2(new_n558), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n514), .A2(new_n620), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n629), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n447), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT85), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n342), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n330), .A2(KEYINPUT85), .A3(new_n332), .A4(new_n341), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n385), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT86), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(new_n647), .A3(new_n395), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n383), .A2(new_n384), .B1(new_n643), .B2(new_n644), .ZN(new_n649));
  INV_X1    g0449(.A(new_n387), .ZN(new_n650));
  OAI21_X1  g0450(.A(G169), .B1(new_n357), .B2(new_n358), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n650), .B1(KEYINPUT14), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n380), .B1(new_n652), .B2(new_n393), .ZN(new_n653));
  OAI21_X1  g0453(.A(KEYINPUT86), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n648), .A2(new_n654), .A3(new_n435), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n443), .A2(new_n418), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT18), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n443), .A2(KEYINPUT18), .A3(new_n418), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n655), .A2(KEYINPUT87), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n321), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT87), .B1(new_n655), .B2(new_n660), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n346), .B(new_n641), .C1(new_n662), .C2(new_n663), .ZN(G369));
  INV_X1    g0464(.A(G13), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n333), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n256), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT27), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n666), .A2(new_n669), .A3(new_n256), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n668), .A2(G213), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n598), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n610), .A2(new_n611), .ZN(new_n675));
  INV_X1    g0475(.A(new_n673), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n585), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n674), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n624), .A2(new_n676), .ZN(new_n679));
  XOR2_X1   g0479(.A(new_n679), .B(KEYINPUT88), .Z(new_n680));
  NOR2_X1   g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n676), .A2(new_n478), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n492), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n624), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n678), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n598), .A2(new_n676), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n682), .A2(new_n688), .A3(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n233), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n507), .A2(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n231), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  INV_X1    g0498(.A(new_n537), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n481), .A2(new_n331), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n593), .A2(new_n594), .A3(new_n515), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n699), .A2(KEYINPUT30), .A3(new_n700), .A4(new_n701), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n490), .A2(G179), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n557), .A2(new_n596), .A3(new_n618), .A4(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n676), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(KEYINPUT31), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n710), .B1(new_n612), .B2(new_n673), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT31), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G330), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n523), .A2(new_n632), .A3(new_n633), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n632), .A2(new_n621), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n637), .B(new_n717), .C1(new_n718), .C2(new_n633), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n622), .B1(new_n598), .B2(new_n624), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT29), .B(new_n673), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n676), .B1(new_n629), .B2(new_n639), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(KEYINPUT29), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n716), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n698), .B1(new_n724), .B2(G1), .ZN(G364));
  INV_X1    g0525(.A(new_n686), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT89), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n256), .B1(new_n666), .B2(G45), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n727), .B1(new_n729), .B2(new_n693), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n728), .A2(KEYINPUT89), .A3(new_n694), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n726), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(G330), .B2(new_n685), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n292), .A2(new_n233), .ZN(new_n736));
  INV_X1    g0536(.A(G355), .ZN(new_n737));
  OAI22_X1  g0537(.A1(new_n736), .A2(new_n737), .B1(G116), .B2(new_n233), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n251), .A2(G45), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n692), .A2(new_n292), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(new_n305), .B2(new_n232), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n738), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n227), .B1(G20), .B2(new_n329), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n733), .B1(new_n743), .B2(new_n749), .ZN(new_n750));
  NOR4_X1   g0550(.A1(new_n226), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G159), .ZN(new_n752));
  XOR2_X1   g0552(.A(new_n752), .B(KEYINPUT32), .Z(new_n753));
  NOR2_X1   g0553(.A1(new_n426), .A2(G179), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT90), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n222), .A2(new_n314), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G87), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n755), .A2(new_n314), .A3(new_n333), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G107), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n314), .A2(G179), .A3(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n226), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n285), .B1(new_n765), .B2(G97), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n753), .A2(new_n759), .A3(new_n762), .A4(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n226), .A2(new_n331), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G190), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n426), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(G200), .ZN(new_n771));
  AOI22_X1  g0571(.A1(G50), .A2(new_n770), .B1(new_n771), .B2(G58), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n768), .A2(new_n314), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n426), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n773), .A2(G200), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n772), .B1(new_n209), .B2(new_n775), .C1(new_n202), .C2(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(G322), .A2(new_n771), .B1(new_n770), .B2(G326), .ZN(new_n779));
  INV_X1    g0579(.A(G311), .ZN(new_n780));
  XNOR2_X1  g0580(.A(KEYINPUT91), .B(KEYINPUT33), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(G317), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n779), .B1(new_n780), .B2(new_n777), .C1(new_n775), .C2(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n761), .A2(G283), .B1(G329), .B2(new_n751), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n292), .B1(new_n765), .B2(G294), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n784), .B(new_n785), .C1(new_n450), .C2(new_n757), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n767), .A2(new_n778), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n787), .A2(KEYINPUT92), .ZN(new_n788));
  INV_X1    g0588(.A(new_n747), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(new_n787), .B2(KEYINPUT92), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n750), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n746), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n791), .B1(new_n685), .B2(new_n792), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n735), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(G396));
  NOR2_X1   g0595(.A1(new_n747), .A2(new_n744), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n733), .B1(G77), .B2(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G143), .A2(new_n771), .B1(new_n776), .B2(G159), .ZN(new_n799));
  INV_X1    g0599(.A(G137), .ZN(new_n800));
  INV_X1    g0600(.A(new_n770), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n799), .B1(new_n800), .B2(new_n801), .C1(new_n271), .C2(new_n775), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT94), .Z(new_n803));
  OR2_X1    g0603(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n760), .A2(new_n209), .ZN(new_n806));
  INV_X1    g0606(.A(new_n751), .ZN(new_n807));
  INV_X1    g0607(.A(G132), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n292), .B1(new_n229), .B2(new_n764), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n806), .B(new_n809), .C1(G50), .C2(new_n758), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n804), .A2(new_n805), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n761), .A2(G87), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n780), .B2(new_n807), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT93), .ZN(new_n814));
  INV_X1    g0614(.A(G97), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n285), .B1(new_n815), .B2(new_n764), .C1(new_n757), .C2(new_n541), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(G294), .B2(new_n771), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n776), .A2(G116), .ZN(new_n818));
  AOI22_X1  g0618(.A1(G283), .A2(new_n774), .B1(new_n770), .B2(G303), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n814), .A2(new_n817), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n789), .B1(new_n811), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n676), .A2(new_n341), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n344), .A2(new_n342), .A3(new_n822), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n643), .A2(new_n644), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n824), .B2(new_n822), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n798), .B(new_n821), .C1(new_n744), .C2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n716), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n722), .B(new_n826), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n733), .B1(new_n828), .B2(new_n829), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n827), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G384));
  OAI211_X1 g0634(.A(G116), .B(new_n228), .C1(new_n543), .C2(KEYINPUT35), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(KEYINPUT35), .B2(new_n543), .ZN(new_n836));
  XOR2_X1   g0636(.A(KEYINPUT95), .B(KEYINPUT36), .Z(new_n837));
  NAND3_X1  g0637(.A1(new_n232), .A2(G77), .A3(new_n409), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT96), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n838), .A2(new_n839), .B1(new_n259), .B2(G68), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n256), .A2(G13), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n836), .A2(new_n837), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n380), .A2(new_n673), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT97), .ZN(new_n845));
  AND3_X1   g0645(.A1(new_n385), .A2(new_n395), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n845), .B1(new_n385), .B2(new_n395), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n848), .A2(new_n826), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n715), .B(new_n849), .C1(KEYINPUT101), .C2(KEYINPUT40), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT16), .B1(new_n407), .B2(new_n411), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n399), .B1(new_n413), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n672), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n431), .A2(new_n432), .A3(new_n403), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n407), .A2(new_n411), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT16), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n858), .A2(new_n262), .A3(new_n412), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n439), .A2(new_n442), .B1(new_n859), .B2(new_n399), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT37), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n418), .A2(new_n672), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n656), .A2(new_n862), .A3(new_n854), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT98), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n861), .A2(new_n864), .A3(KEYINPUT98), .ZN(new_n868));
  INV_X1    g0668(.A(new_n853), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n446), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n867), .A2(KEYINPUT38), .A3(new_n868), .A4(new_n870), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AND4_X1   g0675(.A1(new_n558), .A2(new_n492), .A3(new_n523), .A4(new_n565), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(new_n675), .A3(new_n673), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n714), .B1(new_n877), .B2(new_n709), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n878), .A2(new_n711), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n879), .A2(new_n826), .A3(new_n848), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n850), .B(new_n875), .C1(new_n880), .C2(KEYINPUT101), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT99), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n435), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n429), .A2(KEYINPUT99), .A3(new_n434), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n660), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n863), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n656), .A2(new_n854), .A3(new_n863), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n885), .A2(new_n886), .B1(new_n864), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n889), .A2(KEYINPUT38), .ZN(new_n890));
  INV_X1    g0690(.A(new_n874), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT40), .B1(new_n850), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n881), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n447), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n895), .A2(new_n879), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(G330), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n881), .B2(new_n893), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n716), .A2(new_n895), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n395), .A2(new_n676), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n865), .A2(new_n866), .B1(new_n446), .B2(new_n869), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n904), .B2(new_n868), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT39), .B1(new_n891), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n874), .B(new_n907), .C1(new_n889), .C2(KEYINPUT38), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n903), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n673), .B(new_n825), .C1(new_n628), .C2(new_n638), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n342), .A2(new_n676), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n848), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n875), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n660), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n671), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT100), .B1(new_n909), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n908), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n907), .B1(new_n873), .B2(new_n874), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n902), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT100), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n875), .A2(new_n913), .B1(new_n915), .B2(new_n671), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n918), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n901), .B(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n447), .B(new_n721), .C1(new_n722), .C2(KEYINPUT29), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n928), .B(new_n346), .C1(new_n662), .C2(new_n663), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n927), .A2(new_n929), .B1(new_n256), .B2(new_n666), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n927), .A2(new_n929), .ZN(new_n931));
  OAI221_X1 g0731(.A(new_n843), .B1(new_n836), .B2(new_n837), .C1(new_n930), .C2(new_n931), .ZN(G367));
  OAI211_X1 g0732(.A(new_n565), .B(new_n558), .C1(new_n560), .C2(new_n673), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n558), .B2(new_n673), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT103), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n682), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT42), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n558), .B1(new_n935), .B2(new_n598), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n673), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n512), .A2(new_n521), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n676), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n621), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n637), .B2(new_n942), .ZN(new_n944));
  XOR2_X1   g0744(.A(KEYINPUT102), .B(KEYINPUT43), .Z(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(KEYINPUT43), .B2(new_n944), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n940), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n937), .A2(new_n939), .A3(new_n946), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n688), .A2(new_n935), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n950), .B(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n693), .B(KEYINPUT41), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  OR3_X1    g0754(.A1(new_n681), .A2(KEYINPUT106), .A3(new_n726), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n678), .A2(new_n680), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n726), .B1(new_n681), .B2(KEYINPUT106), .ZN(new_n957));
  AND3_X1   g0757(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n956), .B1(new_n955), .B2(new_n957), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n724), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n960), .A2(KEYINPUT107), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(KEYINPUT107), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT105), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n934), .B(KEYINPUT103), .Z(new_n964));
  NAND3_X1  g0764(.A1(new_n964), .A2(new_n682), .A3(new_n690), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(KEYINPUT45), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n935), .B1(new_n681), .B2(new_n689), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT44), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n968), .A2(KEYINPUT104), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n966), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n965), .A2(KEYINPUT45), .B1(new_n967), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n963), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n688), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n963), .B(new_n687), .C1(new_n971), .C2(new_n974), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n961), .A2(new_n962), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n954), .B1(new_n978), .B2(new_n724), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n952), .B1(new_n979), .B2(new_n729), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n246), .A2(new_n741), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n748), .B1(new_n233), .B2(new_n336), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n733), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n760), .A2(new_n202), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n765), .A2(G68), .ZN(new_n986));
  AND3_X1   g0786(.A1(new_n985), .A2(new_n292), .A3(new_n986), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n758), .A2(G58), .B1(G137), .B2(new_n751), .ZN(new_n988));
  AOI22_X1  g0788(.A1(G50), .A2(new_n776), .B1(new_n771), .B2(G150), .ZN(new_n989));
  AOI22_X1  g0789(.A1(G143), .A2(new_n770), .B1(new_n774), .B2(G159), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n760), .A2(new_n815), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n292), .B(new_n992), .C1(G317), .C2(new_n751), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n758), .A2(G116), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT46), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n771), .A2(G303), .ZN(new_n996));
  AOI22_X1  g0796(.A1(G294), .A2(new_n774), .B1(new_n770), .B2(G311), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n993), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n776), .A2(G283), .B1(G107), .B2(new_n765), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT108), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n991), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT47), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n789), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n983), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n792), .B2(new_n944), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n980), .A2(new_n1006), .ZN(G387));
  NAND2_X1  g0807(.A1(new_n961), .A2(new_n962), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n958), .A2(new_n959), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n724), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1011), .A2(KEYINPUT110), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(KEYINPUT110), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1008), .A2(new_n1012), .A3(new_n693), .A4(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1009), .A2(new_n728), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n243), .A2(G45), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n1016), .A2(new_n741), .B1(new_n695), .B2(new_n736), .ZN(new_n1017));
  OR3_X1    g0817(.A1(new_n268), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1018));
  OAI21_X1  g0818(.A(KEYINPUT50), .B1(new_n268), .B2(G50), .ZN(new_n1019));
  AOI21_X1  g0819(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1018), .A2(new_n695), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1017), .A2(new_n1021), .B1(new_n541), .B2(new_n692), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n758), .A2(G77), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n271), .B2(new_n807), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1025), .A2(KEYINPUT109), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1025), .A2(KEYINPUT109), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G50), .A2(new_n771), .B1(new_n770), .B2(G159), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n268), .B2(new_n775), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n992), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n776), .A2(G68), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n765), .A2(new_n335), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n292), .A4(new_n1032), .ZN(new_n1033));
  NOR4_X1   g0833(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .A4(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G303), .A2(new_n776), .B1(new_n771), .B2(G317), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G311), .A2(new_n774), .B1(new_n770), .B2(G322), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT48), .Z(new_n1038));
  INV_X1    g0838(.A(G294), .ZN(new_n1039));
  INV_X1    g0839(.A(G283), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n757), .A2(new_n1039), .B1(new_n1040), .B2(new_n764), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1042), .A2(KEYINPUT49), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n292), .B1(new_n751), .B2(G326), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n467), .B2(new_n760), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1042), .A2(KEYINPUT49), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1034), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n733), .B1(new_n749), .B2(new_n1022), .C1(new_n1048), .C2(new_n789), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n678), .B2(new_n746), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1015), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1014), .A2(new_n1051), .ZN(G393));
  OAI221_X1 g0852(.A(new_n748), .B1(new_n815), .B2(new_n233), .C1(new_n254), .C2(new_n741), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT112), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n733), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT113), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n777), .A2(new_n1039), .B1(new_n467), .B2(new_n764), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G311), .A2(new_n771), .B1(new_n770), .B2(G317), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT52), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1057), .B(new_n1059), .C1(G303), .C2(new_n774), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n758), .A2(G283), .B1(G322), .B2(new_n751), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1061), .A2(new_n285), .A3(new_n762), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT114), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G150), .A2(new_n770), .B1(new_n771), .B2(G159), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT51), .Z(new_n1065));
  AOI22_X1  g0865(.A1(G50), .A2(new_n774), .B1(new_n776), .B2(new_n267), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n285), .B1(new_n765), .B2(G77), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n758), .A2(new_n366), .B1(G143), .B2(new_n751), .ZN(new_n1068));
  AND4_X1   g0868(.A1(new_n812), .A2(new_n1066), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1060), .A2(new_n1063), .B1(new_n1065), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1056), .B1(new_n1070), .B2(new_n789), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n935), .B2(new_n746), .ZN(new_n1072));
  OR3_X1    g0872(.A1(new_n971), .A2(new_n974), .A3(new_n687), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n687), .B1(new_n971), .B2(new_n974), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n1075), .A2(KEYINPUT111), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n728), .B1(new_n1075), .B2(KEYINPUT111), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1072), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1008), .A2(new_n1075), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1079), .A2(new_n693), .A3(new_n978), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1080), .ZN(G390));
  INV_X1    g0881(.A(new_n848), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n715), .A2(G330), .A3(new_n825), .A4(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n906), .A2(new_n908), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n913), .A2(new_n902), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n673), .B(new_n825), .C1(new_n719), .C2(new_n720), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n848), .B1(new_n1088), .B2(new_n912), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n892), .A2(new_n1089), .A3(new_n902), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1084), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n903), .B1(new_n890), .B2(new_n891), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1083), .B1(new_n1089), .B2(new_n1092), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n929), .A2(new_n900), .ZN(new_n1096));
  OAI211_X1 g0896(.A(G330), .B(new_n825), .C1(new_n878), .C2(new_n711), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n848), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1088), .A2(new_n912), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1083), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1083), .A2(new_n1098), .B1(new_n910), .B2(new_n912), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1096), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n694), .B1(new_n1095), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n1095), .B2(new_n1103), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1095), .A2(new_n729), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n733), .B1(new_n267), .B2(new_n797), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n757), .A2(new_n271), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT53), .ZN(new_n1109));
  XOR2_X1   g0909(.A(KEYINPUT54), .B(G143), .Z(new_n1110));
  AOI22_X1  g0910(.A1(G137), .A2(new_n774), .B1(new_n776), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n285), .B1(new_n765), .B2(G159), .ZN(new_n1113));
  INV_X1    g0913(.A(G125), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1113), .B1(new_n807), .B2(new_n1114), .C1(new_n259), .C2(new_n760), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n770), .A2(G128), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n771), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1116), .B1(new_n1117), .B2(new_n808), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n1112), .A2(new_n1115), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n759), .A2(new_n285), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n806), .B(new_n1120), .C1(G294), .C2(new_n751), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n771), .A2(G116), .B1(G77), .B2(new_n765), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT115), .Z(new_n1123));
  NAND2_X1  g0923(.A1(new_n776), .A2(G97), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G107), .A2(new_n774), .B1(new_n770), .B2(G283), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1121), .A2(new_n1123), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1119), .B1(new_n1126), .B2(KEYINPUT116), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(KEYINPUT116), .B2(new_n1126), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1107), .B1(new_n1128), .B2(new_n747), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT117), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n1085), .B2(new_n745), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1105), .A2(new_n1106), .A3(new_n1131), .ZN(G378));
  INV_X1    g0932(.A(new_n899), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n321), .A2(new_n346), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n276), .A2(new_n671), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1134), .B(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1136), .B(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n918), .A2(new_n924), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1139), .B1(new_n918), .B2(new_n924), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1133), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NOR3_X1   g0942(.A1(new_n909), .A2(new_n917), .A3(KEYINPUT100), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n922), .B1(new_n921), .B2(new_n923), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1138), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n918), .A2(new_n924), .A3(new_n1139), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1145), .A2(new_n899), .A3(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1142), .A2(new_n729), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n732), .B1(new_n259), .B2(new_n796), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G116), .A2(new_n770), .B1(new_n776), .B2(new_n335), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n815), .B2(new_n775), .ZN(new_n1151));
  AND4_X1   g0951(.A1(new_n304), .A2(new_n1023), .A3(new_n285), .A4(new_n986), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n761), .A2(G58), .B1(G283), .B2(new_n751), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n771), .A2(G107), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1152), .B(new_n1153), .C1(KEYINPUT118), .C2(new_n1154), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1151), .B(new_n1155), .C1(KEYINPUT118), .C2(new_n1154), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT58), .Z(new_n1157));
  AOI21_X1  g0957(.A(G50), .B1(new_n281), .B2(new_n304), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n292), .B2(G41), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n758), .A2(new_n1110), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n1114), .A2(new_n801), .B1(new_n1160), .B2(KEYINPUT119), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1160), .A2(KEYINPUT119), .B1(G128), .B2(new_n771), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1162), .B1(new_n800), .B2(new_n777), .C1(new_n271), .C2(new_n764), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1161), .B(new_n1163), .C1(G132), .C2(new_n774), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(KEYINPUT59), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n761), .A2(G159), .ZN(new_n1167));
  AOI211_X1 g0967(.A(G33), .B(G41), .C1(new_n751), .C2(G124), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1165), .A2(KEYINPUT59), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1157), .B(new_n1159), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT120), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n747), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1149), .B1(new_n1174), .B2(new_n1175), .C1(new_n745), .C2(new_n1139), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n1148), .A2(KEYINPUT121), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(KEYINPUT121), .B1(new_n1148), .B2(new_n1176), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1096), .B1(new_n1094), .B2(new_n1102), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1142), .A2(new_n1180), .A3(new_n1147), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT57), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1142), .A2(new_n1180), .A3(new_n1147), .A4(KEYINPUT57), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1183), .A2(new_n693), .A3(new_n1184), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1179), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(G375));
  OR2_X1    g0987(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1188), .A2(new_n1096), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1189), .A2(new_n954), .A3(new_n1103), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT122), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n758), .A2(G97), .B1(G303), .B2(new_n751), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1192), .A2(new_n985), .A3(new_n285), .A4(new_n1032), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(G283), .A2(new_n771), .B1(new_n770), .B2(G294), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1194), .B1(new_n541), .B2(new_n777), .C1(new_n467), .C2(new_n775), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G137), .A2(new_n771), .B1(new_n774), .B2(new_n1110), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1196), .B1(new_n808), .B2(new_n801), .C1(new_n271), .C2(new_n777), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n758), .A2(G159), .B1(G128), .B2(new_n751), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n285), .B1(new_n765), .B2(G50), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(new_n229), .C2(new_n760), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n1193), .A2(new_n1195), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n747), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1202), .B(new_n733), .C1(G68), .C2(new_n797), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n848), .B2(new_n744), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n1188), .B2(new_n729), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1191), .A2(new_n1205), .ZN(G381));
  INV_X1    g1006(.A(G378), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1186), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(G390), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(G393), .A2(G396), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1209), .A2(new_n833), .A3(new_n1210), .ZN(new_n1211));
  OR4_X1    g1011(.A1(G387), .A2(new_n1208), .A3(G381), .A4(new_n1211), .ZN(G407));
  OAI211_X1 g1012(.A(G407), .B(G213), .C1(G343), .C2(new_n1208), .ZN(G409));
  AOI21_X1  g1013(.A(G390), .B1(new_n980), .B2(new_n1006), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n794), .B1(new_n1014), .B2(new_n1051), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1210), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(G390), .A2(new_n980), .A3(new_n1006), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1215), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1218), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n1220), .A2(new_n1214), .B1(new_n1210), .B2(new_n1216), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT61), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1219), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1185), .B(G378), .C1(new_n1178), .C2(new_n1177), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1148), .B(new_n1176), .C1(new_n1181), .C2(new_n954), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1207), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(G343), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1224), .A2(new_n1226), .B1(G213), .B2(new_n1227), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1189), .A2(KEYINPUT60), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1189), .A2(KEYINPUT60), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1229), .A2(new_n693), .A3(new_n1102), .A4(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1231), .A2(G384), .A3(new_n1205), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(G384), .B1(new_n1231), .B2(new_n1205), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1228), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1223), .B1(KEYINPUT63), .B2(new_n1236), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1227), .A2(G213), .A3(G2897), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1238), .B(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT123), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1227), .A2(G213), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT123), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1224), .A2(new_n1226), .A3(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1240), .A2(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1238), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1237), .B(new_n1247), .C1(new_n1248), .C2(new_n1249), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1235), .B(new_n1239), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1222), .B1(new_n1251), .B2(new_n1228), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1241), .A2(KEYINPUT62), .A3(new_n1235), .A4(new_n1243), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(KEYINPUT125), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT125), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1228), .A2(new_n1255), .A3(KEYINPUT62), .A4(new_n1235), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT62), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n1246), .B2(new_n1238), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1252), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1250), .B1(new_n1260), .B2(new_n1261), .ZN(G405));
  NAND2_X1  g1062(.A1(new_n1235), .A2(KEYINPUT126), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1219), .A2(new_n1221), .A3(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1263), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(G375), .A2(G378), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1267), .B(new_n1208), .C1(KEYINPUT126), .C2(new_n1235), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1266), .B(new_n1268), .ZN(G402));
endmodule


