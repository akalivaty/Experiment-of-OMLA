//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n857, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986;
  INV_X1    g000(.A(KEYINPUT41), .ZN(new_n202));
  INV_X1    g001(.A(G232gat), .ZN(new_n203));
  INV_X1    g002(.A(G233gat), .ZN(new_n204));
  NOR3_X1   g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(KEYINPUT97), .B(G92gat), .Z(new_n206));
  INV_X1    g005(.A(G85gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n206), .A2(new_n207), .B1(KEYINPUT8), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT7), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G99gat), .B(G106gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(KEYINPUT98), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT99), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT98), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n213), .B(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(new_n209), .A3(new_n211), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n215), .A2(new_n216), .A3(new_n219), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n218), .A2(KEYINPUT99), .A3(new_n209), .A4(new_n211), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g021(.A(G43gat), .B(G50gat), .Z(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT15), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT15), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT14), .ZN(new_n228));
  INV_X1    g027(.A(G29gat), .ZN(new_n229));
  INV_X1    g028(.A(G36gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n231), .A2(new_n232), .B1(G29gat), .B2(G36gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n225), .A2(new_n227), .A3(new_n233), .ZN(new_n234));
  NOR3_X1   g033(.A1(new_n233), .A2(new_n226), .A3(new_n223), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n205), .B1(new_n222), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G190gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT17), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n234), .A2(new_n236), .A3(KEYINPUT17), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n241), .A2(new_n220), .A3(new_n221), .A4(new_n242), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n238), .A2(new_n239), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n239), .B1(new_n238), .B2(new_n243), .ZN(new_n245));
  INV_X1    g044(.A(G218gat), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n222), .A2(new_n237), .ZN(new_n248));
  INV_X1    g047(.A(new_n205), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n243), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G190gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n238), .A2(new_n239), .A3(new_n243), .ZN(new_n252));
  AOI21_X1  g051(.A(G218gat), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT100), .B1(new_n247), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n246), .B1(new_n244), .B2(new_n245), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n251), .A2(G218gat), .A3(new_n252), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT100), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G134gat), .B(G162gat), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n254), .A2(new_n258), .A3(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n255), .A2(new_n256), .A3(new_n257), .A4(new_n261), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G231gat), .A2(G233gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT19), .ZN(new_n267));
  XOR2_X1   g066(.A(KEYINPUT96), .B(G183gat), .Z(new_n268));
  XOR2_X1   g067(.A(new_n267), .B(new_n268), .Z(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G57gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(KEYINPUT95), .ZN(new_n272));
  INV_X1    g071(.A(G64gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  AND2_X1   g073(.A1(G71gat), .A2(G78gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(G71gat), .A2(G78gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n275), .A2(KEYINPUT9), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n281), .B1(new_n271), .B2(new_n273), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n274), .A2(new_n279), .B1(new_n282), .B2(new_n277), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(KEYINPUT21), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(G15gat), .B(G22gat), .Z(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G1gat), .ZN(new_n287));
  INV_X1    g086(.A(G8gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT90), .ZN(new_n289));
  XNOR2_X1  g088(.A(G15gat), .B(G22gat), .ZN(new_n290));
  INV_X1    g089(.A(G1gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(KEYINPUT16), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n287), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n288), .A2(KEYINPUT90), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n294), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n287), .A2(new_n292), .A3(new_n296), .A4(new_n289), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(KEYINPUT92), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT92), .B1(new_n295), .B2(new_n297), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G211gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n283), .A2(KEYINPUT21), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n302), .B1(new_n301), .B2(new_n303), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n285), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n301), .A2(new_n303), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G211gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n309), .A2(new_n284), .A3(new_n304), .ZN(new_n310));
  XNOR2_X1  g109(.A(G127gat), .B(G155gat), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n311), .B(KEYINPUT20), .Z(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n307), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n313), .B1(new_n307), .B2(new_n310), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n270), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n316), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n318), .A2(new_n269), .A3(new_n314), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n265), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT101), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT101), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n265), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G197gat), .B(G204gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT22), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n327), .B1(new_n302), .B2(new_n246), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  XOR2_X1   g128(.A(G211gat), .B(G218gat), .Z(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT3), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT78), .B(G162gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G155gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT2), .ZN(new_n337));
  XNOR2_X1  g136(.A(G155gat), .B(G162gat), .ZN(new_n338));
  INV_X1    g137(.A(G148gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(G141gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(KEYINPUT77), .B(G141gat), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n340), .B1(new_n341), .B2(new_n339), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n337), .A2(new_n338), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n344));
  INV_X1    g143(.A(G141gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G148gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n340), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT2), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT74), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(KEYINPUT74), .A2(G155gat), .A3(G162gat), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n347), .A2(new_n349), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n354));
  INV_X1    g153(.A(G155gat), .ZN(new_n355));
  INV_X1    g154(.A(G162gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n344), .B1(new_n353), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n345), .A2(G148gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n339), .A2(G141gat), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n349), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n351), .A2(new_n352), .ZN(new_n364));
  AND4_X1   g163(.A1(new_n344), .A2(new_n363), .A3(new_n359), .A4(new_n364), .ZN(new_n365));
  OAI211_X1 g164(.A(KEYINPUT79), .B(new_n343), .C1(new_n360), .C2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n349), .ZN(new_n368));
  XNOR2_X1  g167(.A(G141gat), .B(G148gat), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n359), .B(new_n364), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT76), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n353), .A2(new_n344), .A3(new_n359), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT79), .B1(new_n373), .B2(new_n343), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n334), .B1(new_n367), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G228gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(new_n204), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT3), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n378), .B(new_n343), .C1(new_n360), .C2(new_n365), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n332), .ZN(new_n380));
  INV_X1    g179(.A(new_n331), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n375), .A2(new_n377), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n331), .B1(new_n379), .B2(new_n332), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n345), .A2(KEYINPUT77), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n345), .A2(KEYINPUT77), .ZN(new_n386));
  OAI21_X1  g185(.A(G148gat), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n340), .A2(new_n387), .B1(new_n336), .B2(KEYINPUT2), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n371), .A2(new_n372), .B1(new_n388), .B2(new_n338), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n389), .A2(new_n333), .ZN(new_n390));
  OAI22_X1  g189(.A1(new_n384), .A2(new_n390), .B1(new_n376), .B2(new_n204), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n383), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(G22gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT85), .ZN(new_n394));
  XNOR2_X1  g193(.A(G78gat), .B(G106gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(KEYINPUT31), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(G50gat), .ZN(new_n397));
  INV_X1    g196(.A(G22gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n398), .A3(new_n391), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT86), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n394), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT84), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n399), .A2(KEYINPUT83), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n393), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n392), .A2(KEYINPUT83), .A3(G22gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(new_n397), .B(KEYINPUT82), .Z(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n402), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  AOI211_X1 g208(.A(KEYINPUT84), .B(new_n407), .C1(new_n404), .C2(new_n405), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n401), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(G120gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(G113gat), .ZN(new_n413));
  INV_X1    g212(.A(G113gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(G120gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G127gat), .B(G134gat), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT1), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT68), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n418), .A2(new_n416), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G134gat), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n422), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT69), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n416), .A2(new_n418), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n422), .A2(G127gat), .ZN(new_n426));
  INV_X1    g225(.A(G127gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(G134gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n428), .A3(new_n420), .ZN(new_n429));
  AND4_X1   g228(.A1(KEYINPUT69), .A2(new_n425), .A3(new_n423), .A4(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n419), .B1(new_n424), .B2(new_n430), .ZN(new_n431));
  AND2_X1   g230(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n432));
  NOR2_X1   g231(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n239), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT66), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n435), .A2(KEYINPUT28), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(KEYINPUT28), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n434), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT67), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n440), .A2(G169gat), .A3(G176gat), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n441), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT26), .ZN(new_n443));
  NAND2_X1  g242(.A1(G169gat), .A2(G176gat), .ZN(new_n444));
  INV_X1    g243(.A(G169gat), .ZN(new_n445));
  INV_X1    g244(.A(G176gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n443), .B(new_n444), .C1(new_n447), .C2(new_n440), .ZN(new_n448));
  XNOR2_X1  g247(.A(KEYINPUT27), .B(G183gat), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n449), .A2(new_n239), .A3(new_n436), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n439), .A2(new_n442), .A3(new_n448), .A4(new_n450), .ZN(new_n451));
  OR2_X1    g250(.A1(G183gat), .A2(G190gat), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT24), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT65), .ZN(new_n454));
  NAND2_X1  g253(.A1(G183gat), .A2(G190gat), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n452), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n444), .A2(KEYINPUT23), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n447), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n445), .A2(new_n446), .A3(KEYINPUT23), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n460), .B1(new_n455), .B2(new_n454), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT25), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT64), .ZN(new_n463));
  OR2_X1    g262(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT25), .B1(new_n457), .B2(new_n447), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n455), .A2(new_n453), .ZN(new_n466));
  NAND3_X1  g265(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n452), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n460), .A2(new_n463), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n464), .A2(new_n465), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n451), .A2(new_n462), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT70), .B1(new_n431), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n419), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n425), .A2(new_n423), .A3(new_n429), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT69), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n421), .A2(KEYINPUT69), .A3(new_n423), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n451), .A2(new_n462), .A3(new_n470), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT70), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n431), .A2(new_n471), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n472), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  AND2_X1   g282(.A1(G227gat), .A2(G233gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT32), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT71), .ZN(new_n487));
  XNOR2_X1  g286(.A(G15gat), .B(G43gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(G71gat), .ZN(new_n489));
  INV_X1    g288(.A(G99gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT33), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n492), .B1(new_n485), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT32), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(new_n483), .B2(new_n484), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT71), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n487), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT72), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT72), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n487), .A2(new_n501), .A3(new_n494), .A4(new_n498), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n486), .B1(KEYINPUT33), .B2(new_n491), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n483), .A2(new_n484), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT34), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n503), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n496), .A2(new_n497), .ZN(new_n510));
  AOI211_X1 g309(.A(KEYINPUT71), .B(new_n495), .C1(new_n483), .C2(new_n484), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n501), .B1(new_n512), .B2(new_n494), .ZN(new_n513));
  INV_X1    g312(.A(new_n502), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n505), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n507), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n411), .A2(new_n509), .A3(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(G1gat), .B(G29gat), .Z(new_n518));
  XNOR2_X1  g317(.A(G57gat), .B(G85gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT3), .B1(new_n367), .B2(new_n374), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n379), .A2(new_n431), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n389), .A2(new_n478), .A3(KEYINPUT4), .ZN(new_n528));
  AOI21_X1  g327(.A(KEYINPUT4), .B1(new_n389), .B2(new_n478), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G225gat), .A2(G233gat), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT4), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n527), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n373), .A2(new_n343), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT79), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n478), .B1(new_n537), .B2(new_n366), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n535), .A2(new_n431), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n532), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n534), .A2(KEYINPUT5), .A3(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n532), .A2(KEYINPUT5), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n527), .A2(new_n530), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n523), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT6), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT81), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n544), .A2(KEYINPUT81), .A3(KEYINPUT6), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n541), .A2(new_n543), .A3(new_n523), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT6), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n547), .B(new_n548), .C1(new_n544), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G226gat), .A2(G233gat), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(new_n479), .B2(KEYINPUT29), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n471), .A2(G226gat), .A3(G233gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(new_n381), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n554), .A2(new_n331), .A3(new_n555), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G8gat), .B(G36gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(G92gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT73), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(G64gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT30), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n567), .B1(new_n559), .B2(new_n564), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n560), .A2(new_n567), .A3(new_n565), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n552), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT35), .B1(new_n517), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT89), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n541), .A2(new_n543), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n522), .B(KEYINPUT87), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n578), .A2(new_n550), .A3(new_n549), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n547), .A2(new_n579), .A3(new_n548), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT35), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(new_n581), .A3(new_n571), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n574), .B1(new_n517), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n571), .A2(new_n581), .ZN(new_n584));
  INV_X1    g383(.A(new_n548), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT81), .B1(new_n544), .B2(KEYINPUT6), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n584), .B1(new_n587), .B2(new_n579), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n508), .B1(new_n503), .B2(new_n505), .ZN(new_n589));
  AOI211_X1 g388(.A(new_n504), .B(new_n507), .C1(new_n500), .C2(new_n502), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n588), .A2(new_n591), .A3(KEYINPUT89), .A4(new_n411), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n573), .A2(new_n583), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n411), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n572), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n378), .B1(new_n537), .B2(new_n366), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n596), .A2(new_n525), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT4), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n598), .B1(new_n535), .B2(new_n431), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n389), .A2(new_n478), .A3(KEYINPUT4), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n532), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  OR3_X1    g401(.A1(new_n538), .A2(new_n532), .A3(new_n539), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(KEYINPUT39), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n531), .B1(new_n527), .B2(new_n530), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT39), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n577), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT40), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n608), .A2(KEYINPUT88), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n608), .A2(KEYINPUT88), .B1(new_n575), .B2(new_n577), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n604), .A2(new_n607), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT40), .ZN(new_n612));
  INV_X1    g411(.A(new_n571), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n609), .A2(new_n610), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n559), .B(KEYINPUT37), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n615), .A2(new_n565), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT38), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n547), .A2(new_n618), .A3(new_n579), .A4(new_n548), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n566), .B1(new_n616), .B2(new_n617), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n614), .B(new_n411), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n516), .A2(KEYINPUT36), .A3(new_n509), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT36), .B1(new_n516), .B2(new_n509), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n595), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n325), .B1(new_n593), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n237), .B1(new_n299), .B2(new_n300), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n295), .A2(new_n297), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n241), .A2(new_n627), .A3(new_n242), .ZN(new_n628));
  NAND2_X1  g427(.A1(G229gat), .A2(G233gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT91), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n626), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(KEYINPUT93), .A2(KEYINPUT18), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n630), .B(KEYINPUT13), .Z(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n237), .ZN(new_n637));
  INV_X1    g436(.A(new_n300), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n637), .B1(new_n638), .B2(new_n298), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n299), .A2(new_n300), .A3(new_n237), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n636), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n633), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n626), .A2(new_n628), .A3(new_n631), .A4(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n634), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT11), .B(G169gat), .ZN(new_n645));
  INV_X1    g444(.A(G197gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g446(.A(G113gat), .B(G141gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(KEYINPUT12), .Z(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n644), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n634), .A2(new_n641), .A3(new_n650), .A4(new_n643), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT94), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n652), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(G230gat), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n659), .A2(new_n204), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n215), .A2(new_n283), .A3(new_n219), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n215), .A2(new_n283), .A3(new_n219), .A4(KEYINPUT102), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT10), .ZN(new_n666));
  INV_X1    g465(.A(new_n283), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n220), .A2(new_n221), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n222), .A2(KEYINPUT10), .A3(new_n283), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n660), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n660), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n672), .B1(new_n665), .B2(new_n668), .ZN(new_n673));
  XNOR2_X1  g472(.A(G120gat), .B(G148gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(new_n446), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(G204gat), .Z(new_n676));
  OR3_X1    g475(.A1(new_n671), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n676), .B1(new_n671), .B2(new_n673), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n658), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n625), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(KEYINPUT103), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n625), .A2(new_n683), .A3(new_n680), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n552), .B(KEYINPUT104), .Z(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g488(.A(new_n571), .B1(new_n682), .B2(new_n684), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT16), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(new_n288), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n288), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n690), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT42), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n690), .A2(KEYINPUT42), .A3(new_n693), .A4(new_n694), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n697), .B(new_n698), .C1(new_n288), .C2(new_n690), .ZN(G1325gat));
  AOI21_X1  g498(.A(G15gat), .B1(new_n685), .B2(new_n591), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n701));
  INV_X1    g500(.A(new_n622), .ZN(new_n702));
  INV_X1    g501(.A(new_n623), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n622), .A2(new_n623), .A3(KEYINPUT105), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(G15gat), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT106), .Z(new_n708));
  AOI21_X1  g507(.A(new_n700), .B1(new_n685), .B2(new_n708), .ZN(G1326gat));
  NAND2_X1  g508(.A1(new_n685), .A2(new_n594), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT43), .B(G22gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1327gat));
  AOI21_X1  g511(.A(new_n265), .B1(new_n593), .B2(new_n624), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n320), .A2(new_n658), .A3(new_n679), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n715), .A2(G29gat), .A3(new_n686), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n716), .B(KEYINPUT45), .Z(new_n717));
  NAND2_X1  g516(.A1(new_n593), .A2(new_n624), .ZN(new_n718));
  INV_X1    g517(.A(new_n265), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n713), .A2(KEYINPUT44), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n714), .ZN(new_n725));
  OAI21_X1  g524(.A(G29gat), .B1(new_n725), .B2(new_n686), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n717), .A2(new_n726), .ZN(G1328gat));
  OAI21_X1  g526(.A(G36gat), .B1(new_n725), .B2(new_n571), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n715), .A2(G36gat), .A3(new_n571), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT46), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1329gat));
  INV_X1    g530(.A(new_n591), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n715), .A2(G43gat), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n702), .A2(new_n703), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n722), .A2(new_n735), .A3(new_n714), .A4(new_n723), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n733), .B1(new_n736), .B2(G43gat), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT47), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n722), .A2(new_n706), .A3(new_n714), .A4(new_n723), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n739), .A2(KEYINPUT108), .A3(G43gat), .ZN(new_n740));
  AOI21_X1  g539(.A(KEYINPUT108), .B1(new_n739), .B2(G43gat), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n740), .A2(new_n741), .A3(new_n733), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n743));
  OAI21_X1  g542(.A(new_n738), .B1(new_n742), .B2(new_n743), .ZN(G1330gat));
  NAND4_X1  g543(.A1(new_n724), .A2(G50gat), .A3(new_n594), .A4(new_n714), .ZN(new_n745));
  INV_X1    g544(.A(G50gat), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(new_n715), .B2(new_n411), .ZN(new_n747));
  AND3_X1   g546(.A1(new_n745), .A2(KEYINPUT48), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT48), .B1(new_n745), .B2(new_n747), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(G1331gat));
  INV_X1    g549(.A(new_n325), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n718), .A2(new_n679), .A3(new_n658), .A4(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n686), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(new_n271), .ZN(G1332gat));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n625), .A2(KEYINPUT109), .A3(new_n679), .A4(new_n658), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  AND2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n758), .B(new_n613), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  XOR2_X1   g560(.A(KEYINPUT110), .B(KEYINPUT111), .Z(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n571), .B1(new_n756), .B2(new_n757), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n761), .B(new_n763), .C1(new_n764), .C2(new_n759), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n764), .A2(new_n759), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n760), .A2(new_n759), .ZN(new_n767));
  AOI211_X1 g566(.A(new_n571), .B(new_n767), .C1(new_n756), .C2(new_n757), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n762), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n765), .A2(new_n769), .ZN(G1333gat));
  NAND3_X1  g569(.A1(new_n758), .A2(G71gat), .A3(new_n706), .ZN(new_n771));
  INV_X1    g570(.A(G71gat), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n752), .B2(new_n732), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n594), .ZN(new_n776));
  XNOR2_X1  g575(.A(KEYINPUT112), .B(G78gat), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1335gat));
  AND2_X1   g577(.A1(new_n677), .A2(new_n678), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n320), .A2(new_n779), .A3(new_n657), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n722), .A2(new_n723), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n782), .A2(new_n207), .A3(new_n686), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n320), .A2(new_n657), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n713), .A2(KEYINPUT51), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n779), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n718), .A2(new_n719), .A3(new_n784), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n791), .A2(new_n786), .A3(new_n785), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n788), .A2(new_n687), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n783), .B1(new_n793), .B2(new_n207), .ZN(G1336gat));
  AOI21_X1  g593(.A(new_n206), .B1(new_n781), .B2(new_n613), .ZN(new_n795));
  INV_X1    g594(.A(G92gat), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n613), .A2(new_n796), .ZN(new_n797));
  AOI211_X1 g596(.A(new_n779), .B(new_n797), .C1(new_n791), .C2(new_n785), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT52), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n788), .A2(new_n792), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n801), .B2(new_n797), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n799), .B1(new_n802), .B2(new_n795), .ZN(G1337gat));
  INV_X1    g602(.A(new_n706), .ZN(new_n804));
  OAI21_X1  g603(.A(G99gat), .B1(new_n782), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n490), .A3(new_n792), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n732), .B2(new_n806), .ZN(G1338gat));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n722), .A2(new_n594), .A3(new_n723), .A4(new_n780), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G106gat), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n411), .A2(G106gat), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n808), .B(new_n810), .C1(new_n801), .C2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n809), .A2(new_n814), .A3(G106gat), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n814), .B1(new_n809), .B2(G106gat), .ZN(new_n816));
  AOI211_X1 g615(.A(new_n779), .B(new_n812), .C1(new_n791), .C2(new_n785), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n813), .B1(new_n818), .B2(new_n808), .ZN(G1339gat));
  NOR2_X1   g618(.A1(new_n686), .A2(new_n613), .ZN(new_n820));
  INV_X1    g619(.A(new_n517), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n322), .A2(new_n779), .A3(new_n658), .A4(new_n324), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823));
  INV_X1    g622(.A(new_n649), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n639), .A2(new_n640), .A3(new_n636), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n631), .B1(new_n626), .B2(new_n628), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n827), .B1(new_n655), .B2(new_n656), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n823), .B1(new_n828), .B2(new_n779), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n669), .A2(new_n660), .A3(new_n670), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT54), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(new_n671), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n669), .A2(new_n670), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n835), .A3(new_n672), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n676), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n830), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n676), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n839), .B1(new_n671), .B2(new_n835), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n840), .B(KEYINPUT55), .C1(new_n671), .C2(new_n832), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n657), .A2(new_n677), .A3(new_n838), .A4(new_n841), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n653), .B(new_n654), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n843), .A2(new_n679), .A3(KEYINPUT115), .A4(new_n827), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n838), .A2(new_n841), .A3(new_n677), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n265), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n828), .ZN(new_n848));
  AOI22_X1  g647(.A1(new_n845), .A2(new_n265), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n822), .B1(new_n849), .B2(new_n320), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n820), .A2(new_n821), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n657), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n679), .ZN(new_n854));
  XOR2_X1   g653(.A(KEYINPUT116), .B(G120gat), .Z(new_n855));
  XNOR2_X1  g654(.A(new_n854), .B(new_n855), .ZN(G1341gat));
  NAND2_X1  g655(.A1(new_n851), .A2(new_n320), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g657(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n851), .A2(new_n719), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n861));
  XOR2_X1   g660(.A(new_n860), .B(new_n861), .Z(G1343gat));
  OAI21_X1  g661(.A(new_n687), .B1(new_n704), .B2(new_n705), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n850), .A2(new_n594), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT120), .B1(new_n863), .B2(new_n864), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n613), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n658), .A2(G141gat), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT58), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n341), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n820), .A2(new_n734), .ZN(new_n873));
  INV_X1    g672(.A(new_n320), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n843), .A2(new_n679), .A3(new_n827), .ZN(new_n875));
  AOI22_X1  g674(.A1(new_n842), .A2(new_n875), .B1(new_n264), .B2(new_n263), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n265), .A2(new_n846), .A3(new_n828), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT117), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n880), .B(new_n874), .C1(new_n876), .C2(new_n877), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n879), .A2(new_n822), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(KEYINPUT57), .A3(new_n594), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n864), .A2(new_n884), .ZN(new_n885));
  AOI211_X1 g684(.A(new_n658), .B(new_n873), .C1(new_n883), .C2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n871), .B1(new_n872), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n864), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n734), .A2(KEYINPUT105), .ZN(new_n889));
  INV_X1    g688(.A(new_n705), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n686), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n888), .A2(new_n891), .A3(new_n571), .A4(new_n870), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n865), .A2(KEYINPUT118), .A3(new_n571), .A4(new_n870), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n873), .B1(new_n883), .B2(new_n885), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n872), .B1(new_n897), .B2(new_n657), .ZN(new_n898));
  OAI211_X1 g697(.A(KEYINPUT119), .B(KEYINPUT58), .C1(new_n896), .C2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n894), .B(new_n895), .C1(new_n886), .C2(new_n872), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT119), .B1(new_n901), .B2(KEYINPUT58), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n887), .B1(new_n900), .B2(new_n902), .ZN(G1344gat));
  NAND3_X1  g702(.A1(new_n869), .A2(new_n339), .A3(new_n679), .ZN(new_n904));
  AOI211_X1 g703(.A(KEYINPUT59), .B(new_n339), .C1(new_n897), .C2(new_n679), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906));
  INV_X1    g705(.A(new_n873), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n864), .A2(KEYINPUT57), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n847), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT121), .B1(new_n265), .B2(new_n846), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n848), .A3(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n876), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n320), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n822), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n884), .B(new_n594), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n907), .A2(new_n908), .A3(new_n679), .A4(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n906), .B1(new_n917), .B2(G148gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n904), .B1(new_n905), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT122), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n904), .B(new_n921), .C1(new_n905), .C2(new_n918), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1345gat));
  AOI21_X1  g722(.A(G155gat), .B1(new_n869), .B2(new_n320), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n874), .A2(new_n355), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n897), .B2(new_n925), .ZN(G1346gat));
  NAND2_X1  g725(.A1(new_n897), .A2(new_n719), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n335), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n265), .A2(new_n335), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n869), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n929), .B1(new_n869), .B2(new_n930), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n928), .B1(new_n931), .B2(new_n932), .ZN(G1347gat));
  AND2_X1   g732(.A1(new_n850), .A2(new_n686), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n517), .A2(new_n571), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT125), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT125), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n934), .A2(new_n938), .A3(new_n935), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n445), .B1(new_n940), .B2(new_n657), .ZN(new_n941));
  INV_X1    g740(.A(new_n935), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n942), .A2(KEYINPUT124), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(KEYINPUT124), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n934), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n945), .A2(G169gat), .A3(new_n658), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n941), .A2(new_n946), .ZN(G1348gat));
  NAND3_X1  g746(.A1(new_n940), .A2(G176gat), .A3(new_n679), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n446), .B1(new_n945), .B2(new_n779), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(G1349gat));
  NAND2_X1  g749(.A1(new_n320), .A2(new_n449), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n945), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n937), .A2(new_n320), .A3(new_n939), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n952), .B1(new_n953), .B2(G183gat), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(KEYINPUT60), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n954), .B(new_n956), .ZN(G1350gat));
  OR3_X1    g756(.A1(new_n945), .A2(G190gat), .A3(new_n265), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT61), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n940), .A2(new_n719), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n959), .B1(new_n960), .B2(G190gat), .ZN(new_n961));
  AOI211_X1 g760(.A(KEYINPUT61), .B(new_n239), .C1(new_n940), .C2(new_n719), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(G1351gat));
  NOR3_X1   g762(.A1(new_n706), .A2(new_n571), .A3(new_n687), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n965), .A2(new_n864), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n966), .A2(new_n646), .A3(new_n657), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n908), .A2(new_n916), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n968), .A2(new_n964), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n969), .A2(new_n657), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n970), .B2(new_n646), .ZN(G1352gat));
  XNOR2_X1  g770(.A(KEYINPUT127), .B(G204gat), .ZN(new_n972));
  NOR4_X1   g771(.A1(new_n965), .A2(new_n779), .A3(new_n864), .A4(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n968), .A2(new_n679), .A3(new_n964), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(new_n972), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n973), .A2(new_n974), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n975), .A2(new_n977), .A3(new_n978), .ZN(G1353gat));
  NAND3_X1  g778(.A1(new_n966), .A2(new_n302), .A3(new_n320), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n969), .A2(new_n320), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n981), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n982));
  AOI21_X1  g781(.A(KEYINPUT63), .B1(new_n981), .B2(G211gat), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(G1354gat));
  AOI21_X1  g783(.A(G218gat), .B1(new_n966), .B2(new_n719), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n265), .A2(new_n246), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n985), .B1(new_n969), .B2(new_n986), .ZN(G1355gat));
endmodule


