//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985;
  XNOR2_X1  g000(.A(KEYINPUT67), .B(G237), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT28), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT11), .ZN(new_n195));
  INV_X1    g009(.A(G134), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n195), .B1(new_n196), .B2(G137), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(G137), .ZN(new_n198));
  INV_X1    g012(.A(G137), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT11), .A3(G134), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(new_n198), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G131), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n197), .A2(new_n200), .A3(new_n203), .A4(new_n198), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OR2_X1    g024(.A1(KEYINPUT0), .A2(G128), .ZN(new_n211));
  NAND2_X1  g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n208), .A2(G146), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n217), .B1(new_n206), .B2(G143), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n208), .A2(KEYINPUT65), .A3(G146), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n216), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(KEYINPUT0), .A3(G128), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n210), .A2(KEYINPUT64), .A3(new_n211), .A4(new_n212), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n205), .A2(new_n215), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT1), .B1(new_n208), .B2(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G128), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n220), .A2(new_n226), .B1(new_n228), .B2(new_n210), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n199), .A2(G134), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n196), .A2(G137), .ZN(new_n231));
  OAI21_X1  g045(.A(G131), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n204), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n224), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n218), .A2(new_n219), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(new_n207), .A3(new_n226), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n228), .A2(new_n210), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n204), .A2(new_n232), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(new_n239), .A3(KEYINPUT66), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n223), .A2(new_n234), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G116), .ZN(new_n243));
  INV_X1    g057(.A(G116), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G119), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT2), .B(G113), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n238), .A2(new_n239), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n249), .B1(new_n223), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n241), .A2(new_n249), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n223), .A2(new_n250), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT68), .B1(new_n254), .B2(new_n249), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n194), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT28), .B1(new_n254), .B2(new_n249), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n193), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n241), .A2(new_n249), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT30), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n223), .A2(new_n260), .A3(new_n250), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n223), .A2(new_n234), .A3(new_n240), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n261), .B1(KEYINPUT30), .B2(new_n262), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n259), .B(new_n192), .C1(new_n263), .C2(new_n249), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT31), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n254), .A2(new_n260), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n262), .A2(KEYINPUT30), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n248), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT31), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n269), .A2(new_n270), .A3(new_n259), .A4(new_n192), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n258), .A2(new_n265), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT69), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT69), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n258), .A2(new_n265), .A3(new_n274), .A4(new_n271), .ZN(new_n275));
  NOR2_X1   g089(.A1(G472), .A2(G902), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT32), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT32), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n273), .A2(new_n279), .A3(new_n275), .A4(new_n276), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G472), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n251), .A2(new_n252), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n255), .A2(new_n259), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n257), .B1(new_n284), .B2(KEYINPUT28), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT29), .B1(new_n285), .B2(new_n192), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n269), .A2(new_n259), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n193), .ZN(new_n288));
  AOI21_X1  g102(.A(G902), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n262), .A2(new_n248), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n259), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT70), .B1(new_n291), .B2(KEYINPUT28), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n293));
  AOI211_X1 g107(.A(new_n293), .B(new_n194), .C1(new_n259), .C2(new_n290), .ZN(new_n294));
  OR2_X1    g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n257), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n295), .A2(KEYINPUT29), .A3(new_n296), .A4(new_n192), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n282), .B1(new_n289), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT71), .B1(new_n281), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT71), .ZN(new_n301));
  AOI211_X1 g115(.A(new_n301), .B(new_n298), .C1(new_n278), .C2(new_n280), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G221), .ZN(new_n304));
  XOR2_X1   g118(.A(KEYINPUT9), .B(G234), .Z(new_n305));
  INV_X1    g119(.A(G902), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(G110), .B(G140), .ZN(new_n308));
  INV_X1    g122(.A(G227), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(G953), .ZN(new_n310));
  XOR2_X1   g124(.A(new_n308), .B(new_n310), .Z(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n205), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT3), .ZN(new_n314));
  INV_X1    g128(.A(G104), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(G107), .ZN(new_n316));
  INV_X1    g130(.A(G107), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(KEYINPUT3), .A3(G104), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G101), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n315), .A2(G107), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n317), .B2(G104), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n317), .A2(G104), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n315), .A2(KEYINPUT77), .A3(G107), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G101), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT10), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n329), .A2(new_n229), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n319), .A2(new_n321), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G101), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n332), .B1(new_n334), .B2(KEYINPUT4), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n316), .A2(new_n318), .B1(new_n315), .B2(G107), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(new_n320), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(KEYINPUT76), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n338), .B1(new_n336), .B2(new_n320), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n335), .A2(new_n339), .B1(new_n334), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n215), .A2(new_n221), .A3(new_n222), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n331), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n322), .A2(new_n328), .ZN(new_n345));
  INV_X1    g159(.A(new_n236), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n220), .B1(G128), .B2(new_n227), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n330), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n313), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n340), .A2(new_n334), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT76), .B1(new_n337), .B2(new_n338), .ZN(new_n352));
  NOR4_X1   g166(.A1(new_n336), .A2(new_n332), .A3(KEYINPUT4), .A4(new_n320), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n343), .B(new_n351), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n331), .ZN(new_n355));
  AND4_X1   g169(.A1(new_n313), .A2(new_n354), .A3(new_n349), .A4(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n312), .B1(new_n350), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n344), .A2(new_n313), .A3(new_n349), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT78), .B1(new_n345), .B2(new_n238), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n329), .A2(new_n360), .A3(new_n229), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(new_n348), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n205), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT12), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT12), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n362), .A2(new_n365), .A3(new_n205), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n358), .A2(new_n364), .A3(new_n311), .A4(new_n366), .ZN(new_n367));
  AOI211_X1 g181(.A(G469), .B(G902), .C1(new_n357), .C2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G469), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(new_n306), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  OR3_X1    g185(.A1(new_n350), .A2(new_n356), .A3(new_n312), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n358), .A2(new_n364), .A3(new_n366), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n312), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G469), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n307), .B1(new_n371), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G125), .B(G140), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n206), .ZN(new_n379));
  NAND2_X1  g193(.A1(KEYINPUT74), .A2(G125), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(G140), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT16), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT16), .ZN(new_n383));
  INV_X1    g197(.A(G125), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n383), .B1(new_n384), .B2(G140), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n206), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  XOR2_X1   g201(.A(G119), .B(G128), .Z(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(KEYINPUT73), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT24), .B(G110), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n242), .A2(G128), .ZN(new_n393));
  OR2_X1    g207(.A1(new_n393), .A2(KEYINPUT23), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(KEYINPUT23), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n394), .B(new_n395), .C1(G119), .C2(new_n225), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(G110), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n379), .B(new_n387), .C1(new_n392), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n389), .A2(new_n391), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n396), .A2(G110), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n382), .A2(new_n385), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(G146), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n399), .B(new_n400), .C1(new_n402), .C2(new_n386), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT22), .B(G137), .ZN(new_n405));
  INV_X1    g219(.A(G234), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n304), .A2(new_n406), .A3(G953), .ZN(new_n407));
  XOR2_X1   g221(.A(new_n405), .B(new_n407), .Z(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  OR2_X1    g224(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n398), .A2(new_n403), .A3(new_n408), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n410), .A2(new_n306), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  AND2_X1   g227(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(KEYINPUT75), .A3(KEYINPUT25), .ZN(new_n416));
  OAI21_X1  g230(.A(G217), .B1(new_n406), .B2(G902), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n417), .B(KEYINPUT72), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n410), .A2(new_n412), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n418), .A2(G902), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n303), .A2(new_n377), .A3(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(G113), .B(G122), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT83), .B(G104), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n426), .B(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  MUX2_X1   g243(.A(new_n378), .B(new_n381), .S(KEYINPUT19), .Z(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(G146), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n188), .A2(G214), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(new_n208), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G131), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n432), .B(G143), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n203), .ZN(new_n436));
  AOI211_X1 g250(.A(new_n386), .B(new_n431), .C1(new_n434), .C2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(KEYINPUT18), .A2(G131), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n381), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n379), .B1(new_n440), .B2(new_n206), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT18), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n439), .B(new_n441), .C1(new_n434), .C2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n429), .B1(new_n437), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT17), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n434), .A2(new_n436), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n433), .A2(KEYINPUT17), .A3(G131), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT84), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n449), .B1(new_n402), .B2(new_n386), .ZN(new_n450));
  OR3_X1    g264(.A1(new_n402), .A2(new_n386), .A3(new_n449), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n447), .A2(new_n448), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n443), .A3(new_n428), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n445), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G475), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n455), .A3(new_n306), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT20), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(G475), .B1(new_n445), .B2(new_n453), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(KEYINPUT20), .A3(new_n306), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(G234), .A2(G237), .ZN(new_n462));
  INV_X1    g276(.A(G953), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(G952), .A3(new_n463), .ZN(new_n464));
  XOR2_X1   g278(.A(new_n464), .B(KEYINPUT87), .Z(new_n465));
  XOR2_X1   g279(.A(KEYINPUT21), .B(G898), .Z(new_n466));
  NAND3_X1  g280(.A1(new_n462), .A2(G902), .A3(G953), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n305), .A2(G217), .A3(new_n463), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(G116), .B(G122), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n317), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n244), .A2(KEYINPUT14), .A3(G122), .ZN(new_n473));
  INV_X1    g287(.A(new_n471), .ZN(new_n474));
  OAI211_X1 g288(.A(G107), .B(new_n473), .C1(new_n474), .C2(KEYINPUT14), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n208), .A2(G128), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n225), .A2(G143), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT85), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT85), .B1(new_n476), .B2(new_n477), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n479), .A2(G134), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n476), .A2(new_n477), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT85), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n196), .B1(new_n484), .B2(new_n478), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n472), .B(new_n475), .C1(new_n481), .C2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT86), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(G134), .B1(new_n479), .B2(new_n480), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n484), .A2(new_n478), .A3(new_n196), .ZN(new_n490));
  AOI22_X1  g304(.A1(new_n489), .A2(new_n490), .B1(new_n317), .B2(new_n471), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(KEYINPUT86), .A3(new_n475), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n471), .B(new_n317), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT13), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n495), .B(G134), .C1(KEYINPUT13), .C2(new_n476), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n490), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n470), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n497), .ZN(new_n499));
  AOI211_X1 g313(.A(new_n499), .B(new_n469), .C1(new_n488), .C2(new_n492), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n306), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G478), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(KEYINPUT15), .ZN(new_n503));
  XOR2_X1   g317(.A(new_n501), .B(new_n503), .Z(new_n504));
  INV_X1    g318(.A(new_n453), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n428), .B1(new_n452), .B2(new_n443), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n306), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G475), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n461), .A2(new_n468), .A3(new_n504), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT88), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n458), .A2(new_n508), .A3(new_n460), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT88), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n512), .A2(new_n513), .A3(new_n468), .A4(new_n504), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(G214), .B1(G237), .B2(G902), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(G210), .B1(G237), .B2(G902), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n229), .A2(new_n384), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n343), .B2(new_n384), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n463), .A2(G224), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n243), .A2(new_n245), .A3(KEYINPUT5), .ZN(new_n524));
  OR3_X1    g338(.A1(new_n244), .A2(KEYINPUT5), .A3(G119), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(G113), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT79), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n524), .A2(new_n525), .A3(KEYINPUT79), .A4(G113), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n246), .A2(new_n247), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(new_n345), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT80), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n351), .B(new_n248), .C1(new_n352), .C2(new_n353), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n531), .B1(new_n528), .B2(new_n529), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT80), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n537), .A3(new_n345), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n534), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  XOR2_X1   g353(.A(G110), .B(G122), .Z(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT6), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT81), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n540), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n534), .A2(new_n548), .A3(new_n535), .A4(new_n538), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n549), .A2(KEYINPUT6), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n535), .A2(new_n538), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n537), .B1(new_n536), .B2(new_n345), .ZN(new_n552));
  OAI211_X1 g366(.A(KEYINPUT81), .B(new_n540), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n547), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT82), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n547), .A2(new_n550), .A3(KEYINPUT82), .A4(new_n553), .ZN(new_n557));
  AOI211_X1 g371(.A(new_n523), .B(new_n545), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n521), .A2(G224), .A3(new_n463), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n536), .A2(new_n329), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n540), .B(KEYINPUT8), .Z(new_n561));
  AND2_X1   g375(.A1(new_n532), .A2(new_n526), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n560), .B(new_n561), .C1(new_n329), .C2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT7), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n520), .B(new_n522), .C1(new_n343), .C2(new_n384), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n559), .B(new_n563), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n521), .A2(new_n564), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n549), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n306), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n519), .B1(new_n558), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n523), .ZN(new_n571));
  INV_X1    g385(.A(new_n553), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT81), .B1(new_n539), .B2(new_n540), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT82), .B1(new_n574), .B2(new_n550), .ZN(new_n575));
  INV_X1    g389(.A(new_n557), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n544), .B(new_n571), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n569), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n518), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n517), .B1(new_n570), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n515), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n425), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(new_n320), .ZN(G3));
  INV_X1    g397(.A(KEYINPUT89), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT33), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(KEYINPUT89), .A2(KEYINPUT33), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n586), .B(new_n587), .C1(new_n498), .C2(new_n500), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n486), .A2(new_n487), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT86), .B1(new_n491), .B2(new_n475), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n497), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n469), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n493), .A2(new_n497), .A3(new_n470), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n592), .A2(new_n584), .A3(new_n585), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(G478), .A3(new_n306), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT90), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n501), .A2(new_n502), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT90), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n595), .A2(new_n599), .A3(G478), .A4(new_n306), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT91), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT91), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n597), .A2(new_n603), .A3(new_n598), .A4(new_n600), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n512), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n605), .A2(new_n468), .A3(new_n580), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n273), .A2(new_n306), .A3(new_n275), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(G472), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n277), .ZN(new_n609));
  INV_X1    g423(.A(new_n377), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n609), .A2(new_n610), .A3(new_n423), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT34), .B(G104), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G6));
  AOI21_X1  g428(.A(new_n545), .B1(new_n556), .B2(new_n557), .ZN(new_n615));
  AOI211_X1 g429(.A(new_n519), .B(new_n569), .C1(new_n615), .C2(new_n571), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n518), .B1(new_n577), .B2(new_n578), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n468), .B(new_n516), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n511), .A2(new_n504), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n611), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT35), .B(G107), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G9));
  XOR2_X1   g438(.A(new_n404), .B(KEYINPUT92), .Z(new_n625));
  NOR2_X1   g439(.A1(new_n409), .A2(KEYINPUT36), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n404), .B(KEYINPUT92), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n628), .B1(KEYINPUT36), .B2(new_n409), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n627), .A2(new_n629), .A3(new_n421), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n419), .A2(new_n630), .A3(KEYINPUT93), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT93), .B1(new_n419), .B2(new_n630), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n609), .A2(new_n610), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n515), .A2(new_n580), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT37), .B(G110), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT94), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n635), .B(new_n637), .ZN(G12));
  OAI21_X1  g452(.A(new_n465), .B1(G900), .B2(new_n467), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n620), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n516), .B1(new_n616), .B2(new_n617), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n633), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n303), .A2(new_n377), .A3(new_n641), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G128), .ZN(G30));
  AND2_X1   g459(.A1(new_n419), .A2(new_n630), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT95), .B(KEYINPUT39), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n639), .B(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n377), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT40), .ZN(new_n651));
  NOR4_X1   g465(.A1(new_n651), .A2(new_n504), .A3(new_n512), .A4(new_n517), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n570), .A2(new_n579), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT38), .ZN(new_n654));
  INV_X1    g468(.A(new_n287), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n193), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n306), .B1(new_n291), .B2(new_n192), .ZN(new_n657));
  OAI21_X1  g471(.A(G472), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n281), .A2(new_n658), .ZN(new_n659));
  AND4_X1   g473(.A1(new_n646), .A2(new_n652), .A3(new_n654), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(new_n208), .ZN(G45));
  AOI211_X1 g475(.A(new_n640), .B(new_n512), .C1(new_n602), .C2(new_n604), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n303), .A2(new_n377), .A3(new_n643), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G146), .ZN(G48));
  NAND2_X1  g478(.A1(new_n357), .A2(new_n367), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n306), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(G469), .ZN(new_n667));
  INV_X1    g481(.A(new_n307), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n665), .A2(new_n369), .A3(new_n306), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT96), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n369), .B1(new_n665), .B2(new_n306), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n368), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT96), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n673), .A2(new_n674), .A3(new_n668), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT97), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(KEYINPUT97), .B1(new_n671), .B2(new_n675), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n303), .A2(new_n606), .A3(new_n680), .A4(new_n424), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  NAND4_X1  g497(.A1(new_n303), .A2(new_n680), .A3(new_n424), .A4(new_n621), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G116), .ZN(G18));
  INV_X1    g499(.A(KEYINPUT98), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(new_n642), .B2(new_n676), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n674), .B1(new_n673), .B2(new_n668), .ZN(new_n688));
  NOR4_X1   g502(.A1(new_n672), .A2(new_n368), .A3(KEYINPUT96), .A4(new_n307), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n580), .A2(new_n690), .A3(KEYINPUT98), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n633), .B1(new_n510), .B2(new_n514), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n692), .A2(new_n303), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT99), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT99), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n692), .A2(new_n303), .A3(new_n696), .A4(new_n693), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G119), .ZN(G21));
  NOR3_X1   g513(.A1(new_n642), .A2(new_n504), .A3(new_n512), .ZN(new_n700));
  INV_X1    g514(.A(new_n276), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n296), .B1(new_n292), .B2(new_n294), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n193), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n265), .A2(new_n271), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n701), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AOI211_X1 g519(.A(new_n423), .B(new_n705), .C1(new_n607), .C2(G472), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n680), .A2(new_n468), .A3(new_n700), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G122), .ZN(G24));
  AOI211_X1 g522(.A(new_n705), .B(new_n646), .C1(G472), .C2(new_n607), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n605), .A2(new_n709), .A3(new_n639), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n692), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G125), .ZN(G27));
  NAND2_X1  g526(.A1(new_n281), .A2(new_n299), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT101), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(new_n714), .A3(new_n424), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n298), .B1(new_n278), .B2(new_n280), .ZN(new_n716));
  OAI21_X1  g530(.A(KEYINPUT101), .B1(new_n716), .B2(new_n423), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT100), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n374), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n373), .A2(KEYINPUT100), .A3(new_n312), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(G469), .A3(new_n372), .A4(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n307), .B1(new_n371), .B2(new_n722), .ZN(new_n723));
  AND4_X1   g537(.A1(new_n516), .A2(new_n570), .A3(new_n723), .A4(new_n579), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n718), .A2(new_n662), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n713), .A2(new_n301), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n716), .A2(KEYINPUT71), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n424), .A4(new_n724), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n605), .A2(new_n639), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(KEYINPUT42), .ZN(new_n731));
  AOI22_X1  g545(.A1(new_n725), .A2(KEYINPUT42), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT102), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT42), .ZN(new_n735));
  INV_X1    g549(.A(new_n724), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n736), .B1(new_n715), .B2(new_n717), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n735), .B1(new_n737), .B2(new_n662), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n728), .A2(KEYINPUT42), .A3(new_n730), .ZN(new_n739));
  OAI21_X1  g553(.A(KEYINPUT102), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n734), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G131), .ZN(G33));
  NAND4_X1  g556(.A1(new_n303), .A2(new_n424), .A3(new_n641), .A4(new_n724), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G134), .ZN(G36));
  OR2_X1    g558(.A1(new_n375), .A2(KEYINPUT45), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n720), .A2(KEYINPUT45), .A3(new_n372), .A4(new_n721), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(G469), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT103), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n745), .A2(KEYINPUT103), .A3(G469), .A4(new_n746), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n370), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n751), .A2(KEYINPUT46), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n669), .B1(new_n751), .B2(KEYINPUT46), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n668), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n754), .A2(new_n648), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n653), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n516), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n602), .A2(new_n604), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n512), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n646), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n609), .A3(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n756), .A2(new_n759), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G137), .ZN(G39));
  NOR2_X1   g584(.A1(KEYINPUT104), .A2(KEYINPUT47), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n754), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n772), .B1(new_n754), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n758), .A2(new_n424), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n303), .A2(new_n730), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XOR2_X1   g592(.A(KEYINPUT105), .B(G140), .Z(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(G42));
  NOR2_X1   g594(.A1(G952), .A2(G953), .ZN(new_n781));
  XOR2_X1   g595(.A(new_n781), .B(KEYINPUT114), .Z(new_n782));
  INV_X1    g596(.A(new_n465), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n763), .A2(new_n783), .A3(new_n706), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n692), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n758), .A2(new_n676), .ZN(new_n787));
  INV_X1    g601(.A(new_n659), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n787), .A2(new_n783), .A3(new_n424), .A4(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n605), .ZN(new_n790));
  OAI211_X1 g604(.A(G952), .B(new_n463), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n763), .A2(new_n783), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n718), .A3(new_n787), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n793), .A2(KEYINPUT48), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(KEYINPUT48), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n672), .A2(new_n368), .A3(new_n668), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n785), .B(new_n759), .C1(new_n774), .C2(new_n797), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n654), .A2(new_n516), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n784), .A2(new_n676), .A3(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT50), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n792), .A2(new_n709), .A3(new_n787), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n789), .A2(new_n511), .A3(new_n760), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n804), .B1(new_n800), .B2(new_n801), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n798), .A2(new_n802), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n806), .A2(KEYINPUT112), .A3(KEYINPUT51), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT51), .B1(new_n806), .B2(KEYINPUT112), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n786), .B(new_n796), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT113), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n809), .B(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n812));
  OAI21_X1  g626(.A(KEYINPUT107), .B1(new_n618), .B2(new_n620), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT107), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n580), .A2(new_n814), .A3(new_n468), .A4(new_n619), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n611), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT108), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n635), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n612), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n817), .B1(new_n816), .B2(new_n635), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n819), .A2(new_n582), .A3(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n681), .A2(new_n684), .A3(new_n707), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT106), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n698), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n823), .B1(new_n698), .B2(new_n822), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n741), .B(new_n821), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT109), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n605), .A2(new_n709), .A3(new_n639), .A4(new_n723), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n300), .A2(new_n302), .A3(new_n610), .ZN(new_n829));
  INV_X1    g643(.A(new_n504), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n633), .A2(new_n511), .A3(new_n830), .A4(new_n640), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n828), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n827), .B(new_n743), .C1(new_n832), .C2(new_n758), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n726), .A2(new_n377), .A3(new_n727), .A4(new_n831), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n662), .A2(new_n709), .A3(new_n723), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n758), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n641), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n728), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT109), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n833), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n764), .A2(new_n640), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n700), .A2(new_n659), .A3(new_n723), .A4(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n644), .A2(new_n663), .A3(new_n711), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT52), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n829), .B(new_n643), .C1(new_n641), .C2(new_n662), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n845), .A2(new_n846), .A3(new_n711), .A4(new_n842), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n840), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n812), .B1(new_n826), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n582), .ZN(new_n850));
  INV_X1    g664(.A(new_n820), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n850), .A2(new_n851), .A3(new_n612), .A4(new_n818), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n698), .A2(new_n822), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT106), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n698), .A2(new_n822), .A3(new_n823), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n833), .A2(new_n839), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n844), .A2(new_n847), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n856), .A2(KEYINPUT53), .A3(new_n741), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n849), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT54), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT110), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT111), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n698), .A2(new_n732), .A3(new_n822), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(new_n852), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n859), .A2(new_n864), .A3(KEYINPUT53), .A4(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n840), .A2(KEYINPUT53), .A3(new_n844), .A4(new_n847), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n821), .A2(new_n698), .A3(new_n732), .A4(new_n822), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT111), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n872), .A3(new_n849), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT110), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n861), .A2(new_n874), .A3(KEYINPUT54), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n863), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n782), .B1(new_n811), .B2(new_n876), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n673), .B(KEYINPUT49), .Z(new_n878));
  NOR3_X1   g692(.A1(new_n654), .A2(new_n423), .A3(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n761), .A2(new_n659), .A3(new_n307), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n516), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n877), .A2(new_n881), .ZN(G75));
  NOR2_X1   g696(.A1(new_n463), .A2(G952), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n849), .A2(new_n870), .A3(new_n867), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(G902), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(KEYINPUT116), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT116), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n885), .A2(new_n888), .A3(G902), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n887), .A2(new_n519), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n615), .A2(new_n571), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n558), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT55), .ZN(new_n893));
  XNOR2_X1  g707(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n884), .B1(new_n890), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n885), .A2(G210), .A3(G902), .ZN(new_n897));
  OR2_X1    g711(.A1(new_n897), .A2(KEYINPUT115), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT56), .B1(new_n897), .B2(KEYINPUT115), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n893), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n896), .A2(new_n900), .ZN(G51));
  NAND2_X1  g715(.A1(new_n885), .A2(KEYINPUT54), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n873), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n370), .B(KEYINPUT118), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT57), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n904), .A2(KEYINPUT57), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n665), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n887), .A2(new_n749), .A3(new_n750), .A4(new_n889), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n883), .B1(new_n908), .B2(new_n909), .ZN(G54));
  AND2_X1   g724(.A1(KEYINPUT58), .A2(G475), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n887), .A2(new_n889), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n912), .A2(new_n453), .A3(new_n445), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n887), .A2(new_n454), .A3(new_n889), .A4(new_n911), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n913), .A2(new_n884), .A3(new_n914), .ZN(G60));
  XNOR2_X1  g729(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n916));
  NAND2_X1  g730(.A1(G478), .A2(G902), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n916), .B(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n872), .B1(new_n871), .B2(new_n849), .ZN(new_n919));
  AND4_X1   g733(.A1(new_n872), .A2(new_n849), .A3(new_n870), .A4(new_n867), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n595), .B(new_n918), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT120), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n903), .A2(KEYINPUT120), .A3(new_n595), .A4(new_n918), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n595), .B1(new_n876), .B2(new_n918), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n925), .A2(new_n883), .A3(new_n926), .ZN(G63));
  NAND2_X1  g741(.A1(G217), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT60), .Z(new_n929));
  NAND2_X1  g743(.A1(new_n627), .A2(new_n629), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT121), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n885), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n885), .A2(new_n929), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n884), .B(new_n932), .C1(new_n933), .C2(new_n420), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g749(.A(new_n463), .B1(new_n466), .B2(G224), .ZN(new_n936));
  INV_X1    g750(.A(new_n856), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n936), .B1(new_n937), .B2(new_n463), .ZN(new_n938));
  INV_X1    g752(.A(G898), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n615), .B1(new_n939), .B2(G953), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n938), .B(new_n940), .ZN(G69));
  XNOR2_X1  g755(.A(new_n268), .B(new_n430), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n767), .A2(new_n759), .A3(new_n768), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n718), .A2(new_n700), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n756), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n845), .A2(new_n711), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n776), .B2(new_n777), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n945), .A2(new_n947), .A3(new_n741), .A4(new_n743), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n942), .B1(new_n948), .B2(new_n463), .ZN(new_n949));
  INV_X1    g763(.A(G900), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(G953), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT126), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n425), .A2(new_n648), .A3(new_n758), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n790), .A2(new_n620), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT123), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n769), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT124), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n769), .A2(KEYINPUT124), .A3(new_n956), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT62), .ZN(new_n962));
  OR3_X1    g776(.A1(new_n660), .A2(new_n962), .A3(new_n946), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n962), .B1(new_n660), .B2(new_n946), .ZN(new_n964));
  AOI22_X1  g778(.A1(new_n963), .A2(new_n964), .B1(new_n777), .B2(new_n776), .ZN(new_n965));
  AOI21_X1  g779(.A(G953), .B1(new_n961), .B2(new_n965), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n949), .B(new_n952), .C1(new_n966), .C2(KEYINPUT122), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT122), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n942), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(KEYINPUT125), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(G953), .B1(new_n309), .B2(new_n950), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(G72));
  NAND2_X1  g786(.A1(new_n655), .A2(new_n193), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n948), .A2(new_n937), .ZN(new_n974));
  NAND2_X1  g788(.A1(G472), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT63), .Z(new_n976));
  AOI21_X1  g790(.A(new_n973), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n961), .A2(new_n965), .A3(new_n856), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n978), .A2(new_n976), .ZN(new_n979));
  INV_X1    g793(.A(new_n656), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n884), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n861), .A2(new_n980), .A3(new_n976), .A4(new_n973), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n982), .A2(new_n983), .ZN(new_n985));
  AOI211_X1 g799(.A(new_n977), .B(new_n981), .C1(new_n984), .C2(new_n985), .ZN(G57));
endmodule


