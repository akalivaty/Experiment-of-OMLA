

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603;

  INV_X1 U323 ( .A(G106GAT), .ZN(n311) );
  XNOR2_X1 U324 ( .A(n437), .B(n436), .ZN(n438) );
  AND2_X1 U325 ( .A1(n564), .A2(n540), .ZN(n486) );
  XNOR2_X1 U326 ( .A(n324), .B(n323), .ZN(n329) );
  XNOR2_X1 U327 ( .A(n346), .B(n345), .ZN(n349) );
  XNOR2_X1 U328 ( .A(n344), .B(KEYINPUT96), .ZN(n345) );
  XNOR2_X1 U329 ( .A(n466), .B(KEYINPUT111), .ZN(n467) );
  NOR2_X1 U330 ( .A1(n601), .A2(n573), .ZN(n476) );
  XNOR2_X1 U331 ( .A(n316), .B(n315), .ZN(n319) );
  XNOR2_X1 U332 ( .A(n298), .B(KEYINPUT17), .ZN(n299) );
  XNOR2_X1 U333 ( .A(n347), .B(KEYINPUT26), .ZN(n588) );
  XNOR2_X1 U334 ( .A(n483), .B(KEYINPUT48), .ZN(n484) );
  INV_X1 U335 ( .A(KEYINPUT64), .ZN(n483) );
  XNOR2_X1 U336 ( .A(n340), .B(n304), .ZN(n305) );
  XNOR2_X1 U337 ( .A(n303), .B(G99GAT), .ZN(n304) );
  NOR2_X1 U338 ( .A1(n428), .A2(n601), .ZN(n429) );
  XNOR2_X1 U339 ( .A(n409), .B(n408), .ZN(n428) );
  INV_X1 U340 ( .A(KEYINPUT101), .ZN(n408) );
  XNOR2_X1 U341 ( .A(n439), .B(n438), .ZN(n444) );
  NOR2_X1 U342 ( .A1(n491), .A2(n490), .ZN(n580) );
  AND2_X1 U343 ( .A1(n586), .A2(n294), .ZN(n489) );
  XNOR2_X1 U344 ( .A(n423), .B(n422), .ZN(n424) );
  INV_X1 U345 ( .A(n576), .ZN(n558) );
  XNOR2_X1 U346 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U347 ( .A(n437), .B(n292), .ZN(n337) );
  AND2_X1 U348 ( .A1(G232GAT), .A2(G233GAT), .ZN(n291) );
  XOR2_X1 U349 ( .A(G190GAT), .B(G176GAT), .Z(n292) );
  XOR2_X1 U350 ( .A(n321), .B(n320), .Z(n293) );
  NOR2_X1 U351 ( .A1(n487), .A2(n538), .ZN(n294) );
  INV_X1 U352 ( .A(KEYINPUT95), .ZN(n341) );
  INV_X1 U353 ( .A(KEYINPUT25), .ZN(n344) );
  INV_X1 U354 ( .A(KEYINPUT46), .ZN(n466) );
  INV_X1 U355 ( .A(KEYINPUT45), .ZN(n475) );
  XNOR2_X1 U356 ( .A(n468), .B(n467), .ZN(n469) );
  XOR2_X1 U357 ( .A(G22GAT), .B(G155GAT), .Z(n394) );
  XOR2_X1 U358 ( .A(G78GAT), .B(KEYINPUT22), .Z(n314) );
  XNOR2_X1 U359 ( .A(n312), .B(n311), .ZN(n316) );
  XNOR2_X1 U360 ( .A(n412), .B(n291), .ZN(n413) );
  INV_X1 U361 ( .A(G64GAT), .ZN(n403) );
  XNOR2_X1 U362 ( .A(n414), .B(n413), .ZN(n418) );
  XNOR2_X1 U363 ( .A(n322), .B(n293), .ZN(n323) );
  XNOR2_X1 U364 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U365 ( .A(n300), .B(n299), .ZN(n302) );
  XNOR2_X1 U366 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U367 ( .A(n425), .B(n424), .ZN(n427) );
  XNOR2_X1 U368 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U369 ( .A(n505), .B(G106GAT), .ZN(n506) );
  XNOR2_X1 U370 ( .A(n463), .B(G43GAT), .ZN(n464) );
  XNOR2_X1 U371 ( .A(n502), .B(n501), .ZN(G1351GAT) );
  XNOR2_X1 U372 ( .A(n498), .B(n497), .ZN(G1331GAT) );
  XOR2_X1 U373 ( .A(G71GAT), .B(KEYINPUT80), .Z(n296) );
  NAND2_X1 U374 ( .A1(G227GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U375 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U376 ( .A(KEYINPUT20), .B(n297), .ZN(n310) );
  XNOR2_X1 U377 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n300) );
  INV_X1 U378 ( .A(KEYINPUT79), .ZN(n298) );
  XNOR2_X1 U379 ( .A(G169GAT), .B(G183GAT), .ZN(n301) );
  XNOR2_X1 U380 ( .A(n302), .B(n301), .ZN(n340) );
  XOR2_X1 U381 ( .A(G113GAT), .B(KEYINPUT0), .Z(n360) );
  XOR2_X1 U382 ( .A(n360), .B(KEYINPUT78), .Z(n303) );
  XOR2_X1 U383 ( .A(G15GAT), .B(G127GAT), .Z(n395) );
  XOR2_X1 U384 ( .A(n305), .B(n395), .Z(n308) );
  XNOR2_X1 U385 ( .A(G43GAT), .B(G190GAT), .ZN(n306) );
  XNOR2_X1 U386 ( .A(n306), .B(G134GAT), .ZN(n422) );
  XOR2_X1 U387 ( .A(G176GAT), .B(G120GAT), .Z(n433) );
  XNOR2_X1 U388 ( .A(n422), .B(n433), .ZN(n307) );
  XNOR2_X1 U389 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U390 ( .A(n310), .B(n309), .ZN(n491) );
  XNOR2_X1 U391 ( .A(n394), .B(G218GAT), .ZN(n312) );
  XNOR2_X1 U392 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n313) );
  XNOR2_X1 U393 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U394 ( .A(G211GAT), .B(KEYINPUT21), .Z(n318) );
  XNOR2_X1 U395 ( .A(G197GAT), .B(KEYINPUT83), .ZN(n317) );
  XNOR2_X1 U396 ( .A(n318), .B(n317), .ZN(n334) );
  XOR2_X1 U397 ( .A(n319), .B(n334), .Z(n324) );
  XOR2_X1 U398 ( .A(G50GAT), .B(G162GAT), .Z(n412) );
  XOR2_X1 U399 ( .A(G204GAT), .B(G148GAT), .Z(n432) );
  XNOR2_X1 U400 ( .A(n412), .B(n432), .ZN(n322) );
  XOR2_X1 U401 ( .A(KEYINPUT87), .B(KEYINPUT82), .Z(n321) );
  NAND2_X1 U402 ( .A1(G228GAT), .A2(G233GAT), .ZN(n320) );
  XOR2_X1 U403 ( .A(KEYINPUT85), .B(KEYINPUT2), .Z(n326) );
  XNOR2_X1 U404 ( .A(KEYINPUT3), .B(KEYINPUT84), .ZN(n325) );
  XNOR2_X1 U405 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U406 ( .A(G141GAT), .B(n327), .Z(n364) );
  XNOR2_X1 U407 ( .A(n364), .B(KEYINPUT86), .ZN(n328) );
  XNOR2_X1 U408 ( .A(n329), .B(n328), .ZN(n487) );
  XOR2_X1 U409 ( .A(G204GAT), .B(KEYINPUT94), .Z(n331) );
  NAND2_X1 U410 ( .A1(G226GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U411 ( .A(n331), .B(n330), .ZN(n333) );
  XNOR2_X1 U412 ( .A(G36GAT), .B(G218GAT), .ZN(n332) );
  XNOR2_X1 U413 ( .A(KEYINPUT75), .B(n332), .ZN(n426) );
  XOR2_X1 U414 ( .A(n333), .B(n426), .Z(n336) );
  XNOR2_X1 U415 ( .A(G8GAT), .B(n334), .ZN(n335) );
  XNOR2_X1 U416 ( .A(n336), .B(n335), .ZN(n338) );
  XOR2_X1 U417 ( .A(G92GAT), .B(G64GAT), .Z(n437) );
  XOR2_X1 U418 ( .A(n340), .B(n339), .Z(n540) );
  INV_X1 U419 ( .A(n540), .ZN(n524) );
  NOR2_X1 U420 ( .A1(n524), .A2(n491), .ZN(n342) );
  XNOR2_X1 U421 ( .A(n342), .B(n341), .ZN(n343) );
  NOR2_X1 U422 ( .A1(n487), .A2(n343), .ZN(n346) );
  XOR2_X1 U423 ( .A(KEYINPUT27), .B(n540), .Z(n376) );
  NAND2_X1 U424 ( .A1(n487), .A2(n491), .ZN(n347) );
  NOR2_X1 U425 ( .A1(n376), .A2(n588), .ZN(n348) );
  NOR2_X1 U426 ( .A1(n349), .A2(n348), .ZN(n350) );
  XNOR2_X1 U427 ( .A(n350), .B(KEYINPUT97), .ZN(n375) );
  XOR2_X1 U428 ( .A(KEYINPUT91), .B(KEYINPUT4), .Z(n352) );
  XNOR2_X1 U429 ( .A(G1GAT), .B(KEYINPUT90), .ZN(n351) );
  XNOR2_X1 U430 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U431 ( .A(G57GAT), .B(KEYINPUT1), .Z(n354) );
  XNOR2_X1 U432 ( .A(KEYINPUT89), .B(KEYINPUT6), .ZN(n353) );
  XNOR2_X1 U433 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U434 ( .A(n356), .B(n355), .Z(n366) );
  XOR2_X1 U435 ( .A(G85GAT), .B(G162GAT), .Z(n358) );
  XNOR2_X1 U436 ( .A(G29GAT), .B(G134GAT), .ZN(n357) );
  XNOR2_X1 U437 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U438 ( .A(n360), .B(n359), .Z(n362) );
  NAND2_X1 U439 ( .A1(G225GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U440 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U441 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U442 ( .A(n366), .B(n365), .ZN(n374) );
  XOR2_X1 U443 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n368) );
  XNOR2_X1 U444 ( .A(KEYINPUT88), .B(KEYINPUT92), .ZN(n367) );
  XNOR2_X1 U445 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U446 ( .A(G155GAT), .B(G148GAT), .Z(n370) );
  XNOR2_X1 U447 ( .A(G120GAT), .B(G127GAT), .ZN(n369) );
  XNOR2_X1 U448 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U449 ( .A(n372), .B(n371), .Z(n373) );
  XOR2_X1 U450 ( .A(n374), .B(n373), .Z(n538) );
  INV_X1 U451 ( .A(n538), .ZN(n585) );
  NAND2_X1 U452 ( .A1(n375), .A2(n585), .ZN(n382) );
  OR2_X1 U453 ( .A1(n585), .A2(n376), .ZN(n563) );
  XOR2_X1 U454 ( .A(n487), .B(KEYINPUT28), .Z(n495) );
  INV_X1 U455 ( .A(n495), .ZN(n533) );
  NOR2_X1 U456 ( .A1(n563), .A2(n533), .ZN(n547) );
  INV_X1 U457 ( .A(n491), .ZN(n546) );
  XNOR2_X1 U458 ( .A(n546), .B(KEYINPUT81), .ZN(n377) );
  NAND2_X1 U459 ( .A1(n547), .A2(n377), .ZN(n380) );
  NAND2_X1 U460 ( .A1(n382), .A2(n380), .ZN(n378) );
  NAND2_X1 U461 ( .A1(n378), .A2(KEYINPUT98), .ZN(n384) );
  INV_X1 U462 ( .A(KEYINPUT98), .ZN(n379) );
  AND2_X1 U463 ( .A1(n380), .A2(n379), .ZN(n381) );
  NAND2_X1 U464 ( .A1(n382), .A2(n381), .ZN(n383) );
  NAND2_X1 U465 ( .A1(n384), .A2(n383), .ZN(n509) );
  INV_X1 U466 ( .A(KEYINPUT13), .ZN(n385) );
  NAND2_X1 U467 ( .A1(n385), .A2(KEYINPUT67), .ZN(n388) );
  INV_X1 U468 ( .A(KEYINPUT67), .ZN(n386) );
  NAND2_X1 U469 ( .A1(n386), .A2(KEYINPUT13), .ZN(n387) );
  NAND2_X1 U470 ( .A1(n388), .A2(n387), .ZN(n390) );
  XNOR2_X1 U471 ( .A(G71GAT), .B(G78GAT), .ZN(n389) );
  XNOR2_X1 U472 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U473 ( .A(G57GAT), .B(n391), .Z(n431) );
  XOR2_X1 U474 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n393) );
  XNOR2_X1 U475 ( .A(KEYINPUT77), .B(KEYINPUT76), .ZN(n392) );
  XNOR2_X1 U476 ( .A(n393), .B(n392), .ZN(n399) );
  XOR2_X1 U477 ( .A(n394), .B(G211GAT), .Z(n397) );
  XNOR2_X1 U478 ( .A(G183GAT), .B(n395), .ZN(n396) );
  XNOR2_X1 U479 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U480 ( .A(n399), .B(n398), .Z(n401) );
  NAND2_X1 U481 ( .A1(G231GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U482 ( .A(n401), .B(n400), .ZN(n406) );
  XNOR2_X1 U483 ( .A(G1GAT), .B(KEYINPUT66), .ZN(n402) );
  XNOR2_X1 U484 ( .A(n402), .B(G8GAT), .ZN(n445) );
  XNOR2_X1 U485 ( .A(n445), .B(KEYINPUT15), .ZN(n404) );
  XOR2_X1 U486 ( .A(n431), .B(n407), .Z(n595) );
  INV_X1 U487 ( .A(n595), .ZN(n573) );
  NAND2_X1 U488 ( .A1(n509), .A2(n573), .ZN(n409) );
  XOR2_X1 U489 ( .A(KEYINPUT73), .B(KEYINPUT72), .Z(n411) );
  XNOR2_X1 U490 ( .A(KEYINPUT9), .B(KEYINPUT74), .ZN(n410) );
  XNOR2_X1 U491 ( .A(n411), .B(n410), .ZN(n414) );
  XOR2_X1 U492 ( .A(G92GAT), .B(KEYINPUT65), .Z(n416) );
  XNOR2_X1 U493 ( .A(KEYINPUT10), .B(KEYINPUT11), .ZN(n415) );
  XOR2_X1 U494 ( .A(n416), .B(n415), .Z(n417) );
  XNOR2_X1 U495 ( .A(n418), .B(n417), .ZN(n425) );
  XNOR2_X1 U496 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n419) );
  XNOR2_X1 U497 ( .A(n419), .B(KEYINPUT7), .ZN(n446) );
  XOR2_X1 U498 ( .A(KEYINPUT68), .B(G85GAT), .Z(n421) );
  XNOR2_X1 U499 ( .A(G99GAT), .B(G106GAT), .ZN(n420) );
  XNOR2_X1 U500 ( .A(n421), .B(n420), .ZN(n430) );
  XNOR2_X1 U501 ( .A(n446), .B(n430), .ZN(n423) );
  XNOR2_X1 U502 ( .A(n427), .B(n426), .ZN(n576) );
  XOR2_X1 U503 ( .A(n558), .B(KEYINPUT36), .Z(n601) );
  XNOR2_X1 U504 ( .A(KEYINPUT37), .B(n429), .ZN(n503) );
  XOR2_X1 U505 ( .A(n431), .B(n430), .Z(n435) );
  XNOR2_X1 U506 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U507 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U508 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n436) );
  XOR2_X1 U509 ( .A(KEYINPUT31), .B(KEYINPUT69), .Z(n441) );
  NAND2_X1 U510 ( .A1(G230GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U511 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U512 ( .A(KEYINPUT70), .B(n442), .Z(n443) );
  XNOR2_X1 U513 ( .A(n444), .B(n443), .ZN(n592) );
  XNOR2_X1 U514 ( .A(n446), .B(n445), .ZN(n459) );
  XOR2_X1 U515 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n448) );
  NAND2_X1 U516 ( .A1(G229GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U517 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U518 ( .A(n449), .B(G22GAT), .Z(n457) );
  XOR2_X1 U519 ( .A(G36GAT), .B(G43GAT), .Z(n451) );
  XNOR2_X1 U520 ( .A(G169GAT), .B(G50GAT), .ZN(n450) );
  XNOR2_X1 U521 ( .A(n451), .B(n450), .ZN(n455) );
  XOR2_X1 U522 ( .A(G197GAT), .B(G141GAT), .Z(n453) );
  XNOR2_X1 U523 ( .A(G15GAT), .B(G113GAT), .ZN(n452) );
  XNOR2_X1 U524 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U525 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U526 ( .A(n457), .B(n456), .ZN(n458) );
  XOR2_X1 U527 ( .A(n459), .B(n458), .Z(n589) );
  INV_X1 U528 ( .A(n589), .ZN(n566) );
  NOR2_X1 U529 ( .A1(n592), .A2(n566), .ZN(n460) );
  XNOR2_X1 U530 ( .A(n460), .B(KEYINPUT71), .ZN(n511) );
  NOR2_X1 U531 ( .A1(n503), .A2(n511), .ZN(n462) );
  XOR2_X1 U532 ( .A(KEYINPUT102), .B(KEYINPUT38), .Z(n461) );
  XNOR2_X1 U533 ( .A(n462), .B(n461), .ZN(n523) );
  NOR2_X1 U534 ( .A1(n491), .A2(n523), .ZN(n465) );
  XNOR2_X1 U535 ( .A(KEYINPUT40), .B(KEYINPUT103), .ZN(n463) );
  XNOR2_X1 U536 ( .A(n465), .B(n464), .ZN(G1330GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT110), .B(n573), .Z(n579) );
  XOR2_X1 U538 ( .A(KEYINPUT41), .B(n592), .Z(n568) );
  AND2_X1 U539 ( .A1(n589), .A2(n568), .ZN(n468) );
  NOR2_X1 U540 ( .A1(n579), .A2(n469), .ZN(n471) );
  INV_X1 U541 ( .A(KEYINPUT112), .ZN(n470) );
  XNOR2_X1 U542 ( .A(n471), .B(n470), .ZN(n472) );
  NOR2_X1 U543 ( .A1(n472), .A2(n558), .ZN(n474) );
  INV_X1 U544 ( .A(KEYINPUT47), .ZN(n473) );
  XNOR2_X1 U545 ( .A(n474), .B(n473), .ZN(n482) );
  XNOR2_X1 U546 ( .A(n476), .B(n475), .ZN(n477) );
  NOR2_X1 U547 ( .A1(n592), .A2(n477), .ZN(n478) );
  XNOR2_X1 U548 ( .A(n478), .B(KEYINPUT113), .ZN(n479) );
  NOR2_X1 U549 ( .A1(n479), .A2(n589), .ZN(n480) );
  XNOR2_X1 U550 ( .A(n480), .B(KEYINPUT114), .ZN(n481) );
  NOR2_X1 U551 ( .A1(n482), .A2(n481), .ZN(n485) );
  XNOR2_X1 U552 ( .A(n485), .B(n484), .ZN(n564) );
  XNOR2_X1 U553 ( .A(n486), .B(KEYINPUT54), .ZN(n586) );
  XNOR2_X1 U554 ( .A(KEYINPUT55), .B(KEYINPUT120), .ZN(n488) );
  XNOR2_X1 U555 ( .A(n489), .B(n488), .ZN(n490) );
  NAND2_X1 U556 ( .A1(n580), .A2(n568), .ZN(n494) );
  XOR2_X1 U557 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n492) );
  XNOR2_X1 U558 ( .A(n492), .B(G176GAT), .ZN(n493) );
  XNOR2_X1 U559 ( .A(n494), .B(n493), .ZN(G1349GAT) );
  NOR2_X1 U560 ( .A1(n495), .A2(n523), .ZN(n498) );
  INV_X1 U561 ( .A(G50GAT), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n496), .B(KEYINPUT104), .ZN(n497) );
  NAND2_X1 U563 ( .A1(n580), .A2(n558), .ZN(n502) );
  XOR2_X1 U564 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n500) );
  XNOR2_X1 U565 ( .A(G190GAT), .B(KEYINPUT122), .ZN(n499) );
  NAND2_X1 U566 ( .A1(n566), .A2(n568), .ZN(n527) );
  NOR2_X1 U567 ( .A1(n503), .A2(n527), .ZN(n504) );
  XOR2_X1 U568 ( .A(KEYINPUT107), .B(n504), .Z(n543) );
  NAND2_X1 U569 ( .A1(n543), .A2(n533), .ZN(n507) );
  XOR2_X1 U570 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n505) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(G1339GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT34), .B(KEYINPUT99), .Z(n513) );
  NOR2_X1 U573 ( .A1(n558), .A2(n573), .ZN(n508) );
  XNOR2_X1 U574 ( .A(KEYINPUT16), .B(n508), .ZN(n510) );
  NAND2_X1 U575 ( .A1(n510), .A2(n509), .ZN(n526) );
  NOR2_X1 U576 ( .A1(n511), .A2(n526), .ZN(n519) );
  NAND2_X1 U577 ( .A1(n519), .A2(n538), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G1GAT), .B(n514), .ZN(G1324GAT) );
  NAND2_X1 U580 ( .A1(n519), .A2(n540), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n515), .B(KEYINPUT100), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G8GAT), .B(n516), .ZN(G1325GAT) );
  XOR2_X1 U583 ( .A(G15GAT), .B(KEYINPUT35), .Z(n518) );
  NAND2_X1 U584 ( .A1(n519), .A2(n546), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(G1326GAT) );
  NAND2_X1 U586 ( .A1(n533), .A2(n519), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n520), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U588 ( .A1(n585), .A2(n523), .ZN(n522) );
  XNOR2_X1 U589 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n521) );
  XNOR2_X1 U590 ( .A(n522), .B(n521), .ZN(G1328GAT) );
  NOR2_X1 U591 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U592 ( .A(G36GAT), .B(n525), .Z(G1329GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n529) );
  NOR2_X1 U594 ( .A1(n527), .A2(n526), .ZN(n534) );
  NAND2_X1 U595 ( .A1(n534), .A2(n538), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U597 ( .A(G57GAT), .B(n530), .ZN(G1332GAT) );
  NAND2_X1 U598 ( .A1(n534), .A2(n540), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n531), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U600 ( .A1(n546), .A2(n534), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n532), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT43), .B(KEYINPUT106), .Z(n536) );
  NAND2_X1 U603 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U604 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U605 ( .A(G78GAT), .B(n537), .ZN(G1335GAT) );
  NAND2_X1 U606 ( .A1(n538), .A2(n543), .ZN(n539) );
  XNOR2_X1 U607 ( .A(G85GAT), .B(n539), .ZN(G1336GAT) );
  XNOR2_X1 U608 ( .A(G92GAT), .B(KEYINPUT108), .ZN(n542) );
  NAND2_X1 U609 ( .A1(n540), .A2(n543), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(G1337GAT) );
  NAND2_X1 U611 ( .A1(n543), .A2(n546), .ZN(n544) );
  XNOR2_X1 U612 ( .A(G99GAT), .B(n544), .ZN(G1338GAT) );
  XOR2_X1 U613 ( .A(G113GAT), .B(KEYINPUT115), .Z(n550) );
  INV_X1 U614 ( .A(n564), .ZN(n545) );
  NAND2_X1 U615 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U616 ( .A1(n545), .A2(n548), .ZN(n559) );
  NAND2_X1 U617 ( .A1(n559), .A2(n589), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(G1340GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n552) );
  NAND2_X1 U620 ( .A1(n559), .A2(n568), .ZN(n551) );
  XNOR2_X1 U621 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U622 ( .A(G120GAT), .B(n553), .ZN(G1341GAT) );
  XNOR2_X1 U623 ( .A(G127GAT), .B(KEYINPUT118), .ZN(n557) );
  XOR2_X1 U624 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n555) );
  NAND2_X1 U625 ( .A1(n559), .A2(n579), .ZN(n554) );
  XNOR2_X1 U626 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U627 ( .A(n557), .B(n556), .ZN(G1342GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n561) );
  NAND2_X1 U629 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U630 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U631 ( .A(G134GAT), .B(n562), .Z(G1343GAT) );
  NOR2_X1 U632 ( .A1(n588), .A2(n563), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n565), .A2(n564), .ZN(n575) );
  NOR2_X1 U634 ( .A1(n566), .A2(n575), .ZN(n567) );
  XOR2_X1 U635 ( .A(G141GAT), .B(n567), .Z(G1344GAT) );
  INV_X1 U636 ( .A(n568), .ZN(n569) );
  NOR2_X1 U637 ( .A1(n569), .A2(n575), .ZN(n571) );
  XNOR2_X1 U638 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n570) );
  XNOR2_X1 U639 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U640 ( .A(G148GAT), .B(n572), .ZN(G1345GAT) );
  NOR2_X1 U641 ( .A1(n573), .A2(n575), .ZN(n574) );
  XOR2_X1 U642 ( .A(G155GAT), .B(n574), .Z(G1346GAT) );
  NOR2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U644 ( .A(G162GAT), .B(n577), .Z(G1347GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n589), .ZN(n578) );
  XNOR2_X1 U646 ( .A(G169GAT), .B(n578), .ZN(G1348GAT) );
  XOR2_X1 U647 ( .A(G183GAT), .B(KEYINPUT121), .Z(n582) );
  NAND2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U649 ( .A(n582), .B(n581), .ZN(G1350GAT) );
  XNOR2_X1 U650 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n583) );
  XNOR2_X1 U651 ( .A(n583), .B(KEYINPUT59), .ZN(n584) );
  XOR2_X1 U652 ( .A(KEYINPUT60), .B(n584), .Z(n591) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n599) );
  NAND2_X1 U655 ( .A1(n599), .A2(n589), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n591), .B(n590), .ZN(G1352GAT) );
  XOR2_X1 U657 ( .A(G204GAT), .B(KEYINPUT61), .Z(n594) );
  NAND2_X1 U658 ( .A1(n599), .A2(n592), .ZN(n593) );
  XNOR2_X1 U659 ( .A(n594), .B(n593), .ZN(G1353GAT) );
  NAND2_X1 U660 ( .A1(n599), .A2(n595), .ZN(n596) );
  XNOR2_X1 U661 ( .A(n596), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U662 ( .A(KEYINPUT62), .B(KEYINPUT125), .Z(n598) );
  XNOR2_X1 U663 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n597) );
  XNOR2_X1 U664 ( .A(n598), .B(n597), .ZN(n603) );
  INV_X1 U665 ( .A(n599), .ZN(n600) );
  NOR2_X1 U666 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U667 ( .A(n603), .B(n602), .Z(G1355GAT) );
endmodule

