//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT23), .B1(new_n187), .B2(G119), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  OAI211_X1 g003(.A(new_n188), .B(KEYINPUT73), .C1(new_n189), .C2(G128), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT73), .ZN(new_n191));
  OAI211_X1 g005(.A(G119), .B(new_n187), .C1(new_n191), .C2(KEYINPUT23), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(G119), .B(G128), .ZN(new_n194));
  XOR2_X1   g008(.A(KEYINPUT24), .B(G110), .Z(new_n195));
  AOI22_X1  g009(.A1(new_n193), .A2(G110), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(G125), .B(G140), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT16), .ZN(new_n198));
  INV_X1    g012(.A(G125), .ZN(new_n199));
  NOR3_X1   g013(.A1(new_n199), .A2(KEYINPUT16), .A3(G140), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(G146), .B1(new_n198), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  AOI211_X1 g017(.A(new_n203), .B(new_n200), .C1(KEYINPUT16), .C2(new_n197), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n196), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  OAI22_X1  g019(.A1(new_n193), .A2(G110), .B1(new_n194), .B2(new_n195), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n197), .A2(new_n203), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n198), .A2(G146), .A3(new_n201), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT74), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT74), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n205), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G953), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(G221), .A3(G234), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n215), .B(KEYINPUT22), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n216), .B(G137), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n211), .A2(new_n213), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n210), .A2(KEYINPUT74), .A3(new_n217), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G902), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT25), .ZN(new_n224));
  XOR2_X1   g038(.A(KEYINPUT72), .B(G217), .Z(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n226), .B1(G234), .B2(new_n222), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT25), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n221), .A2(new_n228), .A3(new_n222), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n224), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n227), .A2(G902), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n221), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  XOR2_X1   g047(.A(KEYINPUT71), .B(KEYINPUT32), .Z(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  XOR2_X1   g049(.A(KEYINPUT2), .B(G113), .Z(new_n236));
  XNOR2_X1  g050(.A(G116), .B(G119), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n189), .A2(G116), .ZN(new_n239));
  INV_X1    g053(.A(G116), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT2), .B(G113), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n238), .A2(KEYINPUT66), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT66), .B1(new_n238), .B2(new_n244), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT30), .ZN(new_n248));
  NAND2_X1  g062(.A1(G134), .A2(G137), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT65), .B(G137), .ZN(new_n250));
  OAI211_X1 g064(.A(G131), .B(new_n249), .C1(new_n250), .C2(G134), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT11), .ZN(new_n252));
  INV_X1    g066(.A(G134), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(KEYINPUT11), .A2(G134), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G137), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n254), .B(new_n256), .C1(new_n250), .C2(new_n255), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n251), .B1(new_n257), .B2(G131), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(G143), .B(G146), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n187), .A2(new_n203), .A3(G143), .ZN(new_n264));
  INV_X1    g078(.A(G143), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n265), .B(G146), .C1(new_n187), .C2(KEYINPUT1), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n263), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n255), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(G137), .ZN(new_n270));
  INV_X1    g084(.A(G137), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(KEYINPUT65), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n268), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G131), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n273), .A2(new_n274), .A3(new_n254), .A4(new_n256), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(KEYINPUT67), .A3(new_n251), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n260), .A2(new_n267), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n261), .A2(KEYINPUT0), .A3(G128), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT0), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(new_n187), .A3(KEYINPUT64), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT64), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n281), .B1(KEYINPUT0), .B2(G128), .ZN(new_n282));
  NAND2_X1  g096(.A1(KEYINPUT0), .A2(G128), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n278), .B1(new_n261), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n257), .A2(G131), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n285), .B1(new_n286), .B2(new_n275), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n248), .B1(new_n277), .B2(new_n288), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n275), .A2(new_n267), .A3(new_n251), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n287), .A2(new_n290), .A3(KEYINPUT30), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n247), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n247), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n277), .A2(new_n293), .A3(new_n288), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n295), .B(G101), .ZN(new_n296));
  NOR2_X1   g110(.A1(G237), .A2(G953), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G210), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n296), .B(new_n298), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT31), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n292), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT68), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT68), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n292), .A2(new_n300), .A3(new_n304), .A4(new_n301), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n301), .B1(new_n292), .B2(new_n300), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n247), .B1(new_n287), .B2(new_n290), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT69), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT69), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n247), .B(new_n310), .C1(new_n287), .C2(new_n290), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n294), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT28), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT28), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n294), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n299), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n307), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n306), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(G472), .A2(G902), .ZN(new_n320));
  AOI21_X1  g134(.A(KEYINPUT70), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT70), .ZN(new_n322));
  INV_X1    g136(.A(new_n320), .ZN(new_n323));
  AOI211_X1 g137(.A(new_n322), .B(new_n323), .C1(new_n306), .C2(new_n318), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n235), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n317), .B1(new_n313), .B2(new_n315), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n292), .A2(new_n294), .A3(new_n317), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n277), .A2(new_n288), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n247), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n294), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT28), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n333), .A2(new_n315), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n317), .A2(new_n326), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n329), .A2(new_n336), .A3(new_n222), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n323), .B1(new_n306), .B2(new_n318), .ZN(new_n338));
  AOI22_X1  g152(.A1(G472), .A2(new_n337), .B1(new_n338), .B2(KEYINPUT32), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n233), .B1(new_n325), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n341));
  INV_X1    g155(.A(G104), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT75), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT75), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G104), .ZN(new_n345));
  INV_X1    g159(.A(G107), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT3), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n345), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G107), .ZN(new_n350));
  XOR2_X1   g164(.A(KEYINPUT76), .B(G101), .Z(new_n351));
  NOR3_X1   g165(.A1(new_n342), .A2(KEYINPUT3), .A3(G107), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n348), .A2(new_n350), .A3(new_n351), .A4(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G101), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n352), .B1(new_n347), .B2(KEYINPUT3), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n356), .B1(new_n357), .B2(new_n350), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT4), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n355), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n348), .A2(new_n350), .A3(new_n353), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n359), .A3(G101), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n238), .A2(KEYINPUT66), .A3(new_n244), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n238), .A2(new_n244), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT66), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n362), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n341), .B1(new_n360), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n239), .A2(KEYINPUT5), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n369), .B1(new_n237), .B2(KEYINPUT5), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n370), .A2(G113), .B1(new_n237), .B2(new_n236), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n347), .B1(G104), .B2(new_n346), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G101), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n354), .A2(new_n373), .A3(KEYINPUT78), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(KEYINPUT78), .B1(new_n354), .B2(new_n373), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n371), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n361), .A2(G101), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(KEYINPUT4), .A3(new_n354), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n379), .A2(KEYINPUT80), .A3(new_n247), .A4(new_n362), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n368), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  XOR2_X1   g195(.A(G110), .B(G122), .Z(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n382), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n368), .A2(new_n384), .A3(new_n377), .A4(new_n380), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(KEYINPUT6), .A3(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n267), .A2(G125), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n387), .B1(G125), .B2(new_n285), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n214), .A2(G224), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n388), .B(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT6), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n381), .A2(new_n391), .A3(new_n382), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n386), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n388), .A2(KEYINPUT7), .A3(new_n389), .ZN(new_n394));
  XOR2_X1   g208(.A(new_n394), .B(KEYINPUT81), .Z(new_n395));
  NOR2_X1   g209(.A1(new_n388), .A2(new_n389), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n354), .A2(new_n373), .ZN(new_n397));
  XOR2_X1   g211(.A(new_n397), .B(new_n371), .Z(new_n398));
  XOR2_X1   g212(.A(new_n382), .B(KEYINPUT8), .Z(new_n399));
  AOI21_X1  g213(.A(new_n396), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n388), .A2(KEYINPUT7), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n395), .A2(new_n385), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n393), .A2(new_n222), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(G210), .B1(G237), .B2(G902), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(KEYINPUT82), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n405), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n393), .A2(new_n222), .A3(new_n407), .A4(new_n402), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n204), .A2(new_n202), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n297), .A2(G143), .A3(G214), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(G143), .B1(new_n297), .B2(G214), .ZN(new_n413));
  OAI21_X1  g227(.A(G131), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT17), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT84), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n297), .A2(G214), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n265), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(new_n274), .A3(new_n411), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n414), .A2(new_n419), .A3(new_n415), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n274), .B1(new_n418), .B2(new_n411), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT84), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n422), .A3(KEYINPUT17), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n410), .A2(new_n416), .A3(new_n420), .A4(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n197), .B(new_n203), .ZN(new_n425));
  NAND2_X1  g239(.A1(KEYINPUT18), .A2(G131), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n418), .A2(new_n411), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT18), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n425), .B(new_n427), .C1(new_n428), .C2(new_n414), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(G113), .B(G122), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(new_n342), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(KEYINPUT85), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n424), .A2(new_n429), .A3(new_n433), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n222), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT86), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n435), .A2(KEYINPUT86), .A3(new_n222), .A4(new_n436), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(G475), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT19), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n197), .A2(new_n442), .ZN(new_n443));
  OR2_X1    g257(.A1(G125), .A2(G140), .ZN(new_n444));
  NAND2_X1  g258(.A1(G125), .A2(G140), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(KEYINPUT19), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n443), .A2(new_n203), .A3(new_n446), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n412), .A2(new_n413), .A3(G131), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n208), .B(new_n447), .C1(new_n448), .C2(new_n421), .ZN(new_n449));
  INV_X1    g263(.A(new_n432), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n429), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(new_n430), .B2(new_n432), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT20), .ZN(new_n453));
  INV_X1    g267(.A(G475), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n452), .A2(new_n453), .A3(new_n454), .A4(new_n222), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n450), .B1(new_n424), .B2(new_n429), .ZN(new_n456));
  NOR4_X1   g270(.A1(new_n456), .A2(new_n451), .A3(G475), .A4(G902), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n455), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n441), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G478), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(KEYINPUT15), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n240), .A2(G122), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n240), .A2(G122), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n465), .B1(KEYINPUT14), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n467), .B(KEYINPUT87), .C1(KEYINPUT14), .C2(new_n466), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n468), .B(G107), .C1(KEYINPUT87), .C2(new_n467), .ZN(new_n469));
  INV_X1    g283(.A(new_n465), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n470), .A2(new_n466), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n346), .ZN(new_n472));
  XNOR2_X1  g286(.A(G128), .B(G143), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(new_n253), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n469), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n471), .B(new_n346), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n473), .A2(KEYINPUT13), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n265), .A2(G128), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n477), .B(G134), .C1(KEYINPUT13), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n473), .A2(new_n253), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n476), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  XOR2_X1   g296(.A(KEYINPUT9), .B(G234), .Z(new_n483));
  NAND3_X1  g297(.A1(new_n225), .A2(new_n483), .A3(new_n214), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n484), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n475), .A2(new_n481), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n464), .B1(new_n488), .B2(new_n222), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n222), .A3(new_n464), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n461), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G952), .ZN(new_n494));
  AOI211_X1 g308(.A(G953), .B(new_n494), .C1(G234), .C2(G237), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AOI211_X1 g310(.A(new_n222), .B(new_n214), .C1(G234), .C2(G237), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  XOR2_X1   g312(.A(KEYINPUT21), .B(G898), .Z(new_n499));
  OAI21_X1  g313(.A(new_n496), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n500), .B(KEYINPUT88), .Z(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(G214), .B1(G237), .B2(G902), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n409), .A2(new_n493), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n483), .A2(new_n222), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n507), .A2(G221), .ZN(new_n508));
  INV_X1    g322(.A(G469), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(new_n222), .ZN(new_n510));
  XNOR2_X1  g324(.A(G110), .B(G140), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n214), .A2(G227), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n511), .B(new_n512), .Z(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n285), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n379), .A2(new_n515), .A3(new_n362), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT77), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT77), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n379), .A2(new_n518), .A3(new_n515), .A4(new_n362), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n286), .A2(new_n275), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n267), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n397), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT10), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT78), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n397), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n523), .B1(new_n528), .B2(new_n374), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n526), .B1(new_n529), .B2(new_n525), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n520), .A2(new_n522), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n522), .B1(new_n520), .B2(new_n530), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n514), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n520), .A2(new_n522), .A3(new_n530), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n267), .B1(new_n354), .B2(new_n373), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n521), .B1(new_n524), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT12), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n534), .A2(new_n540), .A3(new_n513), .ZN(new_n541));
  AOI21_X1  g355(.A(G902), .B1(new_n533), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n510), .B1(new_n542), .B2(new_n509), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n534), .A2(new_n513), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT79), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n520), .A2(new_n530), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n521), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT79), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n534), .A2(new_n548), .A3(new_n513), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n545), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n513), .B1(new_n534), .B2(new_n540), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(G469), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n508), .B1(new_n543), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n340), .A2(new_n506), .A3(new_n554), .ZN(new_n555));
  XOR2_X1   g369(.A(new_n555), .B(new_n351), .Z(G3));
  INV_X1    g370(.A(G472), .ZN(new_n557));
  AOI21_X1  g371(.A(G902), .B1(new_n306), .B2(new_n318), .ZN(new_n558));
  OAI22_X1  g372(.A1(new_n321), .A2(new_n324), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n508), .ZN(new_n560));
  INV_X1    g374(.A(new_n510), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n513), .B1(new_n547), .B2(new_n534), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n534), .A2(new_n540), .A3(new_n513), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n222), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n561), .B1(new_n564), .B2(G469), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n532), .B1(new_n544), .B2(KEYINPUT79), .ZN(new_n566));
  AOI211_X1 g380(.A(new_n509), .B(new_n551), .C1(new_n566), .C2(new_n549), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n560), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n559), .A2(new_n568), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n230), .A2(new_n232), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n403), .A2(new_n404), .ZN(new_n571));
  INV_X1    g385(.A(new_n404), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n393), .A2(new_n222), .A3(new_n572), .A4(new_n402), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n571), .A2(new_n503), .A3(new_n501), .A4(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n488), .A2(KEYINPUT33), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n485), .A2(new_n576), .A3(new_n487), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n577), .A3(G478), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n488), .A2(new_n462), .A3(new_n222), .ZN(new_n579));
  NAND2_X1  g393(.A1(G478), .A2(G902), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n461), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n574), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n569), .A2(new_n570), .A3(new_n583), .ZN(new_n584));
  XOR2_X1   g398(.A(KEYINPUT34), .B(G104), .Z(new_n585));
  XNOR2_X1  g399(.A(new_n584), .B(new_n585), .ZN(G6));
  NAND3_X1  g400(.A1(new_n452), .A2(new_n454), .A3(new_n222), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n458), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n457), .A2(new_n459), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n589), .A3(KEYINPUT89), .ZN(new_n590));
  OR3_X1    g404(.A1(new_n587), .A2(KEYINPUT89), .A3(new_n458), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n492), .A2(new_n590), .A3(new_n591), .A4(new_n441), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n574), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n569), .A2(new_n570), .A3(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT35), .B(G107), .Z(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(G9));
  AOI21_X1  g410(.A(new_n228), .B1(new_n221), .B2(new_n222), .ZN(new_n597));
  AOI211_X1 g411(.A(KEYINPUT25), .B(G902), .C1(new_n219), .C2(new_n220), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n218), .A2(KEYINPUT36), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(new_n210), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n599), .A2(new_n227), .B1(new_n231), .B2(new_n601), .ZN(new_n602));
  AOI211_X1 g416(.A(new_n508), .B(new_n602), .C1(new_n543), .C2(new_n553), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n319), .A2(new_n320), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n322), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n338), .A2(KEYINPUT70), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n319), .A2(new_n222), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n605), .A2(new_n606), .B1(G472), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n603), .A2(new_n506), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(new_n609), .B(KEYINPUT37), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(G110), .ZN(G12));
  OR2_X1    g425(.A1(new_n498), .A2(G900), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n496), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n592), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT90), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n325), .A2(new_n339), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n571), .A2(new_n503), .A3(new_n573), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n616), .A2(new_n617), .A3(new_n619), .A4(new_n603), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G128), .ZN(G30));
  XOR2_X1   g435(.A(KEYINPUT91), .B(KEYINPUT38), .Z(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT92), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n406), .A2(new_n624), .A3(new_n408), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n624), .B1(new_n406), .B2(new_n408), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n409), .A2(KEYINPUT92), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n629), .A2(new_n622), .A3(new_n625), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n504), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT93), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n317), .B1(new_n292), .B2(new_n294), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n332), .A2(new_n299), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n222), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n634), .A2(new_n635), .A3(new_n633), .ZN(new_n638));
  OAI21_X1  g452(.A(G472), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n338), .A2(KEYINPUT32), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n325), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n461), .A2(new_n492), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n613), .B(KEYINPUT94), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT39), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n554), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT95), .B(KEYINPUT40), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n632), .A2(new_n602), .A3(new_n644), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT96), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G143), .ZN(G45));
  NAND3_X1  g466(.A1(new_n581), .A2(new_n461), .A3(new_n613), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT97), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n617), .A2(new_n603), .A3(new_n619), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G146), .ZN(G48));
  NAND2_X1  g470(.A1(KEYINPUT98), .A2(G469), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n564), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n542), .A2(new_n657), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n660), .A3(new_n560), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n617), .A2(new_n570), .A3(new_n583), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT99), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT99), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n340), .A2(new_n665), .A3(new_n583), .A4(new_n662), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT41), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G113), .ZN(G15));
  NAND4_X1  g483(.A1(new_n617), .A2(new_n593), .A3(new_n570), .A4(new_n662), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G116), .ZN(G18));
  AOI21_X1  g485(.A(new_n234), .B1(new_n605), .B2(new_n606), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n337), .A2(G472), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n640), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n493), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n602), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n662), .A2(new_n619), .A3(new_n501), .A4(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(KEYINPUT100), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n493), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n679), .B1(new_n325), .B2(new_n339), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT100), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n661), .A2(new_n618), .A3(new_n602), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n680), .A2(new_n681), .A3(new_n682), .A4(new_n501), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G119), .ZN(G21));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n643), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n461), .A2(new_n492), .A3(KEYINPUT103), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n661), .A2(new_n618), .A3(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT101), .B(G472), .Z(new_n692));
  NAND2_X1  g506(.A1(new_n333), .A2(new_n315), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n317), .ZN(new_n694));
  INV_X1    g508(.A(new_n307), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n306), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n607), .A2(new_n692), .B1(new_n320), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n691), .B1(new_n697), .B2(new_n570), .ZN(new_n698));
  INV_X1    g512(.A(new_n692), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n558), .A2(new_n699), .ZN(new_n700));
  AOI22_X1  g514(.A1(new_n303), .A2(new_n305), .B1(new_n693), .B2(new_n317), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n323), .B1(new_n701), .B2(new_n695), .ZN(new_n702));
  NOR4_X1   g516(.A1(new_n700), .A2(new_n702), .A3(KEYINPUT102), .A4(new_n233), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n690), .B(new_n501), .C1(new_n698), .C2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G122), .ZN(G24));
  NAND3_X1  g519(.A1(new_n682), .A2(new_n654), .A3(new_n697), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G125), .ZN(G27));
  NOR2_X1   g521(.A1(new_n338), .A2(KEYINPUT32), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n570), .B1(new_n674), .B2(new_n708), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n709), .A2(KEYINPUT106), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(KEYINPUT106), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n560), .A2(new_n503), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n409), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n534), .A2(new_n540), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n715), .B1(new_n716), .B2(new_n513), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n551), .A2(KEYINPUT104), .ZN(new_n718));
  AOI22_X1  g532(.A1(new_n717), .A2(new_n718), .B1(new_n566), .B2(new_n549), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(G469), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n543), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n654), .A2(new_n714), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n712), .A2(KEYINPUT42), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n617), .A2(new_n570), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n654), .A2(new_n714), .A3(new_n721), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT105), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n722), .A2(new_n727), .A3(new_n340), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT42), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n723), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G131), .ZN(G33));
  NAND4_X1  g546(.A1(new_n340), .A2(new_n616), .A3(new_n721), .A4(new_n714), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G134), .ZN(G36));
  INV_X1    g548(.A(new_n461), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n581), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT108), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n736), .B(KEYINPUT43), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n739), .A2(new_n742), .A3(new_n559), .A4(new_n676), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT109), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n509), .B1(new_n719), .B2(KEYINPUT45), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n550), .A2(new_n552), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n510), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n748), .B1(new_n753), .B2(KEYINPUT46), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n564), .A2(G469), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n755), .B1(new_n753), .B2(KEYINPUT46), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n551), .A2(KEYINPUT104), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n551), .A2(KEYINPUT104), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n550), .B(KEYINPUT45), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n752), .A2(G469), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n561), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT46), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(KEYINPUT107), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n754), .A2(new_n756), .A3(new_n763), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n764), .A2(new_n560), .A3(new_n646), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n409), .A2(new_n504), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n743), .A2(new_n744), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n747), .A2(new_n765), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G137), .ZN(G39));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n770), .A2(KEYINPUT47), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(new_n764), .B2(new_n560), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n617), .ZN(new_n774));
  XNOR2_X1  g588(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n764), .A2(new_n560), .A3(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n654), .A2(new_n766), .A3(new_n233), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n773), .A2(new_n774), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  AND3_X1   g594(.A1(new_n631), .A2(new_n735), .A3(new_n581), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n642), .A2(new_n570), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n659), .A2(new_n660), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n713), .B1(new_n784), .B2(KEYINPUT49), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n784), .A2(KEYINPUT49), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n781), .A2(new_n783), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT111), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n704), .A2(new_n670), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(new_n666), .B2(new_n664), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n788), .B1(new_n790), .B2(new_n684), .ZN(new_n791));
  AOI211_X1 g605(.A(new_n233), .B(new_n661), .C1(new_n325), .C2(new_n339), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n696), .A2(new_n320), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n570), .B(new_n793), .C1(new_n558), .C2(new_n699), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT102), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n607), .A2(new_n692), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(new_n691), .A3(new_n570), .A4(new_n793), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n502), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  AOI22_X1  g612(.A1(new_n593), .A2(new_n792), .B1(new_n798), .B2(new_n690), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n788), .A2(new_n667), .A3(new_n684), .A4(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n608), .A2(new_n554), .A3(new_n570), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n409), .A2(new_n505), .ZN(new_n802));
  OR3_X1    g616(.A1(new_n801), .A2(new_n802), .A3(new_n582), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT112), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n492), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n490), .A2(KEYINPUT112), .A3(new_n491), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n461), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n409), .A2(new_n505), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT113), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n409), .A2(new_n811), .A3(new_n505), .A4(new_n808), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n804), .B(new_n609), .C1(new_n813), .C2(new_n801), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n569), .A2(new_n570), .A3(new_n810), .A4(new_n812), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n804), .B1(new_n816), .B2(new_n609), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n555), .B(new_n803), .C1(new_n815), .C2(new_n817), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n791), .A2(new_n800), .A3(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n700), .A2(new_n602), .A3(new_n702), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n722), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n590), .A2(new_n591), .ZN(new_n822));
  AND4_X1   g636(.A1(new_n441), .A2(new_n807), .A3(new_n613), .A4(new_n806), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n617), .A2(new_n603), .A3(new_n766), .A4(new_n823), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n821), .B(new_n733), .C1(new_n822), .C2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n641), .A2(new_n560), .A3(new_n602), .A4(new_n613), .ZN(new_n826));
  INV_X1    g640(.A(new_n689), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n721), .A2(new_n619), .A3(new_n827), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n620), .A2(new_n655), .A3(new_n706), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n830), .A3(KEYINPUT52), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n826), .A2(new_n828), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n620), .A2(new_n655), .A3(new_n706), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI221_X4 g649(.A(new_n825), .B1(new_n723), .B2(new_n730), .C1(new_n831), .C2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT53), .B1(new_n819), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n831), .A2(new_n835), .ZN(new_n838));
  INV_X1    g652(.A(new_n825), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n731), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n790), .A2(new_n788), .A3(new_n684), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n667), .A2(new_n799), .A3(new_n684), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT111), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n555), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n816), .A2(new_n609), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT114), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n845), .B1(new_n847), .B2(new_n814), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(KEYINPUT53), .A3(new_n803), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n840), .A2(new_n844), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT54), .B1(new_n837), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT115), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n841), .A2(new_n843), .A3(new_n803), .A4(new_n848), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(new_n854), .B2(new_n840), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n842), .B(KEYINPUT116), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n818), .A2(new_n853), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n836), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n855), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n861), .B(KEYINPUT54), .C1(new_n837), .C2(new_n850), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n852), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n659), .A2(new_n660), .A3(new_n508), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n764), .A2(new_n560), .A3(new_n776), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n865), .B1(new_n866), .B2(new_n772), .ZN(new_n867));
  AOI211_X1 g681(.A(new_n496), .B(new_n740), .C1(new_n795), .C2(new_n797), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n867), .A2(new_n766), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n766), .A2(new_n662), .A3(new_n495), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n782), .A2(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n871), .A2(new_n461), .A3(new_n581), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n628), .A2(new_n630), .A3(new_n504), .A4(new_n662), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n873), .A2(KEYINPUT117), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(KEYINPUT117), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n874), .A2(new_n868), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT50), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n874), .A2(KEYINPUT50), .A3(new_n868), .A4(new_n875), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n872), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n870), .A2(new_n740), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n820), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT118), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n869), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT119), .ZN(new_n886));
  INV_X1    g700(.A(new_n766), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT107), .B1(new_n761), .B2(new_n762), .ZN(new_n888));
  AOI211_X1 g702(.A(new_n748), .B(KEYINPUT46), .C1(new_n760), .C2(new_n561), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n508), .B1(new_n890), .B2(new_n756), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n777), .B1(new_n891), .B2(new_n771), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n887), .B1(new_n892), .B2(new_n865), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n886), .B1(new_n893), .B2(new_n868), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n885), .B1(new_n894), .B2(KEYINPUT51), .ZN(new_n895));
  AOI211_X1 g709(.A(new_n883), .B(new_n872), .C1(new_n878), .C2(new_n879), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT51), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n896), .A2(new_n886), .A3(new_n897), .A4(new_n869), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n712), .A2(new_n881), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT48), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n871), .A2(new_n582), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n661), .A2(new_n618), .ZN(new_n903));
  AOI211_X1 g717(.A(new_n494), .B(G953), .C1(new_n868), .C2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n864), .B1(new_n899), .B2(new_n906), .ZN(new_n907));
  AOI211_X1 g721(.A(KEYINPUT120), .B(new_n905), .C1(new_n895), .C2(new_n898), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n863), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(G952), .A2(G953), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n787), .B1(new_n909), .B2(new_n910), .ZN(G75));
  NAND2_X1  g725(.A1(new_n386), .A2(new_n392), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(new_n390), .ZN(new_n913));
  XNOR2_X1  g727(.A(KEYINPUT121), .B(KEYINPUT55), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n913), .B(new_n914), .Z(new_n915));
  INV_X1    g729(.A(G210), .ZN(new_n916));
  AOI211_X1 g730(.A(new_n916), .B(new_n222), .C1(new_n855), .C2(new_n858), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n917), .B2(KEYINPUT56), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n222), .B1(new_n855), .B2(new_n858), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(G210), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT56), .ZN(new_n921));
  INV_X1    g735(.A(new_n915), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n214), .A2(G952), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n918), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n918), .A2(new_n923), .A3(KEYINPUT122), .A4(new_n925), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(G51));
  NAND2_X1  g744(.A1(new_n561), .A2(KEYINPUT57), .ZN(new_n931));
  INV_X1    g745(.A(new_n860), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n859), .B1(new_n855), .B2(new_n858), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n561), .A2(KEYINPUT57), .ZN(new_n935));
  OAI22_X1  g749(.A1(new_n934), .A2(new_n935), .B1(new_n562), .B2(new_n563), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n919), .A2(new_n752), .A3(new_n749), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n924), .B1(new_n936), .B2(new_n937), .ZN(G54));
  NAND3_X1  g752(.A1(new_n919), .A2(KEYINPUT58), .A3(G475), .ZN(new_n939));
  INV_X1    g753(.A(new_n452), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n941), .A2(new_n942), .A3(new_n924), .ZN(G60));
  NAND2_X1  g757(.A1(new_n575), .A2(new_n577), .ZN(new_n944));
  XNOR2_X1  g758(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(new_n580), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n944), .B1(new_n863), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n932), .A2(new_n933), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n944), .A2(new_n946), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n947), .A2(new_n924), .A3(new_n950), .ZN(G63));
  NAND2_X1  g765(.A1(new_n855), .A2(new_n858), .ZN(new_n952));
  NAND2_X1  g766(.A1(G217), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT60), .Z(new_n954));
  NAND3_X1  g768(.A1(new_n952), .A2(new_n601), .A3(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n952), .A2(new_n954), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n925), .B(new_n955), .C1(new_n956), .C2(new_n221), .ZN(new_n957));
  AOI21_X1  g771(.A(KEYINPUT61), .B1(new_n955), .B2(KEYINPUT124), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(G66));
  AOI21_X1  g773(.A(new_n214), .B1(new_n499), .B2(G224), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n854), .B2(new_n214), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n912), .B1(G898), .B2(new_n214), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n961), .B(new_n962), .Z(G69));
  NAND2_X1  g777(.A1(new_n330), .A2(KEYINPUT30), .ZN(new_n964));
  INV_X1    g778(.A(new_n291), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n443), .A2(new_n446), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n619), .A2(new_n827), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(new_n710), .B2(new_n711), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n891), .A2(new_n646), .A3(new_n971), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n972), .A2(new_n731), .A3(new_n830), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n973), .A2(new_n768), .A3(new_n733), .A4(new_n779), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n214), .A2(G900), .ZN(new_n976));
  AOI22_X1  g790(.A1(new_n974), .A2(new_n214), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(KEYINPUT125), .B1(new_n214), .B2(G900), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n977), .A2(KEYINPUT126), .A3(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(KEYINPUT126), .B1(new_n977), .B2(new_n978), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n969), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n214), .B1(G227), .B2(G900), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n650), .A2(new_n830), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT62), .Z(new_n986));
  AOI21_X1  g800(.A(new_n808), .B1(new_n461), .B2(new_n581), .ZN(new_n987));
  OR4_X1    g801(.A1(new_n724), .A2(new_n647), .A3(new_n887), .A4(new_n987), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n986), .A2(new_n768), .A3(new_n779), .A4(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n969), .B1(new_n989), .B2(new_n214), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n982), .A2(new_n984), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n974), .A2(new_n214), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n976), .A2(new_n975), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n993), .A2(new_n978), .A3(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT126), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n968), .B1(new_n997), .B2(new_n979), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n983), .B1(new_n998), .B2(new_n990), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n992), .A2(new_n999), .ZN(G72));
  NOR2_X1   g814(.A1(new_n328), .A2(new_n634), .ZN(new_n1001));
  NAND2_X1  g815(.A1(G472), .A2(G902), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT63), .Z(new_n1003));
  OAI211_X1 g817(.A(new_n1001), .B(new_n1003), .C1(new_n837), .C2(new_n850), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT127), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1003), .B1(new_n974), .B2(new_n854), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(new_n328), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1003), .B1(new_n989), .B2(new_n854), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n924), .B1(new_n1008), .B2(new_n634), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n1005), .A2(new_n1007), .A3(new_n1009), .ZN(G57));
endmodule


