

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767;

  NOR2_X1 U374 ( .A1(n717), .A2(n716), .ZN(n726) );
  NAND2_X1 U375 ( .A1(n628), .A2(n627), .ZN(n629) );
  AND2_X1 U376 ( .A1(n558), .A2(n553), .ZN(n554) );
  NAND2_X1 U377 ( .A1(n652), .A2(n573), .ZN(n357) );
  XNOR2_X1 U378 ( .A(n416), .B(n415), .ZN(n763) );
  BUF_X1 U379 ( .A(n611), .Z(n356) );
  XNOR2_X1 U380 ( .A(n541), .B(KEYINPUT22), .ZN(n572) );
  AND2_X1 U381 ( .A1(n688), .A2(n427), .ZN(n365) );
  NOR2_X1 U382 ( .A1(G902), .A2(n737), .ZN(n489) );
  INV_X1 U383 ( .A(G953), .ZN(n458) );
  XNOR2_X1 U384 ( .A(n525), .B(n451), .ZN(n752) );
  XNOR2_X1 U385 ( .A(n446), .B(n509), .ZN(n739) );
  XNOR2_X1 U386 ( .A(n515), .B(n431), .ZN(n754) );
  BUF_X1 U387 ( .A(G146), .Z(n353) );
  XOR2_X1 U388 ( .A(KEYINPUT68), .B(G131), .Z(n516) );
  XOR2_X1 U389 ( .A(G122), .B(G107), .Z(n534) );
  INV_X1 U390 ( .A(G128), .ZN(n467) );
  XNOR2_X2 U391 ( .A(n513), .B(KEYINPUT33), .ZN(n720) );
  NAND2_X1 U392 ( .A1(n355), .A2(n354), .ZN(n387) );
  INV_X1 U393 ( .A(n550), .ZN(n354) );
  INV_X1 U394 ( .A(n551), .ZN(n355) );
  AND2_X2 U395 ( .A1(n379), .A2(n378), .ZN(n377) );
  XNOR2_X2 U396 ( .A(n495), .B(n494), .ZN(n525) );
  XNOR2_X2 U397 ( .A(n563), .B(KEYINPUT103), .ZN(n605) );
  XNOR2_X2 U398 ( .A(n677), .B(n626), .ZN(n755) );
  XNOR2_X1 U399 ( .A(n357), .B(KEYINPUT101), .ZN(n575) );
  XNOR2_X2 U400 ( .A(n449), .B(n448), .ZN(n766) );
  XNOR2_X2 U401 ( .A(KEYINPUT32), .B(n549), .ZN(n764) );
  AND2_X1 U402 ( .A1(n616), .A2(n372), .ZN(n371) );
  NOR2_X2 U403 ( .A1(n766), .A2(n767), .ZN(n410) );
  XNOR2_X1 U404 ( .A(n370), .B(n369), .ZN(n368) );
  NAND2_X1 U405 ( .A1(n371), .A2(n617), .ZN(n370) );
  NOR2_X2 U406 ( .A1(n764), .A2(n765), .ZN(n558) );
  XNOR2_X1 U407 ( .A(n462), .B(n461), .ZN(n509) );
  INV_X1 U408 ( .A(KEYINPUT0), .ZN(n440) );
  NOR2_X1 U409 ( .A1(n641), .A2(n738), .ZN(n643) );
  NOR2_X1 U410 ( .A1(n647), .A2(n738), .ZN(n650) );
  NOR2_X1 U411 ( .A1(n636), .A2(n738), .ZN(n637) );
  BUF_X1 U412 ( .A(n731), .Z(n735) );
  NAND2_X1 U413 ( .A1(n359), .A2(n368), .ZN(n677) );
  OR2_X1 U414 ( .A1(n623), .A2(n624), .ZN(n372) );
  OR2_X1 U415 ( .A1(n561), .A2(n514), .ZN(n436) );
  NOR2_X1 U416 ( .A1(n367), .A2(n702), .ZN(n612) );
  XNOR2_X1 U417 ( .A(n568), .B(KEYINPUT99), .ZN(n665) );
  NAND2_X1 U418 ( .A1(n395), .A2(n567), .ZN(n568) );
  NAND2_X2 U419 ( .A1(n377), .A2(n373), .ZN(n563) );
  XNOR2_X1 U420 ( .A(n418), .B(n360), .ZN(n567) );
  XNOR2_X1 U421 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U422 ( .A(n538), .B(n537), .ZN(n570) );
  XNOR2_X1 U423 ( .A(n406), .B(n533), .ZN(n733) );
  NAND2_X1 U424 ( .A1(n477), .A2(n580), .ZN(n442) );
  XNOR2_X1 U425 ( .A(n466), .B(G125), .ZN(n380) );
  XNOR2_X1 U426 ( .A(n394), .B(G104), .ZN(n522) );
  INV_X1 U427 ( .A(G113), .ZN(n394) );
  XOR2_X1 U428 ( .A(KEYINPUT4), .B(G101), .Z(n493) );
  INV_X1 U429 ( .A(G146), .ZN(n466) );
  BUF_X1 U430 ( .A(n700), .Z(n358) );
  XNOR2_X1 U431 ( .A(n619), .B(KEYINPUT38), .ZN(n700) );
  XNOR2_X2 U432 ( .A(n511), .B(n510), .ZN(n638) );
  XNOR2_X2 U433 ( .A(n752), .B(n496), .ZN(n511) );
  AND2_X1 U434 ( .A1(n457), .A2(n610), .ZN(n401) );
  OR2_X1 U435 ( .A1(G237), .A2(G902), .ZN(n471) );
  INV_X1 U436 ( .A(n675), .ZN(n407) );
  XNOR2_X1 U437 ( .A(n597), .B(n505), .ZN(n684) );
  XNOR2_X1 U438 ( .A(n409), .B(n408), .ZN(n702) );
  INV_X1 U439 ( .A(KEYINPUT100), .ZN(n408) );
  XNOR2_X1 U440 ( .A(n411), .B(n508), .ZN(n510) );
  XNOR2_X1 U441 ( .A(n509), .B(n364), .ZN(n411) );
  XNOR2_X1 U442 ( .A(n393), .B(n361), .ZN(n446) );
  XNOR2_X1 U443 ( .A(n534), .B(n522), .ZN(n393) );
  XOR2_X1 U444 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n486) );
  XNOR2_X1 U445 ( .A(n404), .B(n518), .ZN(n644) );
  XNOR2_X1 U446 ( .A(n524), .B(n517), .ZN(n404) );
  NOR2_X1 U447 ( .A1(n434), .A2(n435), .ZN(n433) );
  NOR2_X1 U448 ( .A1(n720), .A2(n514), .ZN(n434) );
  INV_X1 U449 ( .A(n609), .ZN(n438) );
  INV_X1 U450 ( .A(KEYINPUT82), .ZN(n419) );
  NOR2_X1 U451 ( .A1(n665), .A2(n661), .ZN(n703) );
  NAND2_X1 U452 ( .A1(n401), .A2(n402), .ZN(n399) );
  XNOR2_X1 U453 ( .A(n453), .B(KEYINPUT74), .ZN(n452) );
  INV_X1 U454 ( .A(G472), .ZN(n453) );
  XOR2_X1 U455 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n464) );
  XNOR2_X1 U456 ( .A(n380), .B(n392), .ZN(n391) );
  INV_X1 U457 ( .A(KEYINPUT78), .ZN(n392) );
  XNOR2_X1 U458 ( .A(n403), .B(KEYINPUT110), .ZN(n367) );
  XNOR2_X1 U459 ( .A(n425), .B(KEYINPUT70), .ZN(n594) );
  INV_X1 U460 ( .A(G902), .ZN(n375) );
  NAND2_X1 U461 ( .A1(n452), .A2(G902), .ZN(n378) );
  XNOR2_X1 U462 ( .A(n535), .B(KEYINPUT97), .ZN(n536) );
  XNOR2_X1 U463 ( .A(G116), .B(KEYINPUT95), .ZN(n526) );
  XOR2_X1 U464 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n527) );
  INV_X1 U465 ( .A(KEYINPUT43), .ZN(n414) );
  INV_X1 U466 ( .A(n684), .ZN(n624) );
  INV_X1 U467 ( .A(KEYINPUT105), .ZN(n439) );
  XNOR2_X1 U468 ( .A(n473), .B(n472), .ZN(n474) );
  OR2_X1 U469 ( .A1(n644), .A2(G902), .ZN(n418) );
  XNOR2_X1 U470 ( .A(n565), .B(KEYINPUT91), .ZN(n561) );
  BUF_X1 U471 ( .A(n684), .Z(n412) );
  NAND2_X1 U472 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U473 ( .A(n754), .B(n428), .ZN(n488) );
  XNOR2_X1 U474 ( .A(n430), .B(n429), .ZN(n428) );
  NOR2_X1 U475 ( .A1(n756), .A2(G952), .ZN(n738) );
  INV_X1 U476 ( .A(KEYINPUT40), .ZN(n448) );
  AND2_X1 U477 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U478 ( .A1(G953), .A2(G237), .ZN(n519) );
  INV_X1 U479 ( .A(KEYINPUT12), .ZN(n397) );
  XOR2_X1 U480 ( .A(G140), .B(KEYINPUT11), .Z(n521) );
  INV_X1 U481 ( .A(KEYINPUT48), .ZN(n369) );
  XNOR2_X1 U482 ( .A(n400), .B(KEYINPUT20), .ZN(n490) );
  NAND2_X1 U483 ( .A1(n478), .A2(G234), .ZN(n400) );
  XOR2_X1 U484 ( .A(KEYINPUT5), .B(KEYINPUT77), .Z(n507) );
  XNOR2_X1 U485 ( .A(G137), .B(G113), .ZN(n506) );
  INV_X1 U486 ( .A(KEYINPUT10), .ZN(n481) );
  XNOR2_X1 U487 ( .A(n516), .B(KEYINPUT69), .ZN(n451) );
  XNOR2_X1 U488 ( .A(n421), .B(G140), .ZN(n497) );
  INV_X1 U489 ( .A(G137), .ZN(n421) );
  XNOR2_X1 U490 ( .A(n470), .B(KEYINPUT89), .ZN(n627) );
  XNOR2_X1 U491 ( .A(G902), .B(KEYINPUT15), .ZN(n470) );
  AND2_X1 U492 ( .A1(n684), .A2(n365), .ZN(n564) );
  XNOR2_X1 U493 ( .A(n503), .B(n504), .ZN(n597) );
  NOR2_X1 U494 ( .A1(G902), .A2(n730), .ZN(n503) );
  INV_X1 U495 ( .A(KEYINPUT45), .ZN(n384) );
  NAND2_X1 U496 ( .A1(n387), .A2(KEYINPUT44), .ZN(n386) );
  XNOR2_X1 U497 ( .A(n484), .B(n483), .ZN(n430) );
  XNOR2_X1 U498 ( .A(n482), .B(KEYINPUT93), .ZN(n429) );
  XNOR2_X1 U499 ( .A(G119), .B(KEYINPUT24), .ZN(n482) );
  INV_X1 U500 ( .A(n497), .ZN(n431) );
  XNOR2_X1 U501 ( .A(n497), .B(n420), .ZN(n499) );
  INV_X1 U502 ( .A(G110), .ZN(n420) );
  XNOR2_X1 U503 ( .A(n739), .B(n447), .ZN(n631) );
  NAND2_X1 U504 ( .A1(G234), .A2(G237), .ZN(n460) );
  INV_X1 U505 ( .A(KEYINPUT19), .ZN(n443) );
  BUF_X1 U506 ( .A(n597), .Z(n405) );
  XNOR2_X1 U507 ( .A(n596), .B(n595), .ZN(n424) );
  NAND2_X1 U508 ( .A1(n376), .A2(n375), .ZN(n374) );
  XNOR2_X1 U509 ( .A(n532), .B(n536), .ZN(n406) );
  XOR2_X1 U510 ( .A(n644), .B(KEYINPUT59), .Z(n646) );
  XNOR2_X1 U511 ( .A(n589), .B(n413), .ZN(n590) );
  XNOR2_X1 U512 ( .A(n414), .B(KEYINPUT108), .ZN(n413) );
  XNOR2_X1 U513 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U514 ( .A(n620), .B(KEYINPUT36), .ZN(n621) );
  INV_X1 U515 ( .A(KEYINPUT35), .ZN(n415) );
  INV_X1 U516 ( .A(n570), .ZN(n395) );
  NOR2_X1 U517 ( .A1(n608), .A2(n609), .ZN(n664) );
  AND2_X1 U518 ( .A1(n424), .A2(n422), .ZN(n600) );
  NOR2_X1 U519 ( .A1(n417), .A2(n423), .ZN(n422) );
  INV_X1 U520 ( .A(n405), .ZN(n423) );
  BUF_X1 U521 ( .A(n598), .Z(n417) );
  NAND2_X1 U522 ( .A1(n444), .A2(n688), .ZN(n652) );
  XNOR2_X1 U523 ( .A(n445), .B(KEYINPUT86), .ZN(n444) );
  NOR2_X1 U524 ( .A1(n572), .A2(n366), .ZN(n445) );
  INV_X1 U525 ( .A(n738), .ZN(n388) );
  XNOR2_X1 U526 ( .A(n456), .B(n455), .ZN(n454) );
  XNOR2_X1 U527 ( .A(n730), .B(n729), .ZN(n455) );
  INV_X1 U528 ( .A(n582), .ZN(n427) );
  NOR2_X1 U529 ( .A1(n676), .A2(n407), .ZN(n359) );
  XOR2_X1 U530 ( .A(KEYINPUT13), .B(G475), .Z(n360) );
  XNOR2_X1 U531 ( .A(G110), .B(KEYINPUT16), .ZN(n361) );
  AND2_X1 U532 ( .A1(n559), .A2(n556), .ZN(n362) );
  XOR2_X1 U533 ( .A(n480), .B(n479), .Z(n363) );
  AND2_X1 U534 ( .A1(n519), .A2(G210), .ZN(n364) );
  OR2_X1 U535 ( .A1(n583), .A2(n412), .ZN(n366) );
  NOR2_X1 U536 ( .A1(n367), .A2(n703), .ZN(n704) );
  INV_X1 U537 ( .A(n372), .ZN(n673) );
  OR2_X1 U538 ( .A1(n638), .A2(n374), .ZN(n373) );
  INV_X1 U539 ( .A(n452), .ZN(n376) );
  NAND2_X1 U540 ( .A1(n638), .A2(n452), .ZN(n379) );
  NAND2_X1 U541 ( .A1(n605), .A2(n699), .ZN(n398) );
  XNOR2_X1 U542 ( .A(n380), .B(n481), .ZN(n515) );
  NAND2_X1 U543 ( .A1(n381), .A2(n386), .ZN(n385) );
  NOR2_X1 U544 ( .A1(n383), .A2(n382), .ZN(n381) );
  NAND2_X1 U545 ( .A1(n575), .A2(n560), .ZN(n382) );
  NAND2_X1 U546 ( .A1(n557), .A2(n362), .ZN(n383) );
  XNOR2_X2 U547 ( .A(n385), .B(n384), .ZN(n746) );
  AND2_X1 U548 ( .A1(n389), .A2(n388), .ZN(G66) );
  XNOR2_X1 U549 ( .A(n736), .B(n390), .ZN(n389) );
  INV_X1 U550 ( .A(n737), .ZN(n390) );
  XNOR2_X1 U551 ( .A(n398), .B(KEYINPUT30), .ZN(n606) );
  XNOR2_X1 U552 ( .A(n645), .B(n646), .ZN(n647) );
  XNOR2_X1 U553 ( .A(n564), .B(n439), .ZN(n512) );
  XNOR2_X1 U554 ( .A(n639), .B(n640), .ZN(n641) );
  XNOR2_X1 U555 ( .A(n493), .B(n495), .ZN(n468) );
  XNOR2_X1 U556 ( .A(n476), .B(n443), .ZN(n598) );
  XNOR2_X1 U557 ( .A(n468), .B(n391), .ZN(n469) );
  NOR2_X2 U558 ( .A1(n606), .A2(n607), .ZN(n615) );
  INV_X1 U559 ( .A(n567), .ZN(n569) );
  XNOR2_X1 U560 ( .A(n523), .B(n396), .ZN(n524) );
  XNOR2_X1 U561 ( .A(n522), .B(n397), .ZN(n396) );
  XNOR2_X1 U562 ( .A(n399), .B(KEYINPUT75), .ZN(n617) );
  NOR2_X2 U563 ( .A1(n598), .A2(n442), .ZN(n441) );
  NAND2_X1 U564 ( .A1(n611), .A2(n699), .ZN(n476) );
  XNOR2_X2 U565 ( .A(n475), .B(n474), .ZN(n611) );
  NOR2_X1 U566 ( .A1(n763), .A2(KEYINPUT87), .ZN(n551) );
  XNOR2_X1 U567 ( .A(n664), .B(KEYINPUT83), .ZN(n457) );
  NAND2_X1 U568 ( .A1(n599), .A2(n600), .ZN(n402) );
  NOR2_X1 U569 ( .A1(n697), .A2(n613), .ZN(n614) );
  NAND2_X1 U570 ( .A1(n700), .A2(n699), .ZN(n403) );
  XNOR2_X1 U571 ( .A(n511), .B(n502), .ZN(n730) );
  NOR2_X1 U572 ( .A1(n558), .A2(KEYINPUT65), .ZN(n550) );
  NOR2_X1 U573 ( .A1(n570), .A2(n567), .ZN(n409) );
  XNOR2_X1 U574 ( .A(n410), .B(KEYINPUT46), .ZN(n616) );
  XNOR2_X1 U575 ( .A(n528), .B(KEYINPUT98), .ZN(n529) );
  XNOR2_X1 U576 ( .A(n469), .B(n465), .ZN(n447) );
  NAND2_X1 U577 ( .A1(n433), .A2(n432), .ZN(n416) );
  NAND2_X1 U578 ( .A1(n436), .A2(n438), .ZN(n435) );
  XNOR2_X1 U579 ( .A(n703), .B(n419), .ZN(n592) );
  NOR2_X2 U580 ( .A1(n755), .A2(n746), .ZN(n678) );
  NAND2_X1 U581 ( .A1(n600), .A2(n601), .ZN(n602) );
  NAND2_X1 U582 ( .A1(n424), .A2(n405), .ZN(n613) );
  NOR2_X1 U583 ( .A1(n688), .A2(n426), .ZN(n425) );
  NAND2_X1 U584 ( .A1(n427), .A2(n603), .ZN(n426) );
  NAND2_X1 U585 ( .A1(n720), .A2(n437), .ZN(n432) );
  AND2_X1 U586 ( .A1(n561), .A2(n514), .ZN(n437) );
  XNOR2_X2 U587 ( .A(n489), .B(n363), .ZN(n688) );
  XNOR2_X2 U588 ( .A(n441), .B(n440), .ZN(n565) );
  NAND2_X1 U589 ( .A1(n625), .A2(n665), .ZN(n449) );
  XNOR2_X2 U590 ( .A(n450), .B(KEYINPUT39), .ZN(n625) );
  NAND2_X1 U591 ( .A1(n615), .A2(n358), .ZN(n450) );
  XNOR2_X2 U592 ( .A(n467), .B(G143), .ZN(n495) );
  NOR2_X1 U593 ( .A1(n454), .A2(n738), .ZN(G54) );
  NAND2_X1 U594 ( .A1(n735), .A2(G469), .ZN(n456) );
  XNOR2_X1 U595 ( .A(n635), .B(n634), .ZN(n636) );
  INV_X1 U596 ( .A(G134), .ZN(n494) );
  XNOR2_X1 U597 ( .A(KEYINPUT109), .B(KEYINPUT28), .ZN(n595) );
  XNOR2_X1 U598 ( .A(n530), .B(n529), .ZN(n533) );
  INV_X1 U599 ( .A(KEYINPUT90), .ZN(n472) );
  INV_X1 U600 ( .A(KEYINPUT60), .ZN(n648) );
  INV_X1 U601 ( .A(KEYINPUT63), .ZN(n642) );
  XNOR2_X1 U602 ( .A(n648), .B(KEYINPUT123), .ZN(n649) );
  INV_X1 U603 ( .A(KEYINPUT44), .ZN(n553) );
  XNOR2_X1 U604 ( .A(KEYINPUT34), .B(KEYINPUT79), .ZN(n514) );
  NOR2_X1 U605 ( .A1(G898), .A2(n458), .ZN(n741) );
  NAND2_X1 U606 ( .A1(n741), .A2(G902), .ZN(n459) );
  NAND2_X1 U607 ( .A1(G952), .A2(n458), .ZN(n577) );
  NAND2_X1 U608 ( .A1(n459), .A2(n577), .ZN(n477) );
  XNOR2_X1 U609 ( .A(n460), .B(KEYINPUT14), .ZN(n580) );
  INV_X1 U610 ( .A(n580), .ZN(n715) );
  NAND2_X1 U611 ( .A1(G214), .A2(n471), .ZN(n699) );
  XOR2_X1 U612 ( .A(G116), .B(G119), .Z(n462) );
  XNOR2_X1 U613 ( .A(KEYINPUT3), .B(KEYINPUT73), .ZN(n461) );
  XOR2_X2 U614 ( .A(KEYINPUT64), .B(G953), .Z(n756) );
  NAND2_X1 U615 ( .A1(G224), .A2(n756), .ZN(n463) );
  XNOR2_X1 U616 ( .A(n464), .B(n463), .ZN(n465) );
  INV_X1 U617 ( .A(n627), .ZN(n478) );
  NAND2_X1 U618 ( .A1(n631), .A2(n478), .ZN(n475) );
  NAND2_X1 U619 ( .A1(G210), .A2(n471), .ZN(n473) );
  XOR2_X1 U620 ( .A(KEYINPUT25), .B(KEYINPUT94), .Z(n480) );
  NAND2_X1 U621 ( .A1(n490), .A2(G217), .ZN(n479) );
  XOR2_X1 U622 ( .A(KEYINPUT23), .B(KEYINPUT92), .Z(n483) );
  XNOR2_X1 U623 ( .A(G128), .B(G110), .ZN(n484) );
  NAND2_X1 U624 ( .A1(G234), .A2(n756), .ZN(n485) );
  XNOR2_X1 U625 ( .A(n486), .B(n485), .ZN(n531) );
  NAND2_X1 U626 ( .A1(G221), .A2(n531), .ZN(n487) );
  XNOR2_X1 U627 ( .A(n488), .B(n487), .ZN(n737) );
  NAND2_X1 U628 ( .A1(n490), .A2(G221), .ZN(n491) );
  XNOR2_X1 U629 ( .A(n491), .B(KEYINPUT21), .ZN(n582) );
  XNOR2_X1 U630 ( .A(G469), .B(KEYINPUT71), .ZN(n492) );
  XNOR2_X1 U631 ( .A(n492), .B(KEYINPUT72), .ZN(n504) );
  XNOR2_X1 U632 ( .A(n353), .B(n493), .ZN(n496) );
  NAND2_X1 U633 ( .A1(G227), .A2(n756), .ZN(n501) );
  XNOR2_X1 U634 ( .A(G107), .B(G104), .ZN(n498) );
  XNOR2_X1 U635 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U636 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U637 ( .A(KEYINPUT1), .B(KEYINPUT66), .ZN(n505) );
  XNOR2_X1 U638 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U639 ( .A(n563), .B(KEYINPUT6), .Z(n546) );
  INV_X1 U640 ( .A(n546), .ZN(n583) );
  NAND2_X1 U641 ( .A1(n512), .A2(n583), .ZN(n513) );
  XOR2_X1 U642 ( .A(n515), .B(G122), .Z(n518) );
  XNOR2_X1 U643 ( .A(n516), .B(G143), .ZN(n517) );
  NAND2_X1 U644 ( .A1(G214), .A2(n519), .ZN(n520) );
  XNOR2_X1 U645 ( .A(n521), .B(n520), .ZN(n523) );
  XNOR2_X1 U646 ( .A(n525), .B(KEYINPUT96), .ZN(n530) );
  XOR2_X1 U647 ( .A(n527), .B(n526), .Z(n528) );
  NAND2_X1 U648 ( .A1(G217), .A2(n531), .ZN(n532) );
  INV_X1 U649 ( .A(n534), .ZN(n535) );
  NOR2_X1 U650 ( .A1(n733), .A2(G902), .ZN(n538) );
  INV_X1 U651 ( .A(G478), .ZN(n537) );
  NAND2_X1 U652 ( .A1(n567), .A2(n570), .ZN(n609) );
  INV_X1 U653 ( .A(n565), .ZN(n540) );
  NOR2_X1 U654 ( .A1(n582), .A2(n702), .ZN(n539) );
  OR2_X1 U655 ( .A1(n688), .A2(n605), .ZN(n542) );
  OR2_X1 U656 ( .A1(n412), .A2(n542), .ZN(n543) );
  NOR2_X1 U657 ( .A1(n572), .A2(n543), .ZN(n544) );
  XNOR2_X1 U658 ( .A(n544), .B(KEYINPUT104), .ZN(n765) );
  NOR2_X1 U659 ( .A1(n624), .A2(n688), .ZN(n545) );
  XNOR2_X1 U660 ( .A(KEYINPUT102), .B(n545), .ZN(n547) );
  NAND2_X1 U661 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U662 ( .A1(n572), .A2(n548), .ZN(n549) );
  NAND2_X1 U663 ( .A1(n763), .A2(n554), .ZN(n557) );
  NOR2_X1 U664 ( .A1(KEYINPUT87), .A2(KEYINPUT65), .ZN(n555) );
  OR2_X1 U665 ( .A1(KEYINPUT44), .A2(n555), .ZN(n556) );
  NAND2_X1 U666 ( .A1(KEYINPUT87), .A2(n763), .ZN(n560) );
  NAND2_X1 U667 ( .A1(n558), .A2(KEYINPUT65), .ZN(n559) );
  AND2_X1 U668 ( .A1(n405), .A2(n365), .ZN(n604) );
  AND2_X1 U669 ( .A1(n561), .A2(n604), .ZN(n562) );
  NAND2_X1 U670 ( .A1(n563), .A2(n562), .ZN(n655) );
  INV_X1 U671 ( .A(n563), .ZN(n687) );
  NAND2_X1 U672 ( .A1(n564), .A2(n687), .ZN(n693) );
  NOR2_X1 U673 ( .A1(n565), .A2(n693), .ZN(n566) );
  XNOR2_X1 U674 ( .A(KEYINPUT31), .B(n566), .ZN(n670) );
  NAND2_X1 U675 ( .A1(n655), .A2(n670), .ZN(n571) );
  NAND2_X1 U676 ( .A1(n570), .A2(n569), .ZN(n671) );
  INV_X1 U677 ( .A(n671), .ZN(n661) );
  NAND2_X1 U678 ( .A1(n571), .A2(n592), .ZN(n573) );
  NOR2_X1 U679 ( .A1(n756), .A2(G900), .ZN(n576) );
  NAND2_X1 U680 ( .A1(G902), .A2(n576), .ZN(n578) );
  NAND2_X1 U681 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U682 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U683 ( .A(KEYINPUT80), .B(n581), .Z(n603) );
  AND2_X1 U684 ( .A1(n665), .A2(n583), .ZN(n584) );
  NAND2_X1 U685 ( .A1(n594), .A2(n584), .ZN(n586) );
  INV_X1 U686 ( .A(KEYINPUT106), .ZN(n585) );
  XNOR2_X1 U687 ( .A(n586), .B(n585), .ZN(n587) );
  NAND2_X1 U688 ( .A1(n587), .A2(n699), .ZN(n618) );
  XNOR2_X1 U689 ( .A(n618), .B(KEYINPUT107), .ZN(n588) );
  NAND2_X1 U690 ( .A1(n588), .A2(n624), .ZN(n589) );
  NOR2_X1 U691 ( .A1(n356), .A2(n590), .ZN(n676) );
  XNOR2_X1 U692 ( .A(KEYINPUT47), .B(KEYINPUT67), .ZN(n591) );
  XNOR2_X1 U693 ( .A(n593), .B(KEYINPUT76), .ZN(n599) );
  NAND2_X1 U694 ( .A1(n605), .A2(n594), .ZN(n596) );
  INV_X1 U695 ( .A(n703), .ZN(n601) );
  NAND2_X1 U696 ( .A1(n602), .A2(KEYINPUT47), .ZN(n610) );
  NAND2_X1 U697 ( .A1(n604), .A2(n603), .ZN(n607) );
  NAND2_X1 U698 ( .A1(n615), .A2(n356), .ZN(n608) );
  INV_X1 U699 ( .A(n611), .ZN(n619) );
  XNOR2_X1 U700 ( .A(n612), .B(KEYINPUT41), .ZN(n697) );
  XNOR2_X1 U701 ( .A(n614), .B(KEYINPUT42), .ZN(n767) );
  NOR2_X1 U702 ( .A1(n619), .A2(n618), .ZN(n622) );
  INV_X1 U703 ( .A(KEYINPUT88), .ZN(n620) );
  NAND2_X1 U704 ( .A1(n625), .A2(n661), .ZN(n675) );
  INV_X1 U705 ( .A(KEYINPUT85), .ZN(n626) );
  NOR2_X2 U706 ( .A1(n678), .A2(KEYINPUT2), .ZN(n630) );
  NOR2_X1 U707 ( .A1(n677), .A2(n746), .ZN(n680) );
  NAND2_X1 U708 ( .A1(n680), .A2(KEYINPUT2), .ZN(n628) );
  NOR2_X4 U709 ( .A1(n630), .A2(n629), .ZN(n731) );
  NAND2_X1 U710 ( .A1(n731), .A2(G210), .ZN(n635) );
  INV_X1 U711 ( .A(n631), .ZN(n633) );
  XOR2_X1 U712 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n632) );
  XNOR2_X1 U713 ( .A(n637), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U714 ( .A(n638), .B(KEYINPUT62), .ZN(n640) );
  NAND2_X1 U715 ( .A1(n731), .A2(G472), .ZN(n639) );
  XNOR2_X1 U716 ( .A(n643), .B(n642), .ZN(G57) );
  NAND2_X1 U717 ( .A1(n731), .A2(G475), .ZN(n645) );
  XNOR2_X1 U718 ( .A(n650), .B(n649), .ZN(G60) );
  XOR2_X1 U719 ( .A(G101), .B(KEYINPUT111), .Z(n651) );
  XNOR2_X1 U720 ( .A(n652), .B(n651), .ZN(G3) );
  INV_X1 U721 ( .A(n665), .ZN(n667) );
  NOR2_X1 U722 ( .A1(n667), .A2(n655), .ZN(n653) );
  XOR2_X1 U723 ( .A(KEYINPUT112), .B(n653), .Z(n654) );
  XNOR2_X1 U724 ( .A(G104), .B(n654), .ZN(G6) );
  NOR2_X1 U725 ( .A1(n671), .A2(n655), .ZN(n660) );
  XOR2_X1 U726 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n657) );
  XNOR2_X1 U727 ( .A(G107), .B(KEYINPUT26), .ZN(n656) );
  XNOR2_X1 U728 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U729 ( .A(KEYINPUT27), .B(n658), .ZN(n659) );
  XNOR2_X1 U730 ( .A(n660), .B(n659), .ZN(G9) );
  XOR2_X1 U731 ( .A(G128), .B(KEYINPUT29), .Z(n663) );
  NAND2_X1 U732 ( .A1(n600), .A2(n661), .ZN(n662) );
  XNOR2_X1 U733 ( .A(n663), .B(n662), .ZN(G30) );
  XOR2_X1 U734 ( .A(n664), .B(G143), .Z(G45) );
  NAND2_X1 U735 ( .A1(n600), .A2(n665), .ZN(n666) );
  XNOR2_X1 U736 ( .A(n666), .B(n353), .ZN(G48) );
  NOR2_X1 U737 ( .A1(n667), .A2(n670), .ZN(n669) );
  XNOR2_X1 U738 ( .A(G113), .B(KEYINPUT115), .ZN(n668) );
  XNOR2_X1 U739 ( .A(n669), .B(n668), .ZN(G15) );
  NOR2_X1 U740 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U741 ( .A(G116), .B(n672), .Z(G18) );
  XNOR2_X1 U742 ( .A(G125), .B(n673), .ZN(n674) );
  XNOR2_X1 U743 ( .A(n674), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U744 ( .A(G134), .B(n675), .ZN(G36) );
  XOR2_X1 U745 ( .A(G140), .B(n676), .Z(G42) );
  INV_X1 U746 ( .A(KEYINPUT2), .ZN(n718) );
  OR2_X1 U747 ( .A1(n677), .A2(n718), .ZN(n679) );
  NAND2_X1 U748 ( .A1(n679), .A2(n678), .ZN(n683) );
  NOR2_X1 U749 ( .A1(n680), .A2(KEYINPUT81), .ZN(n681) );
  NAND2_X1 U750 ( .A1(n681), .A2(KEYINPUT2), .ZN(n682) );
  NAND2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n717) );
  NOR2_X1 U752 ( .A1(n365), .A2(n412), .ZN(n685) );
  XNOR2_X1 U753 ( .A(n685), .B(KEYINPUT50), .ZN(n686) );
  NOR2_X1 U754 ( .A1(n687), .A2(n686), .ZN(n692) );
  NOR2_X1 U755 ( .A1(n688), .A2(n427), .ZN(n690) );
  XNOR2_X1 U756 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n689) );
  XNOR2_X1 U757 ( .A(n690), .B(n689), .ZN(n691) );
  NAND2_X1 U758 ( .A1(n692), .A2(n691), .ZN(n694) );
  NAND2_X1 U759 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U760 ( .A(n695), .B(KEYINPUT51), .ZN(n696) );
  XNOR2_X1 U761 ( .A(n696), .B(KEYINPUT117), .ZN(n698) );
  INV_X1 U762 ( .A(n697), .ZN(n719) );
  NAND2_X1 U763 ( .A1(n698), .A2(n719), .ZN(n710) );
  NOR2_X1 U764 ( .A1(n358), .A2(n699), .ZN(n701) );
  NOR2_X1 U765 ( .A1(n702), .A2(n701), .ZN(n706) );
  XNOR2_X1 U766 ( .A(n704), .B(KEYINPUT118), .ZN(n705) );
  NOR2_X1 U767 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U768 ( .A(KEYINPUT119), .B(n707), .ZN(n708) );
  NAND2_X1 U769 ( .A1(n708), .A2(n720), .ZN(n709) );
  NAND2_X1 U770 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U771 ( .A(n711), .B(KEYINPUT120), .ZN(n712) );
  XNOR2_X1 U772 ( .A(n712), .B(KEYINPUT52), .ZN(n713) );
  NAND2_X1 U773 ( .A1(n713), .A2(G952), .ZN(n714) );
  NOR2_X1 U774 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U775 ( .A1(KEYINPUT81), .A2(n718), .ZN(n723) );
  AND2_X1 U776 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U777 ( .A(n721), .B(KEYINPUT121), .ZN(n722) );
  NAND2_X1 U778 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U779 ( .A1(n724), .A2(G953), .ZN(n725) );
  NAND2_X1 U780 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U781 ( .A(KEYINPUT122), .B(n727), .ZN(n728) );
  XOR2_X1 U782 ( .A(KEYINPUT53), .B(n728), .Z(G75) );
  XOR2_X1 U783 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n729) );
  NAND2_X1 U784 ( .A1(G478), .A2(n735), .ZN(n732) );
  XNOR2_X1 U785 ( .A(n733), .B(n732), .ZN(n734) );
  NOR2_X1 U786 ( .A1(n738), .A2(n734), .ZN(G63) );
  NAND2_X1 U787 ( .A1(G217), .A2(n735), .ZN(n736) );
  XOR2_X1 U788 ( .A(n739), .B(G101), .Z(n740) );
  XNOR2_X1 U789 ( .A(KEYINPUT125), .B(n740), .ZN(n742) );
  NOR2_X1 U790 ( .A1(n742), .A2(n741), .ZN(n750) );
  NAND2_X1 U791 ( .A1(G224), .A2(G953), .ZN(n743) );
  XNOR2_X1 U792 ( .A(n743), .B(KEYINPUT61), .ZN(n744) );
  XNOR2_X1 U793 ( .A(KEYINPUT124), .B(n744), .ZN(n745) );
  NAND2_X1 U794 ( .A1(G898), .A2(n745), .ZN(n748) );
  OR2_X1 U795 ( .A1(n746), .A2(G953), .ZN(n747) );
  NAND2_X1 U796 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U797 ( .A(n750), .B(n749), .ZN(n751) );
  XNOR2_X1 U798 ( .A(KEYINPUT126), .B(n751), .ZN(G69) );
  XOR2_X1 U799 ( .A(n752), .B(KEYINPUT4), .Z(n753) );
  XNOR2_X1 U800 ( .A(n754), .B(n753), .ZN(n758) );
  XNOR2_X1 U801 ( .A(n758), .B(n755), .ZN(n757) );
  NAND2_X1 U802 ( .A1(n757), .A2(n756), .ZN(n762) );
  XNOR2_X1 U803 ( .A(G227), .B(n758), .ZN(n759) );
  NAND2_X1 U804 ( .A1(n759), .A2(G900), .ZN(n760) );
  NAND2_X1 U805 ( .A1(G953), .A2(n760), .ZN(n761) );
  NAND2_X1 U806 ( .A1(n762), .A2(n761), .ZN(G72) );
  XNOR2_X1 U807 ( .A(n763), .B(G122), .ZN(G24) );
  XOR2_X1 U808 ( .A(G119), .B(n764), .Z(G21) );
  XOR2_X1 U809 ( .A(n765), .B(G110), .Z(G12) );
  XOR2_X1 U810 ( .A(n766), .B(G131), .Z(G33) );
  XOR2_X1 U811 ( .A(n767), .B(G137), .Z(G39) );
endmodule

