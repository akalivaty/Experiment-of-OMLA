//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001;
  NAND2_X1  g000(.A1(G71gat), .A2(G78gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(G71gat), .A2(G78gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT102), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(new_n204), .B2(new_n202), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT103), .ZN(new_n207));
  INV_X1    g006(.A(new_n202), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n208), .A2(KEYINPUT9), .ZN(new_n209));
  OR2_X1    g008(.A1(G57gat), .A2(G64gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G57gat), .A2(G64gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n207), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n208), .A2(new_n203), .ZN(new_n214));
  XOR2_X1   g013(.A(new_n214), .B(KEYINPUT105), .Z(new_n215));
  INV_X1    g014(.A(G57gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(KEYINPUT104), .ZN(new_n217));
  INV_X1    g016(.A(G64gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n215), .A2(new_n209), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n213), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT21), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G231gat), .A2(G233gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(G127gat), .B(G155gat), .Z(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(KEYINPUT106), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n227), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n231), .A2(G1gat), .ZN(new_n232));
  AOI21_X1  g031(.A(G8gat), .B1(new_n232), .B2(KEYINPUT100), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT16), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n231), .B1(new_n234), .B2(G1gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n233), .B(new_n236), .Z(new_n237));
  AND2_X1   g036(.A1(new_n213), .A2(new_n220), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n237), .B1(new_n238), .B2(KEYINPUT21), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n230), .A2(new_n239), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n227), .A2(new_n229), .ZN(new_n241));
  INV_X1    g040(.A(new_n239), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n229), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  XOR2_X1   g043(.A(G183gat), .B(G211gat), .Z(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n240), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n246), .B1(new_n240), .B2(new_n244), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(G43gat), .B(G50gat), .Z(new_n250));
  INV_X1    g049(.A(KEYINPUT15), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G43gat), .B(G50gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT15), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT14), .ZN(new_n255));
  INV_X1    g054(.A(G29gat), .ZN(new_n256));
  INV_X1    g055(.A(G36gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G29gat), .A2(G36gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT98), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n252), .A2(new_n254), .A3(new_n260), .A4(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT99), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n263), .A2(KEYINPUT99), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT96), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n260), .B(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n254), .B1(new_n267), .B2(new_n261), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT97), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n264), .A2(new_n265), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OR2_X1    g069(.A1(new_n268), .A2(new_n269), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(KEYINPUT17), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(G85gat), .A2(G92gat), .ZN(new_n275));
  MUX2_X1   g074(.A(KEYINPUT7), .B(new_n274), .S(new_n275), .Z(new_n276));
  INV_X1    g075(.A(G99gat), .ZN(new_n277));
  INV_X1    g076(.A(G106gat), .ZN(new_n278));
  OR3_X1    g077(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT107), .ZN(new_n279));
  OAI21_X1  g078(.A(KEYINPUT107), .B1(new_n277), .B2(new_n278), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n276), .B1(KEYINPUT8), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G99gat), .B(G106gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT108), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n282), .A2(KEYINPUT108), .A3(new_n283), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n282), .A2(new_n283), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n289), .ZN(new_n291));
  AND2_X1   g090(.A1(G232gat), .A2(G233gat), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n272), .A2(new_n291), .B1(KEYINPUT41), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(G190gat), .B(G218gat), .Z(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(KEYINPUT109), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n294), .B(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n292), .A2(KEYINPUT41), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n298), .ZN(new_n300));
  XOR2_X1   g099(.A(G134gat), .B(G162gat), .Z(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n300), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n297), .A2(new_n298), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G230gat), .ZN(new_n307));
  INV_X1    g106(.A(G233gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n238), .A2(new_n284), .A3(new_n288), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n310), .B1(new_n221), .B2(new_n289), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT10), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n291), .A2(new_n238), .A3(KEYINPUT10), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n309), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n309), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G120gat), .B(G148gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(G176gat), .B(G204gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  OR3_X1    g119(.A1(new_n315), .A2(new_n317), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n320), .B1(new_n315), .B2(new_n317), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(KEYINPUT110), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT110), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n324), .B(new_n320), .C1(new_n315), .C2(new_n317), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n249), .A2(new_n303), .A3(new_n306), .A4(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT111), .ZN(new_n328));
  INV_X1    g127(.A(new_n237), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n273), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n272), .A2(new_n237), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT101), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n273), .A2(KEYINPUT101), .A3(new_n329), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G229gat), .A2(G233gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(KEYINPUT18), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n333), .A2(new_n336), .A3(new_n334), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT18), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n272), .B(new_n237), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n336), .B(KEYINPUT13), .Z(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n337), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G113gat), .B(G141gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(KEYINPUT11), .ZN(new_n346));
  INV_X1    g145(.A(G169gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(G197gat), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n349), .B(KEYINPUT12), .Z(new_n350));
  NAND2_X1  g149(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n350), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n337), .A2(new_n340), .A3(new_n343), .A4(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n306), .A2(new_n303), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT111), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n355), .A2(new_n356), .A3(new_n249), .A4(new_n326), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n328), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G8gat), .B(G36gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT79), .ZN(new_n360));
  XOR2_X1   g159(.A(G64gat), .B(G92gat), .Z(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G226gat), .A2(G233gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(G183gat), .A2(G190gat), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT26), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT26), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n371), .B1(G169gat), .B2(G176gat), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n368), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G183gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT27), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT27), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(G183gat), .ZN(new_n377));
  INV_X1    g176(.A(G190gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n375), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT28), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT27), .B(G183gat), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(KEYINPUT28), .A3(new_n378), .ZN(new_n383));
  AOI211_X1 g182(.A(new_n366), .B(new_n373), .C1(new_n381), .C2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT69), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT68), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT24), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n365), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n374), .A2(new_n378), .ZN(new_n389));
  NAND3_X1  g188(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n392), .A2(new_n386), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n385), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n389), .A2(new_n390), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n365), .A2(new_n387), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT68), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n395), .A2(new_n397), .A3(KEYINPUT69), .A4(new_n388), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(G176gat), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n347), .A2(new_n400), .A3(KEYINPUT23), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n401), .A2(KEYINPUT25), .A3(new_n367), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT67), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(new_n369), .B2(KEYINPUT23), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT23), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n405), .B(KEYINPUT67), .C1(G169gat), .C2(G176gat), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n402), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n399), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT25), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n368), .B1(new_n404), .B2(new_n406), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n401), .A2(KEYINPUT66), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT66), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n369), .A2(new_n412), .A3(KEYINPUT23), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT64), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n390), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n389), .ZN(new_n418));
  NAND4_X1  g217(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n419), .B1(new_n392), .B2(KEYINPUT65), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n365), .A2(KEYINPUT65), .A3(new_n387), .ZN(new_n421));
  NOR3_X1   g220(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n409), .B1(new_n415), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n384), .B1(new_n408), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n364), .B1(new_n424), .B2(KEYINPUT29), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT65), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n396), .A2(new_n426), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n390), .A2(new_n416), .B1(new_n374), .B2(new_n378), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n392), .A2(KEYINPUT65), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n427), .A2(new_n428), .A3(new_n429), .A4(new_n419), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(new_n410), .A3(new_n414), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n399), .A2(new_n407), .B1(new_n431), .B2(new_n409), .ZN(new_n432));
  OAI211_X1 g231(.A(G226gat), .B(G233gat), .C1(new_n432), .C2(new_n384), .ZN(new_n433));
  INV_X1    g232(.A(G204gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(G197gat), .ZN(new_n435));
  INV_X1    g234(.A(G197gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(G204gat), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(new_n437), .A3(KEYINPUT75), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT75), .B1(new_n435), .B2(new_n437), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(G211gat), .ZN(new_n442));
  INV_X1    g241(.A(G218gat), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(G211gat), .A2(G218gat), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(KEYINPUT22), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT76), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT22), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n435), .A2(new_n437), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT75), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n449), .B1(new_n452), .B2(new_n438), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n444), .A2(new_n445), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n448), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT22), .B1(new_n439), .B2(new_n440), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(KEYINPUT76), .A3(new_n454), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n447), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n425), .A2(new_n433), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n447), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n453), .A2(new_n448), .A3(new_n455), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT76), .B1(new_n457), .B2(new_n454), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT77), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT77), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n425), .A2(new_n433), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n363), .B1(new_n460), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT81), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT30), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n425), .A2(new_n433), .A3(new_n459), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n408), .A2(new_n423), .ZN(new_n473));
  INV_X1    g272(.A(new_n384), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n364), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT29), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n476), .B1(new_n432), .B2(new_n384), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n475), .B1(new_n364), .B2(new_n477), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n465), .A2(new_n467), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n472), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT81), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(new_n363), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n470), .A2(new_n471), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT78), .B1(new_n460), .B2(new_n468), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT78), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n485), .B(new_n472), .C1(new_n478), .C2(new_n479), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n362), .B(KEYINPUT80), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n480), .A2(KEYINPUT30), .A3(new_n363), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n483), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  XOR2_X1   g289(.A(G127gat), .B(G134gat), .Z(new_n491));
  XNOR2_X1  g290(.A(G113gat), .B(G120gat), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n491), .B1(KEYINPUT1), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT70), .ZN(new_n494));
  INV_X1    g293(.A(G120gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(G113gat), .ZN(new_n496));
  INV_X1    g295(.A(G113gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(G120gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G127gat), .B(G134gat), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT1), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n493), .A2(new_n494), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n494), .B1(new_n493), .B2(new_n502), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(G148gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(G141gat), .ZN(new_n508));
  INV_X1    g307(.A(G141gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(G148gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(G155gat), .A2(G162gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT2), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(G155gat), .A2(G162gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT82), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n512), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(KEYINPUT82), .A2(G155gat), .A3(G162gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT83), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT83), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n518), .A2(new_n522), .A3(new_n519), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n515), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  XOR2_X1   g323(.A(KEYINPUT84), .B(G141gat), .Z(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(G148gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT2), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n516), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n526), .A2(new_n508), .B1(new_n512), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT4), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n506), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n493), .A2(new_n502), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n518), .A2(new_n522), .A3(new_n519), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n522), .B1(new_n518), .B2(new_n519), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n514), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n528), .A2(new_n512), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT84), .B(G141gat), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n539), .A2(new_n507), .ZN(new_n540));
  INV_X1    g339(.A(new_n508), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n534), .A2(new_n537), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT4), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n537), .A2(new_n542), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n534), .B1(new_n545), .B2(KEYINPUT3), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT3), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n537), .A2(new_n547), .A3(new_n542), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n532), .A2(new_n544), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT5), .ZN(new_n550));
  NAND2_X1  g349(.A1(G225gat), .A2(G233gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT3), .B1(new_n524), .B2(new_n529), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(new_n533), .A3(new_n548), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n551), .ZN(new_n555));
  NOR4_X1   g354(.A1(new_n524), .A2(new_n529), .A3(new_n533), .A4(KEYINPUT4), .ZN(new_n556));
  INV_X1    g355(.A(new_n502), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n500), .B1(new_n501), .B2(new_n499), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT70), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n503), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT4), .B1(new_n560), .B2(new_n545), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT85), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n556), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI211_X1 g362(.A(KEYINPUT85), .B(KEYINPUT4), .C1(new_n560), .C2(new_n545), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n555), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n545), .A2(new_n533), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n566), .A2(new_n543), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT5), .B1(new_n567), .B2(new_n551), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n552), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G1gat), .B(G29gat), .Z(new_n570));
  XNOR2_X1  g369(.A(G57gat), .B(G85gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n569), .A2(KEYINPUT6), .A3(new_n575), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n569), .A2(new_n575), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n552), .B(new_n574), .C1(new_n565), .C2(new_n568), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT87), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT6), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n580), .B1(new_n579), .B2(new_n581), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n578), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n490), .B1(new_n576), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G228gat), .A2(G233gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n548), .A2(new_n476), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n459), .ZN(new_n588));
  OR2_X1    g387(.A1(new_n461), .A2(KEYINPUT88), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n457), .A2(new_n454), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n461), .A2(KEYINPUT88), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT3), .B1(new_n592), .B2(new_n476), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n586), .B(new_n588), .C1(new_n593), .C2(new_n530), .ZN(new_n594));
  XNOR2_X1  g393(.A(G78gat), .B(G106gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT31), .B(G50gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(G22gat), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n547), .B1(new_n459), .B2(KEYINPUT29), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n479), .A2(new_n587), .B1(new_n545), .B2(new_n599), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n594), .B(new_n598), .C1(new_n600), .C2(new_n586), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n594), .B1(new_n600), .B2(new_n586), .ZN(new_n602));
  INV_X1    g401(.A(new_n598), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT73), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n506), .B1(new_n432), .B2(new_n384), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n473), .A2(new_n474), .A3(new_n560), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(G227gat), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n609), .A2(new_n308), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n605), .B(KEYINPUT34), .C1(new_n608), .C2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n610), .B1(new_n606), .B2(new_n607), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT34), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT73), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n611), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n606), .A2(new_n607), .A3(new_n610), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n617), .A2(KEYINPUT32), .ZN(new_n618));
  XOR2_X1   g417(.A(G15gat), .B(G43gat), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT71), .ZN(new_n620));
  XOR2_X1   g419(.A(G71gat), .B(G99gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT72), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT33), .ZN(new_n624));
  INV_X1    g423(.A(new_n622), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n625), .B1(new_n617), .B2(KEYINPUT32), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n617), .A2(new_n627), .ZN(new_n628));
  AOI22_X1  g427(.A1(new_n618), .A2(new_n624), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n616), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n618), .A2(new_n624), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n626), .A2(new_n628), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n611), .A2(new_n614), .A3(new_n615), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AND4_X1   g434(.A1(new_n601), .A2(new_n604), .A3(new_n630), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n585), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n579), .A2(new_n581), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n576), .B1(new_n577), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT35), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n604), .A2(new_n641), .A3(new_n601), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n640), .A2(new_n490), .A3(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n633), .A2(new_n634), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT74), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n645), .B1(new_n616), .B2(new_n629), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n633), .A2(KEYINPUT74), .A3(new_n634), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n637), .A2(KEYINPUT35), .B1(new_n643), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT89), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n604), .A2(new_n601), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n584), .A2(new_n576), .ZN(new_n653));
  INV_X1    g452(.A(new_n490), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n630), .A2(KEYINPUT36), .A3(new_n635), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n616), .A2(new_n629), .A3(new_n645), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT74), .B1(new_n633), .B2(new_n634), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n630), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT36), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n656), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n650), .B1(new_n655), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n630), .A2(new_n635), .A3(KEYINPUT36), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(new_n648), .B2(KEYINPUT36), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n664), .B(KEYINPUT89), .C1(new_n585), .C2(new_n652), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n484), .A2(KEYINPUT37), .A3(new_n486), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT94), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(new_n668), .A3(new_n362), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT93), .B(KEYINPUT37), .Z(new_n670));
  NAND2_X1  g469(.A1(new_n480), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n668), .B1(new_n667), .B2(new_n362), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT38), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT95), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g475(.A(KEYINPUT95), .B(KEYINPUT38), .C1(new_n672), .C2(new_n673), .ZN(new_n677));
  INV_X1    g476(.A(new_n487), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(KEYINPUT38), .ZN(new_n679));
  MUX2_X1   g478(.A(new_n464), .B(new_n479), .S(new_n478), .Z(new_n680));
  INV_X1    g479(.A(KEYINPUT37), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n671), .B(new_n679), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n470), .A2(new_n482), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n640), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n676), .A2(new_n677), .A3(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n549), .A2(new_n551), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT39), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n575), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n566), .A2(new_n543), .A3(new_n551), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT90), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n688), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  OAI221_X1 g491(.A(new_n692), .B1(new_n691), .B2(new_n690), .C1(new_n549), .C2(new_n551), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n689), .A2(KEYINPUT40), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT92), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n689), .A2(KEYINPUT92), .A3(new_n693), .A4(KEYINPUT40), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT91), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT40), .B1(new_n689), .B2(new_n693), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n577), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n700), .A2(new_n699), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n698), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n652), .B1(new_n703), .B2(new_n654), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n686), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n649), .B1(new_n666), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n358), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT112), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n653), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n584), .A2(KEYINPUT112), .A3(new_n576), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g515(.A1(new_n358), .A2(new_n490), .A3(new_n708), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n717), .A2(KEYINPUT113), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(KEYINPUT113), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n718), .A2(G8gat), .A3(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT16), .B(G8gat), .Z(new_n721));
  NAND4_X1  g520(.A1(new_n709), .A2(KEYINPUT42), .A3(new_n490), .A4(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT114), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n718), .A2(new_n719), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n721), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT42), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n723), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n721), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(new_n718), .B2(new_n719), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n729), .A2(KEYINPUT114), .A3(KEYINPUT42), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n720), .B(new_n722), .C1(new_n727), .C2(new_n730), .ZN(G1325gat));
  INV_X1    g530(.A(new_n709), .ZN(new_n732));
  OAI21_X1  g531(.A(G15gat), .B1(new_n732), .B2(new_n664), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n659), .A2(G15gat), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n732), .B2(new_n734), .ZN(G1326gat));
  NAND2_X1  g534(.A1(new_n709), .A2(new_n651), .ZN(new_n736));
  XNOR2_X1  g535(.A(KEYINPUT43), .B(G22gat), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1327gat));
  INV_X1    g537(.A(KEYINPUT115), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n739), .B(KEYINPUT44), .C1(new_n707), .C2(new_n355), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n637), .A2(KEYINPUT35), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n643), .A2(new_n648), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n684), .B1(new_n675), .B2(new_n674), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n704), .B1(new_n744), .B2(new_n677), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n664), .B1(new_n585), .B2(new_n652), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n743), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n306), .A2(new_n303), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n740), .A2(new_n750), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n662), .A2(new_n665), .B1(new_n686), .B2(new_n705), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n749), .B1(new_n752), .B2(new_n649), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n739), .B1(new_n753), .B2(KEYINPUT44), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n354), .ZN(new_n756));
  INV_X1    g555(.A(new_n326), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n756), .A2(new_n249), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n256), .B1(new_n760), .B2(new_n714), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n708), .A2(new_n749), .A3(new_n758), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n762), .A2(G29gat), .A3(new_n713), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT45), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n761), .A2(new_n764), .ZN(G1328gat));
  NAND2_X1  g564(.A1(new_n490), .A2(new_n257), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT116), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT46), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n257), .B1(new_n760), .B2(new_n490), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n769), .A2(new_n770), .ZN(G1329gat));
  NAND3_X1  g570(.A1(new_n760), .A2(G43gat), .A3(new_n661), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n762), .A2(new_n659), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(G43gat), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g574(.A1(new_n760), .A2(G50gat), .A3(new_n651), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n762), .A2(new_n652), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(G50gat), .B2(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g578(.A1(new_n240), .A2(new_n244), .A3(new_n246), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n240), .A2(new_n244), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n245), .ZN(new_n782));
  AND4_X1   g581(.A1(new_n780), .A2(new_n306), .A3(new_n782), .A4(new_n303), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n747), .A2(new_n783), .A3(new_n756), .A4(new_n757), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n714), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g586(.A(new_n654), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n789), .B(new_n790), .Z(G1333gat));
  OAI21_X1  g590(.A(G71gat), .B1(new_n784), .B2(new_n664), .ZN(new_n792));
  OR2_X1    g591(.A1(new_n659), .A2(G71gat), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n792), .B1(new_n784), .B2(new_n793), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n794), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g594(.A1(new_n785), .A2(new_n651), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G78gat), .ZN(G1335gat));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n746), .B1(new_n686), .B2(new_n705), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n799), .B(new_n749), .C1(new_n800), .C2(new_n649), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n249), .A2(new_n354), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n799), .B1(new_n747), .B2(new_n749), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n798), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n746), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n649), .B1(new_n706), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT117), .B1(new_n807), .B2(new_n355), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n808), .A2(KEYINPUT51), .A3(new_n801), .A4(new_n802), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n326), .B1(new_n805), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(G85gat), .B1(new_n810), .B2(new_n714), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n249), .A2(new_n354), .A3(new_n326), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n755), .A2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n714), .A2(G85gat), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n811), .B1(new_n814), .B2(new_n815), .ZN(G1336gat));
  NAND2_X1  g615(.A1(new_n805), .A2(new_n809), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(new_n490), .A3(new_n757), .ZN(new_n818));
  INV_X1    g617(.A(G92gat), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n654), .A2(new_n819), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n812), .B(new_n821), .C1(new_n751), .C2(new_n754), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n820), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(G92gat), .B1(new_n810), .B2(new_n490), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n822), .A2(new_n825), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT119), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n823), .A2(new_n824), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n828), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(new_n828), .B2(new_n831), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(G1337gat));
  AOI21_X1  g634(.A(G99gat), .B1(new_n810), .B2(new_n648), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n664), .A2(new_n277), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n814), .B2(new_n837), .ZN(G1338gat));
  NAND3_X1  g637(.A1(new_n814), .A2(G106gat), .A3(new_n651), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n810), .A2(new_n651), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(G106gat), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n841), .B(new_n842), .ZN(G1339gat));
  OAI21_X1  g642(.A(KEYINPUT120), .B1(new_n327), .B2(new_n354), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n783), .A2(new_n845), .A3(new_n756), .A4(new_n326), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n249), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n313), .A2(new_n314), .A3(new_n309), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n849), .A2(new_n315), .A3(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n320), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n853), .B1(new_n315), .B2(new_n850), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(KEYINPUT55), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT55), .ZN(new_n856));
  INV_X1    g655(.A(new_n854), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(new_n851), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n855), .A2(new_n321), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n354), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n335), .A2(new_n336), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n341), .A2(new_n342), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n349), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n353), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n757), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n749), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n749), .A2(new_n864), .A3(new_n859), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n848), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n847), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n713), .A2(new_n490), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n636), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(G113gat), .B1(new_n873), .B2(new_n354), .ZN(new_n874));
  INV_X1    g673(.A(new_n871), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n659), .A2(new_n651), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n756), .A2(new_n497), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n874), .B1(new_n878), .B2(new_n879), .ZN(G1340gat));
  AOI21_X1  g679(.A(G120gat), .B1(new_n873), .B2(new_n757), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n326), .A2(new_n495), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n878), .B2(new_n882), .ZN(G1341gat));
  OAI21_X1  g682(.A(G127gat), .B1(new_n877), .B2(new_n848), .ZN(new_n884));
  INV_X1    g683(.A(G127gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n873), .A2(new_n885), .A3(new_n249), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(G1342gat));
  OAI21_X1  g686(.A(G134gat), .B1(new_n877), .B2(new_n355), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n871), .A2(new_n355), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n872), .A2(G134gat), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT121), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n889), .A2(new_n893), .A3(new_n890), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n892), .A2(KEYINPUT56), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT56), .B1(new_n892), .B2(new_n894), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n888), .B1(new_n895), .B2(new_n896), .ZN(G1343gat));
  NOR2_X1   g696(.A1(new_n661), .A2(new_n652), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n869), .A2(new_n870), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n354), .A2(new_n509), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT122), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n713), .A2(new_n490), .A3(new_n661), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n869), .A2(KEYINPUT57), .A3(new_n651), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT57), .B1(new_n869), .B2(new_n651), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n354), .B(new_n902), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n901), .B1(new_n906), .B2(new_n539), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT58), .ZN(new_n908));
  INV_X1    g707(.A(new_n902), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT57), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n847), .A2(new_n868), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(new_n652), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n909), .B1(new_n912), .B2(new_n903), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n525), .B1(new_n913), .B2(new_n354), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n901), .A2(KEYINPUT58), .ZN(new_n915));
  OAI22_X1  g714(.A1(new_n907), .A2(new_n908), .B1(new_n914), .B2(new_n915), .ZN(G1344gat));
  INV_X1    g715(.A(new_n899), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(new_n507), .A3(new_n757), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n328), .A2(new_n756), .A3(new_n357), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n652), .B1(new_n920), .B2(new_n868), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n903), .B1(KEYINPUT57), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n757), .A3(new_n902), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n919), .B1(new_n923), .B2(G148gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n919), .A2(G148gat), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n925), .B1(new_n913), .B2(new_n757), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n918), .B1(new_n924), .B2(new_n926), .ZN(G1345gat));
  INV_X1    g726(.A(G155gat), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n917), .A2(new_n928), .A3(new_n249), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n913), .A2(new_n249), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n929), .B1(new_n930), .B2(new_n928), .ZN(G1346gat));
  INV_X1    g730(.A(G162gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n889), .A2(new_n932), .A3(new_n898), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n749), .B(new_n902), .C1(new_n904), .C2(new_n905), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(KEYINPUT123), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G162gat), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n934), .A2(KEYINPUT123), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(G1347gat));
  NOR2_X1   g737(.A1(new_n714), .A2(new_n654), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n939), .A2(new_n876), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n869), .A2(new_n940), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n941), .A2(new_n347), .A3(new_n756), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT124), .B1(new_n911), .B2(new_n714), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n869), .A2(new_n944), .A3(new_n713), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n654), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n946), .A2(new_n636), .A3(new_n354), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n942), .B1(new_n947), .B2(new_n347), .ZN(G1348gat));
  NAND4_X1  g747(.A1(new_n946), .A2(new_n400), .A3(new_n636), .A4(new_n757), .ZN(new_n949));
  OAI21_X1  g748(.A(G176gat), .B1(new_n941), .B2(new_n326), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1349gat));
  NAND2_X1  g750(.A1(new_n943), .A2(new_n945), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n249), .A2(new_n382), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n952), .A2(new_n490), .A3(new_n636), .A4(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(G183gat), .B1(new_n941), .B2(new_n848), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(KEYINPUT60), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT60), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n954), .A2(new_n958), .A3(new_n955), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(G1350gat));
  NOR2_X1   g759(.A1(new_n355), .A2(G190gat), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n952), .A2(new_n490), .A3(new_n636), .A4(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n869), .A2(new_n749), .A3(new_n940), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(G190gat), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(KEYINPUT61), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n963), .A2(new_n966), .A3(G190gat), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n962), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT125), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT125), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n962), .A2(new_n968), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(G1351gat));
  NOR2_X1   g772(.A1(new_n756), .A2(G197gat), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n946), .A2(new_n898), .A3(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n946), .A2(KEYINPUT126), .A3(new_n898), .A4(new_n974), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n939), .A2(new_n664), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n922), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g780(.A(G197gat), .B1(new_n981), .B2(new_n756), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n977), .A2(new_n978), .A3(new_n982), .ZN(G1352gat));
  NOR2_X1   g782(.A1(new_n326), .A2(G204gat), .ZN(new_n984));
  NAND4_X1  g783(.A1(new_n952), .A2(new_n490), .A3(new_n898), .A4(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n946), .A2(KEYINPUT62), .A3(new_n898), .A4(new_n984), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n990), .B1(new_n981), .B2(new_n326), .ZN(new_n991));
  NAND4_X1  g790(.A1(new_n922), .A2(KEYINPUT127), .A3(new_n757), .A4(new_n980), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n991), .A2(new_n992), .A3(G204gat), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n989), .A2(new_n993), .ZN(G1353gat));
  NAND4_X1  g793(.A1(new_n946), .A2(new_n442), .A3(new_n249), .A4(new_n898), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n922), .A2(new_n249), .A3(new_n980), .ZN(new_n996));
  AND3_X1   g795(.A1(new_n996), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n997));
  AOI21_X1  g796(.A(KEYINPUT63), .B1(new_n996), .B2(G211gat), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(G1354gat));
  OAI21_X1  g798(.A(G218gat), .B1(new_n981), .B2(new_n355), .ZN(new_n1000));
  NAND4_X1  g799(.A1(new_n946), .A2(new_n443), .A3(new_n749), .A4(new_n898), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(G1355gat));
endmodule


