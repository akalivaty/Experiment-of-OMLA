//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0008(.A1(new_n206), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G1), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n212), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT0), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n217), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n214), .B(new_n220), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND2_X1  g0046(.A1(G33), .A2(G87), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT79), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  AND2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  OAI211_X1 g0051(.A(G226), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  OAI211_X1 g0053(.A(G223), .B(new_n253), .C1(new_n250), .C2(new_n251), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n249), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G1), .A3(G13), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n215), .B1(G41), .B2(G45), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G274), .ZN(new_n263));
  INV_X1    g0063(.A(new_n211), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n263), .B1(new_n264), .B2(new_n256), .ZN(new_n265));
  INV_X1    g0065(.A(new_n260), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n262), .A2(G232), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G190), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n259), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n266), .A2(new_n257), .A3(G274), .ZN(new_n270));
  INV_X1    g0070(.A(G232), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n270), .B1(new_n271), .B2(new_n261), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n272), .B1(new_n258), .B2(new_n255), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n269), .B1(new_n273), .B2(G200), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT16), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT7), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT3), .B(G33), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n276), .B1(new_n277), .B2(G20), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n250), .A2(new_n251), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n202), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G58), .A2(G68), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n203), .A2(new_n205), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G20), .ZN(new_n284));
  INV_X1    g0084(.A(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n212), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G159), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n275), .B1(new_n281), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(KEYINPUT7), .B1(new_n279), .B2(new_n212), .ZN(new_n291));
  NOR4_X1   g0091(.A1(new_n250), .A2(new_n251), .A3(new_n276), .A4(G20), .ZN(new_n292));
  OAI21_X1  g0092(.A(G68), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n283), .A2(G20), .B1(G159), .B2(new_n287), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(KEYINPUT16), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n211), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n290), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT8), .B(G58), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n215), .A2(G13), .A3(G20), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  XOR2_X1   g0102(.A(KEYINPUT8), .B(G58), .Z(new_n303));
  NAND2_X1  g0103(.A1(new_n215), .A2(G20), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n300), .A2(new_n211), .A3(new_n296), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n302), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT78), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n307), .B(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n274), .A2(new_n298), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT17), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n310), .B(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n298), .A2(new_n309), .ZN(new_n313));
  AOI21_X1  g0113(.A(G169), .B1(new_n259), .B2(new_n267), .ZN(new_n314));
  INV_X1    g0114(.A(G179), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n314), .B1(new_n315), .B2(new_n273), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT18), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n313), .A2(KEYINPUT18), .A3(new_n316), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(KEYINPUT80), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT80), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n313), .A2(new_n316), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT18), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n312), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n202), .A2(G20), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n212), .A2(G33), .ZN(new_n326));
  INV_X1    g0126(.A(G77), .ZN(new_n327));
  INV_X1    g0127(.A(G50), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n325), .B1(new_n326), .B2(new_n327), .C1(new_n328), .C2(new_n286), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n297), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n330), .A2(KEYINPUT75), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(KEYINPUT75), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT11), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n330), .A2(KEYINPUT75), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT11), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n330), .A2(KEYINPUT75), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n215), .A2(G13), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n325), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT12), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n339), .B(new_n340), .C1(KEYINPUT76), .C2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT76), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n342), .B1(new_n343), .B2(KEYINPUT12), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n339), .A2(new_n340), .A3(KEYINPUT76), .A4(new_n341), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n300), .A2(new_n211), .A3(new_n296), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n202), .B1(new_n215), .B2(G20), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n344), .A2(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n333), .A2(new_n337), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n270), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n351), .B1(G238), .B2(new_n262), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G33), .A2(G97), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT73), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT73), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(G33), .A3(G97), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(G226), .B(new_n253), .C1(new_n250), .C2(new_n251), .ZN(new_n358));
  OAI211_X1 g0158(.A(G232), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n360), .A2(KEYINPUT74), .A3(new_n258), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT74), .B1(new_n360), .B2(new_n258), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n352), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT13), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT13), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n365), .B(new_n352), .C1(new_n361), .C2(new_n362), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(G179), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(KEYINPUT77), .A2(G169), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n364), .B2(new_n366), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT14), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n367), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI211_X1 g0171(.A(KEYINPUT14), .B(new_n368), .C1(new_n364), .C2(new_n366), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n350), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n364), .A2(G190), .A3(new_n366), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n349), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G200), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(new_n364), .B2(new_n366), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n324), .A2(new_n373), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n277), .A2(G222), .A3(new_n253), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n277), .A2(G223), .A3(G1698), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n380), .B(new_n381), .C1(new_n327), .C2(new_n277), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n258), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n351), .B1(G226), .B2(new_n262), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G169), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n206), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n212), .B1(new_n388), .B2(new_n328), .ZN(new_n389));
  INV_X1    g0189(.A(G150), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n299), .A2(new_n326), .B1(new_n390), .B2(new_n286), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n297), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n304), .A2(G50), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n306), .A2(new_n393), .B1(G50), .B2(new_n300), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n394), .B(KEYINPUT66), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n387), .B(new_n396), .C1(G179), .C2(new_n385), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT10), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT9), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT71), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n396), .A2(KEYINPUT71), .A3(new_n400), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n392), .A2(new_n395), .A3(KEYINPUT9), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n385), .A2(G200), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n383), .A2(new_n384), .A3(G190), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n399), .B1(new_n405), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n405), .A2(new_n410), .A3(new_n399), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n398), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI211_X1 g0214(.A(G232), .B(new_n253), .C1(new_n250), .C2(new_n251), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT67), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT67), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n277), .A2(new_n417), .A3(G232), .A4(new_n253), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n279), .A2(G107), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n277), .A2(G238), .A3(G1698), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n416), .A2(new_n418), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n258), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n351), .B1(G244), .B2(new_n262), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT68), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n422), .A2(KEYINPUT68), .A3(new_n423), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n426), .A2(G200), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n304), .A2(G77), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n306), .A2(new_n429), .B1(G77), .B2(new_n300), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n303), .A2(new_n287), .B1(G20), .B2(G77), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT15), .B(G87), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n431), .B1(new_n326), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n297), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT69), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT69), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n433), .A2(new_n436), .A3(new_n297), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n430), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT70), .B1(new_n428), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT70), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n426), .A2(new_n427), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n441), .B(new_n438), .C1(new_n442), .C2(new_n376), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(G190), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n440), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n442), .A2(new_n315), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n426), .A2(new_n386), .A3(new_n427), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(new_n439), .A3(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n414), .A2(KEYINPUT72), .A3(new_n445), .A4(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT72), .ZN(new_n450));
  AOI211_X1 g0250(.A(KEYINPUT10), .B(new_n409), .C1(new_n403), .C2(new_n404), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n448), .B(new_n397), .C1(new_n451), .C2(new_n411), .ZN(new_n452));
  INV_X1    g0252(.A(new_n445), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n379), .B1(new_n449), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n432), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(new_n300), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n215), .A2(G33), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n300), .A2(new_n459), .A3(new_n211), .A4(new_n296), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(new_n432), .ZN(new_n461));
  NOR2_X1   g0261(.A1(G97), .A2(G107), .ZN(new_n462));
  INV_X1    g0262(.A(G87), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT19), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n465), .B1(new_n354), .B2(new_n356), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n464), .B1(new_n466), .B2(G20), .ZN(new_n467));
  OR2_X1    g0267(.A1(KEYINPUT3), .A2(G33), .ZN(new_n468));
  NAND2_X1  g0268(.A1(KEYINPUT3), .A2(G33), .ZN(new_n469));
  AOI21_X1  g0269(.A(G20), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n212), .A2(G33), .A3(G97), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n470), .A2(G68), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  AOI211_X1 g0273(.A(new_n458), .B(new_n461), .C1(new_n473), .C2(new_n297), .ZN(new_n474));
  INV_X1    g0274(.A(G45), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(G1), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n257), .A2(G274), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n215), .A2(G45), .ZN(new_n478));
  AND2_X1   g0278(.A1(G33), .A2(G41), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n478), .B(G250), .C1(new_n479), .C2(new_n211), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(G244), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n482));
  OAI211_X1 g0282(.A(G238), .B(new_n253), .C1(new_n250), .C2(new_n251), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G116), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n481), .B1(new_n485), .B2(new_n258), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n315), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n486), .A2(G169), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n474), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n486), .A2(G190), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n485), .A2(new_n258), .ZN(new_n493));
  INV_X1    g0293(.A(new_n481), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G200), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n458), .B1(new_n473), .B2(new_n297), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n346), .A2(G87), .A3(new_n459), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n492), .B1(new_n499), .B2(KEYINPUT84), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT84), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n496), .A2(new_n497), .A3(new_n501), .A4(new_n498), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n490), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(G244), .B(new_n253), .C1(new_n250), .C2(new_n251), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G283), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G250), .A2(G1698), .ZN(new_n509));
  NAND2_X1  g0309(.A1(KEYINPUT4), .A2(G244), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(new_n510), .B2(G1698), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n508), .B1(new_n277), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n258), .ZN(new_n514));
  AND2_X1   g0314(.A1(KEYINPUT5), .A2(G41), .ZN(new_n515));
  NOR2_X1   g0315(.A1(KEYINPUT5), .A2(G41), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(G257), .B(new_n257), .C1(new_n517), .C2(new_n478), .ZN(new_n518));
  XNOR2_X1  g0318(.A(KEYINPUT5), .B(G41), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n519), .A2(G274), .A3(new_n257), .A4(new_n476), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n514), .A2(new_n268), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n257), .B1(new_n506), .B2(new_n512), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n518), .A2(new_n520), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n376), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n297), .ZN(new_n527));
  OAI21_X1  g0327(.A(G107), .B1(new_n291), .B2(new_n292), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT6), .ZN(new_n529));
  AND2_X1   g0329(.A1(G97), .A2(G107), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n529), .B1(new_n530), .B2(new_n462), .ZN(new_n531));
  INV_X1    g0331(.A(G107), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n532), .A2(KEYINPUT6), .A3(G97), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n534), .A2(G20), .B1(G77), .B2(new_n287), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n527), .B1(new_n528), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(G97), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n301), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n460), .B2(new_n537), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT81), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n526), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n541), .B1(new_n526), .B2(new_n540), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n539), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n528), .A2(new_n535), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(new_n527), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT82), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n386), .B1(new_n523), .B2(new_n524), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n514), .A2(new_n315), .A3(new_n521), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n547), .A2(new_n548), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n550), .B(new_n549), .C1(new_n536), .C2(new_n539), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT82), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT83), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n544), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  XNOR2_X1  g0356(.A(new_n552), .B(new_n548), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n526), .A2(new_n540), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT81), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n526), .A2(new_n540), .A3(new_n541), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT83), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n503), .B1(new_n556), .B2(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(G257), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n564));
  OAI211_X1 g0364(.A(G250), .B(new_n253), .C1(new_n250), .C2(new_n251), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G294), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n519), .A2(new_n476), .B1(new_n264), .B2(new_n256), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n567), .A2(new_n258), .B1(new_n568), .B2(G264), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(new_n315), .A3(new_n520), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n520), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n386), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n212), .B(G87), .C1(new_n250), .C2(new_n251), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT22), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT22), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n277), .A2(new_n575), .A3(new_n212), .A4(G87), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n484), .A2(G20), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT23), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n212), .B2(G107), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n532), .A2(KEYINPUT23), .A3(G20), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n578), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT24), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT24), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n577), .A2(new_n585), .A3(new_n582), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n527), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n301), .A2(new_n532), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n588), .B(KEYINPUT25), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n460), .A2(new_n532), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n570), .B(new_n572), .C1(new_n587), .C2(new_n592), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n577), .A2(new_n585), .A3(new_n582), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n585), .B1(new_n577), .B2(new_n582), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n297), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n569), .A2(new_n268), .A3(new_n520), .ZN(new_n597));
  AOI21_X1  g0397(.A(G200), .B1(new_n569), .B2(new_n520), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n596), .B(new_n591), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(G116), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(G20), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n338), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n507), .B(new_n212), .C1(G33), .C2(new_n537), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n604), .A2(new_n297), .A3(new_n602), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT20), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n604), .A2(KEYINPUT20), .A3(new_n297), .A4(new_n602), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n603), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n346), .A2(KEYINPUT86), .A3(G116), .A4(new_n459), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT86), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n460), .B2(new_n601), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(G270), .B(new_n257), .C1(new_n517), .C2(new_n478), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n520), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(G264), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n618));
  OAI211_X1 g0418(.A(G257), .B(new_n253), .C1(new_n250), .C2(new_n251), .ZN(new_n619));
  XNOR2_X1  g0419(.A(KEYINPUT85), .B(G303), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n618), .B(new_n619), .C1(new_n277), .C2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n258), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n614), .A2(new_n623), .A3(G169), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT87), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT21), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n616), .B1(new_n258), .B2(new_n621), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(G190), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n623), .A2(G200), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n629), .A2(new_n630), .A3(new_n613), .A4(new_n609), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n614), .A2(new_n628), .A3(G179), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n625), .A2(new_n626), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n614), .A2(new_n623), .A3(G169), .A4(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n627), .A2(new_n631), .A3(new_n632), .A4(new_n634), .ZN(new_n635));
  NOR4_X1   g0435(.A1(new_n456), .A2(new_n563), .A3(new_n600), .A4(new_n635), .ZN(G372));
  NAND4_X1  g0436(.A1(new_n496), .A2(new_n497), .A3(new_n498), .A4(new_n491), .ZN(new_n637));
  INV_X1    g0437(.A(new_n461), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n497), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT88), .B1(new_n486), .B2(G169), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT88), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n495), .A2(new_n641), .A3(new_n386), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n639), .A2(new_n487), .A3(new_n640), .A4(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n599), .A2(new_n637), .A3(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n634), .A2(new_n632), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n593), .A2(new_n645), .A3(new_n627), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n644), .A2(new_n646), .A3(new_n557), .A4(new_n561), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT89), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n544), .A2(new_n554), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT89), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n649), .A2(new_n650), .A3(new_n646), .A4(new_n644), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n552), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n643), .A2(new_n653), .A3(new_n654), .A4(new_n637), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n643), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n503), .A2(new_n554), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n656), .B1(new_n657), .B2(KEYINPUT26), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n652), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n455), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT90), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n318), .A2(new_n317), .ZN(new_n662));
  INV_X1    g0462(.A(new_n448), .ZN(new_n663));
  INV_X1    g0463(.A(new_n368), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n360), .A2(new_n258), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT74), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n360), .A2(KEYINPUT74), .A3(new_n258), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n365), .B1(new_n669), .B2(new_n352), .ZN(new_n670));
  INV_X1    g0470(.A(new_n366), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n664), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT14), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n369), .A2(new_n370), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n674), .A3(new_n367), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n663), .B1(new_n675), .B2(new_n350), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n310), .B(KEYINPUT17), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n378), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n662), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n412), .A2(new_n413), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n398), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n661), .A2(new_n681), .ZN(G369));
  NOR3_X1   g0482(.A1(new_n338), .A2(KEYINPUT27), .A3(G20), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT91), .Z(new_n684));
  INV_X1    g0484(.A(G213), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT27), .B1(new_n338), .B2(G20), .ZN(new_n687));
  XOR2_X1   g0487(.A(new_n687), .B(KEYINPUT92), .Z(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n691), .A2(new_n614), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n645), .A2(new_n627), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n635), .B2(new_n692), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G330), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n691), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n699), .B1(new_n596), .B2(new_n591), .ZN(new_n700));
  OAI22_X1  g0500(.A1(new_n700), .A2(new_n600), .B1(new_n593), .B2(new_n699), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n693), .A2(new_n699), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n600), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n593), .A2(new_n691), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n702), .A2(new_n706), .ZN(G399));
  INV_X1    g0507(.A(new_n218), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n464), .A2(G116), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G1), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n209), .B2(new_n710), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT26), .B1(new_n503), .B2(new_n554), .ZN(new_n715));
  AND4_X1   g0515(.A1(KEYINPUT26), .A2(new_n643), .A3(new_n653), .A4(new_n637), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n647), .B(new_n643), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n717), .A2(KEYINPUT94), .A3(new_n699), .ZN(new_n718));
  AOI21_X1  g0518(.A(KEYINPUT94), .B1(new_n717), .B2(new_n699), .ZN(new_n719));
  OAI21_X1  g0519(.A(KEYINPUT29), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n657), .A2(KEYINPUT26), .ZN(new_n722));
  INV_X1    g0522(.A(new_n656), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n724), .B1(new_n648), .B2(new_n651), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n721), .B1(new_n725), .B2(new_n691), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n720), .A2(new_n726), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n635), .A2(new_n600), .A3(new_n691), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n503), .B(new_n728), .C1(new_n556), .C2(new_n562), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n514), .A2(new_n569), .A3(new_n486), .A4(new_n521), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n617), .A2(new_n622), .A3(G179), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n486), .A2(G179), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n514), .A2(new_n521), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n734), .A2(new_n571), .A3(new_n735), .A4(new_n623), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n731), .A2(new_n730), .A3(new_n732), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT93), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n733), .B(new_n736), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n514), .A2(new_n486), .A3(new_n521), .ZN(new_n740));
  AND3_X1   g0540(.A1(new_n617), .A2(new_n622), .A3(G179), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n740), .A2(new_n741), .A3(KEYINPUT30), .A4(new_n569), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(KEYINPUT93), .ZN(new_n743));
  OAI211_X1 g0543(.A(KEYINPUT31), .B(new_n691), .C1(new_n739), .C2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n742), .A2(KEYINPUT93), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n731), .A2(new_n732), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(new_n738), .A3(KEYINPUT30), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n746), .A2(new_n748), .A3(new_n733), .A4(new_n736), .ZN(new_n749));
  AOI21_X1  g0549(.A(KEYINPUT31), .B1(new_n749), .B2(new_n691), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n697), .B1(new_n729), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n727), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n714), .B1(new_n755), .B2(G1), .ZN(G364));
  INV_X1    g0556(.A(G13), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n215), .B1(new_n758), .B2(G45), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n709), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n698), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(G330), .B2(new_n695), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n708), .A2(new_n279), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G355), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(G116), .B2(new_n218), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n708), .A2(new_n277), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n768), .B1(new_n210), .B2(new_n475), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n242), .A2(new_n475), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n766), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G13), .A2(G33), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT95), .Z(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n211), .B1(G20), .B2(new_n386), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n761), .B1(new_n771), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G311), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n212), .A2(new_n315), .A3(KEYINPUT96), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT96), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(G20), .B2(G179), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G190), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n268), .A2(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G322), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n779), .A2(new_n786), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n212), .A2(G179), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n785), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n277), .B1(new_n793), .B2(G329), .ZN(new_n794));
  INV_X1    g0594(.A(G283), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n791), .A2(new_n268), .A3(G200), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n787), .A2(new_n315), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G20), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G294), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n791), .A2(G190), .A3(G200), .ZN(new_n802));
  INV_X1    g0602(.A(G303), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n800), .A2(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n790), .A2(new_n797), .A3(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G326), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n783), .A2(new_n376), .ZN(new_n807));
  AND3_X1   g0607(.A1(new_n807), .A2(KEYINPUT97), .A3(G190), .ZN(new_n808));
  AOI21_X1  g0608(.A(KEYINPUT97), .B1(new_n807), .B2(G190), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AND3_X1   g0610(.A1(new_n807), .A2(KEYINPUT98), .A3(new_n268), .ZN(new_n811));
  AOI21_X1  g0611(.A(KEYINPUT98), .B1(new_n807), .B2(new_n268), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(KEYINPUT33), .B(G317), .Z(new_n814));
  OAI221_X1 g0614(.A(new_n805), .B1(new_n806), .B2(new_n810), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n815), .A2(KEYINPUT99), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n279), .B1(new_n799), .B2(G97), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n817), .B1(new_n786), .B2(new_n327), .C1(new_n201), .C2(new_n788), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n796), .A2(new_n532), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n802), .A2(new_n463), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n793), .A2(G159), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT32), .ZN(new_n822));
  NOR4_X1   g0622(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n823), .B1(new_n328), .B2(new_n810), .C1(new_n202), .C2(new_n813), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n815), .A2(KEYINPUT99), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n816), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n778), .B1(new_n826), .B2(new_n775), .ZN(new_n827));
  INV_X1    g0627(.A(new_n774), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n695), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n763), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(G396));
  NAND2_X1  g0631(.A1(new_n448), .A2(KEYINPUT100), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n439), .A2(new_n691), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT100), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n446), .A2(new_n834), .A3(new_n439), .A4(new_n447), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n445), .A2(new_n832), .A3(new_n833), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n663), .A2(new_n691), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n725), .B2(new_n691), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n832), .A2(new_n835), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n453), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n659), .A2(new_n699), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n752), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT101), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n761), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n844), .A2(new_n845), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n840), .A2(new_n752), .A3(new_n843), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n846), .A2(new_n847), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n775), .ZN(new_n851));
  INV_X1    g0651(.A(new_n788), .ZN(new_n852));
  INV_X1    g0652(.A(new_n786), .ZN(new_n853));
  AOI22_X1  g0653(.A1(G143), .A2(new_n852), .B1(new_n853), .B2(G159), .ZN(new_n854));
  INV_X1    g0654(.A(G137), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n854), .B1(new_n813), .B2(new_n390), .C1(new_n855), .C2(new_n810), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT34), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n796), .A2(new_n202), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n279), .B(new_n858), .C1(G132), .C2(new_n793), .ZN(new_n859));
  INV_X1    g0659(.A(new_n802), .ZN(new_n860));
  AOI22_X1  g0660(.A1(G50), .A2(new_n860), .B1(new_n799), .B2(G58), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n857), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n601), .A2(new_n786), .B1(new_n788), .B2(new_n801), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n279), .B1(new_n792), .B2(new_n779), .C1(new_n800), .C2(new_n537), .ZN(new_n864));
  INV_X1    g0664(.A(new_n796), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(G87), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n532), .B2(new_n802), .ZN(new_n867));
  NOR3_X1   g0667(.A1(new_n863), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n868), .B1(new_n795), .B2(new_n813), .C1(new_n803), .C2(new_n810), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n851), .B1(new_n862), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n775), .A2(new_n772), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n847), .B(new_n870), .C1(new_n327), .C2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n773), .B2(new_n838), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n850), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(G384));
  OR2_X1    g0675(.A1(new_n534), .A2(KEYINPUT35), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n534), .A2(KEYINPUT35), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n876), .A2(G116), .A3(new_n213), .A4(new_n877), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT36), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n210), .A2(G77), .A3(new_n282), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(G50), .B2(new_n202), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(G1), .A3(new_n757), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n882), .B(KEYINPUT102), .Z(new_n883));
  NOR2_X1   g0683(.A1(new_n375), .A2(new_n377), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n350), .B(new_n691), .C1(new_n675), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n350), .A2(new_n691), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n373), .A2(new_n378), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n841), .A2(new_n699), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n889), .B1(new_n843), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  INV_X1    g0692(.A(new_n689), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n313), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n313), .A2(KEYINPUT80), .A3(new_n316), .A4(KEYINPUT18), .ZN(new_n895));
  INV_X1    g0695(.A(new_n317), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n323), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n894), .B1(new_n897), .B2(new_n677), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n894), .A2(new_n321), .A3(new_n310), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT37), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT37), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n894), .A2(new_n321), .A3(new_n901), .A4(new_n310), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n892), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n900), .A2(new_n902), .ZN(new_n905));
  OAI211_X1 g0705(.A(KEYINPUT38), .B(new_n905), .C1(new_n324), .C2(new_n894), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n891), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n894), .B1(new_n662), .B2(new_n677), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT104), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n899), .A2(new_n910), .A3(KEYINPUT37), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n910), .B1(new_n899), .B2(KEYINPUT37), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT105), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n902), .B(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n909), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  XOR2_X1   g0716(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n917));
  OAI21_X1  g0717(.A(new_n906), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT39), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n904), .A2(new_n906), .A3(KEYINPUT39), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n675), .A2(new_n350), .A3(new_n699), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n662), .A2(new_n893), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n908), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n720), .A2(new_n455), .A3(new_n726), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n681), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n926), .B(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n729), .A2(new_n751), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(new_n838), .A3(new_n888), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT106), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n729), .A2(new_n751), .B1(new_n836), .B2(new_n837), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(KEYINPUT106), .A3(new_n888), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n933), .A2(KEYINPUT40), .A3(new_n935), .A4(new_n918), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n907), .A2(new_n934), .A3(new_n888), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT40), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n455), .A2(new_n930), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n942), .A2(G330), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n929), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n215), .B2(new_n758), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n929), .A2(new_n944), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n879), .B(new_n883), .C1(new_n946), .C2(new_n947), .ZN(G367));
  INV_X1    g0748(.A(G317), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n279), .B1(new_n792), .B2(new_n949), .C1(new_n537), .C2(new_n796), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n802), .A2(new_n601), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n853), .A2(G283), .B1(KEYINPUT46), .B2(new_n951), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n952), .B1(KEYINPUT46), .B2(new_n951), .C1(new_n620), .C2(new_n788), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n950), .B(new_n953), .C1(G107), .C2(new_n799), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n954), .B1(new_n801), .B2(new_n813), .C1(new_n779), .C2(new_n810), .ZN(new_n955));
  INV_X1    g0755(.A(new_n810), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(G143), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n328), .A2(new_n786), .B1(new_n788), .B2(new_n390), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n277), .B1(new_n792), .B2(new_n855), .C1(new_n201), .C2(new_n802), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n800), .A2(new_n202), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n796), .A2(new_n327), .ZN(new_n961));
  NOR4_X1   g0761(.A1(new_n958), .A2(new_n959), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(G159), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n957), .B(new_n962), .C1(new_n963), .C2(new_n813), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n955), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT47), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n775), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n497), .A2(new_n498), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n691), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n969), .A2(new_n643), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n969), .A2(new_n643), .A3(new_n637), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n970), .A2(new_n774), .A3(new_n971), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n776), .B1(new_n218), .B2(new_n432), .C1(new_n768), .C2(new_n238), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT110), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n973), .A2(new_n974), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n975), .A2(new_n976), .A3(new_n847), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n967), .A2(new_n972), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n649), .B1(new_n540), .B2(new_n699), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n653), .A2(new_n691), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n704), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT42), .Z(new_n983));
  INV_X1    g0783(.A(new_n981), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n557), .B1(new_n984), .B2(new_n593), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n699), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n970), .A2(new_n971), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n983), .A2(new_n986), .B1(KEYINPUT43), .B2(new_n987), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(KEYINPUT43), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n989), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n702), .A2(new_n984), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n990), .B(new_n991), .C1(KEYINPUT107), .C2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(KEYINPUT107), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n993), .B(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n981), .A2(new_n706), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT45), .Z(new_n997));
  NOR2_X1   g0797(.A1(new_n981), .A2(new_n706), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT44), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(new_n702), .Z(new_n1001));
  INV_X1    g0801(.A(new_n704), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n703), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1002), .B(KEYINPUT108), .C1(new_n701), .C2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(KEYINPUT108), .B2(new_n1002), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n698), .A2(KEYINPUT109), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n755), .B1(new_n1001), .B2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n709), .B(KEYINPUT41), .Z(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n760), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n978), .B1(new_n995), .B2(new_n1012), .ZN(G387));
  NAND2_X1  g0813(.A1(new_n755), .A2(new_n1007), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1008), .A2(new_n754), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1014), .A2(new_n709), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n711), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n764), .A2(new_n1017), .B1(new_n532), .B2(new_n708), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n235), .A2(new_n475), .ZN(new_n1019));
  AOI21_X1  g0819(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n303), .A2(new_n328), .ZN(new_n1021));
  XOR2_X1   g0821(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n1022));
  OAI211_X1 g0822(.A(new_n711), .B(new_n1020), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n767), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1018), .B1(new_n1019), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n847), .B1(new_n1026), .B2(new_n776), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n701), .B2(new_n828), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n328), .A2(new_n788), .B1(new_n786), .B2(new_n202), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n277), .B1(new_n792), .B2(new_n390), .C1(new_n537), .C2(new_n796), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n800), .A2(new_n432), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n802), .A2(new_n327), .ZN(new_n1032));
  NOR4_X1   g0832(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n963), .B2(new_n810), .C1(new_n299), .C2(new_n813), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n620), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G317), .A2(new_n852), .B1(new_n853), .B2(new_n1035), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n813), .B2(new_n779), .C1(new_n789), .C2(new_n810), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT48), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G294), .A2(new_n860), .B1(new_n799), .B2(G283), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n279), .B1(new_n792), .B2(new_n806), .C1(new_n601), .C2(new_n796), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1034), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1028), .B1(new_n1048), .B2(new_n775), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n760), .B2(new_n1007), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1016), .A2(new_n1050), .ZN(G393));
  INV_X1    g0851(.A(new_n1014), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1000), .B(new_n702), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n710), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1001), .A2(new_n1014), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1053), .A2(new_n760), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n776), .B1(new_n537), .B2(new_n218), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n768), .A2(new_n245), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n761), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n956), .A2(G150), .B1(G159), .B2(new_n852), .ZN(new_n1061));
  XOR2_X1   g0861(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n800), .A2(new_n327), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G68), .B2(new_n860), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n853), .A2(new_n303), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n279), .B1(new_n793), .B2(G143), .ZN(new_n1067));
  AND4_X1   g0867(.A1(new_n866), .A2(new_n1065), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1063), .B(new_n1068), .C1(new_n328), .C2(new_n813), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n810), .A2(new_n949), .B1(new_n779), .B2(new_n788), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT52), .Z(new_n1072));
  NOR2_X1   g0872(.A1(new_n786), .A2(new_n801), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n800), .A2(new_n601), .B1(new_n802), .B2(new_n795), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n279), .B1(new_n792), .B2(new_n789), .ZN(new_n1075));
  NOR4_X1   g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n819), .A4(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n620), .B2(new_n813), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1069), .A2(new_n1070), .B1(new_n1072), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1060), .B1(new_n1078), .B2(new_n775), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n828), .B2(new_n981), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1056), .A2(new_n1057), .A3(new_n1080), .ZN(G390));
  NAND2_X1  g0881(.A1(new_n752), .A2(new_n838), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n889), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n838), .B1(new_n718), .B2(new_n719), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n930), .A2(G330), .A3(new_n888), .A4(new_n838), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n890), .A4(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n843), .A2(new_n890), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT114), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n888), .B1(new_n752), .B2(new_n838), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1087), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1088), .B(new_n888), .C1(new_n752), .C2(new_n838), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1086), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n455), .A2(new_n752), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n927), .A2(new_n681), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(KEYINPUT115), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT115), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1093), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1085), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1087), .A2(new_n888), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1102), .A2(new_n922), .B1(new_n920), .B2(new_n921), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n918), .A2(new_n922), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1084), .A2(new_n890), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1104), .B1(new_n1105), .B2(new_n888), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1101), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n920), .A2(new_n921), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n923), .B2(new_n891), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n889), .B1(new_n1084), .B2(new_n890), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1109), .B(new_n1085), .C1(new_n1110), .C2(new_n1104), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n710), .B1(new_n1100), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT116), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1093), .A2(new_n1098), .A3(new_n1095), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1098), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1115), .B1(new_n1118), .B2(new_n1112), .ZN(new_n1119));
  AND4_X1   g0919(.A1(new_n1115), .A2(new_n1112), .A3(new_n1097), .A4(new_n1099), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1114), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(G125), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n277), .B1(new_n792), .B2(new_n1122), .C1(new_n800), .C2(new_n963), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n802), .A2(new_n390), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT53), .ZN(new_n1125));
  INV_X1    g0925(.A(G132), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT54), .B(G143), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1125), .B1(new_n1126), .B2(new_n788), .C1(new_n786), .C2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1123), .B(new_n1128), .C1(G50), .C2(new_n865), .ZN(new_n1129));
  INV_X1    g0929(.A(G128), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1129), .B1(new_n1130), .B2(new_n810), .C1(new_n855), .C2(new_n813), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n537), .A2(new_n786), .B1(new_n788), .B2(new_n601), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n279), .B1(new_n792), .B2(new_n801), .C1(new_n463), .C2(new_n802), .ZN(new_n1133));
  NOR4_X1   g0933(.A1(new_n1132), .A2(new_n858), .A3(new_n1064), .A4(new_n1133), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1134), .B1(new_n532), .B2(new_n813), .C1(new_n795), .C2(new_n810), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n851), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n871), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n761), .B1(new_n1137), .B2(new_n303), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n773), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1136), .B(new_n1138), .C1(new_n1108), .C2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n1113), .B2(new_n760), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1121), .A2(new_n1141), .ZN(G378));
  OR2_X1    g0942(.A1(new_n802), .A2(new_n1127), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1143), .A2(KEYINPUT118), .B1(new_n800), .B2(new_n390), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(KEYINPUT118), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n786), .B2(new_n855), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1144), .B(new_n1146), .C1(G128), .C2(new_n852), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1147), .B1(new_n1122), .B2(new_n810), .C1(new_n1126), .C2(new_n813), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(KEYINPUT59), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n865), .A2(G159), .ZN(new_n1150));
  AOI211_X1 g0950(.A(G33), .B(G41), .C1(new_n793), .C2(G124), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n1148), .A2(KEYINPUT59), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n532), .A2(new_n788), .B1(new_n786), .B2(new_n432), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n277), .A2(G41), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1155), .B1(new_n795), .B2(new_n792), .C1(new_n800), .C2(new_n202), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n796), .A2(new_n201), .ZN(new_n1157));
  NOR4_X1   g0957(.A1(new_n1154), .A2(new_n1156), .A3(new_n1032), .A4(new_n1157), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1158), .B1(new_n537), .B2(new_n813), .C1(new_n601), .C2(new_n810), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT117), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1152), .A2(new_n1153), .B1(new_n1160), .B2(KEYINPUT58), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n328), .B1(G33), .B2(G41), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1161), .B1(KEYINPUT58), .B2(new_n1160), .C1(new_n1155), .C2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n775), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n847), .B1(new_n328), .B2(new_n871), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n893), .A2(new_n396), .ZN(new_n1166));
  XOR2_X1   g0966(.A(new_n1166), .B(KEYINPUT119), .Z(new_n1167));
  XOR2_X1   g0967(.A(new_n414), .B(new_n1167), .Z(new_n1168));
  XOR2_X1   g0968(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1169));
  XOR2_X1   g0969(.A(new_n1168), .B(new_n1169), .Z(new_n1170));
  OAI211_X1 g0970(.A(new_n1164), .B(new_n1165), .C1(new_n1170), .C2(new_n773), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n697), .B1(new_n937), .B2(new_n938), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n936), .A2(new_n1172), .A3(KEYINPUT120), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1168), .B(new_n1169), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(KEYINPUT120), .B1(new_n936), .B2(new_n1172), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n936), .A2(new_n1172), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1178), .A2(KEYINPUT120), .A3(new_n1174), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n926), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1176), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1181), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n926), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1180), .A2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1171), .B1(new_n1186), .B2(new_n759), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(new_n1177), .A2(new_n1179), .A3(new_n926), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1183), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1095), .B1(new_n1118), .B2(new_n1112), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT57), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1095), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n1100), .B2(new_n1113), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1180), .A2(KEYINPUT57), .A3(new_n1185), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n709), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1188), .B1(new_n1193), .B2(new_n1197), .ZN(G375));
  AND2_X1   g0998(.A1(new_n1093), .A2(new_n760), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1199), .A2(KEYINPUT121), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(KEYINPUT121), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n855), .A2(new_n788), .B1(new_n786), .B2(new_n390), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n802), .A2(new_n963), .B1(new_n792), .B2(new_n1130), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT122), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n800), .A2(new_n328), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n277), .B1(new_n796), .B2(new_n201), .ZN(new_n1206));
  NOR4_X1   g1006(.A1(new_n1202), .A2(new_n1204), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n1126), .B2(new_n810), .C1(new_n813), .C2(new_n1127), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n532), .A2(new_n786), .B1(new_n788), .B2(new_n795), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n279), .B1(new_n792), .B2(new_n803), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n800), .A2(new_n432), .B1(new_n802), .B2(new_n537), .ZN(new_n1211));
  NOR4_X1   g1011(.A1(new_n1209), .A2(new_n961), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n601), .B2(new_n813), .C1(new_n801), .C2(new_n810), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n851), .B1(new_n1208), .B2(new_n1213), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n847), .B(new_n1214), .C1(new_n202), .C2(new_n871), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n772), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1215), .B1(new_n1216), .B2(new_n888), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1200), .A2(new_n1201), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1097), .A2(new_n1099), .A3(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1219), .B1(new_n1010), .B2(new_n1221), .ZN(G381));
  AND3_X1   g1022(.A1(new_n1056), .A2(new_n1057), .A3(new_n1080), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1016), .A2(new_n830), .A3(new_n1050), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1223), .A2(new_n874), .A3(new_n1225), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n1226), .A2(G387), .A3(G381), .ZN(new_n1227));
  INV_X1    g1027(.A(G375), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1121), .A2(new_n1141), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT123), .Z(G407));
  NAND3_X1  g1031(.A1(new_n1228), .A2(new_n690), .A3(new_n1229), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(G407), .A2(G213), .A3(new_n1232), .ZN(G409));
  NAND2_X1  g1033(.A1(G393), .A2(G396), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1223), .B1(new_n1225), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(G390), .A2(new_n1224), .A3(new_n1234), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(G387), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT126), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n690), .A2(G213), .A3(G2897), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n709), .B1(new_n1242), .B2(KEYINPUT60), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1116), .A2(new_n1117), .A3(new_n1242), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT60), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1244), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT125), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1221), .A2(KEYINPUT60), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1250), .A2(KEYINPUT125), .A3(new_n1244), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(G384), .B1(new_n1252), .B2(new_n1219), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n874), .B(new_n1218), .C1(new_n1249), .C2(new_n1251), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1241), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT125), .B1(new_n1250), .B2(new_n1244), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1248), .B(new_n1243), .C1(new_n1221), .C2(KEYINPUT60), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1219), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n874), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1252), .A2(G384), .A3(new_n1219), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1241), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1195), .A2(new_n1186), .A3(new_n1010), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1121), .B(new_n1141), .C1(new_n1263), .C2(new_n1187), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(G375), .B2(new_n1229), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n690), .A2(G213), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1255), .A2(new_n1262), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1240), .B1(new_n1267), .B2(KEYINPUT61), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1261), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT61), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(KEYINPUT126), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1268), .A2(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1276));
  AND4_X1   g1076(.A1(KEYINPUT62), .A2(new_n1276), .A3(new_n1265), .A4(new_n1266), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT124), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1265), .A2(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(G378), .B(new_n1188), .C1(new_n1193), .C2(new_n1197), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(KEYINPUT124), .A3(new_n1264), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1280), .A2(new_n1276), .A3(new_n1282), .A4(new_n1266), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1277), .B1(new_n1278), .B2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1239), .B1(new_n1275), .B2(new_n1284), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1276), .A2(KEYINPUT63), .A3(new_n1265), .A4(new_n1266), .ZN(new_n1286));
  INV_X1    g1086(.A(G387), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1238), .B(new_n1287), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1286), .A2(new_n1273), .A3(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1283), .A2(new_n1290), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1280), .A2(new_n1282), .A3(new_n1266), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1289), .B(new_n1291), .C1(new_n1292), .C2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1285), .A2(new_n1294), .ZN(G405));
  AND2_X1   g1095(.A1(new_n1288), .A2(new_n1276), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1288), .A2(new_n1276), .ZN(new_n1297));
  OAI21_X1  g1097(.A(KEYINPUT127), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1239), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT127), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1288), .A2(new_n1276), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1298), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(G375), .A2(new_n1229), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1304), .A2(new_n1281), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1303), .A2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1298), .A2(new_n1305), .A3(new_n1302), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(G402));
endmodule


