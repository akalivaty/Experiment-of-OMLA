//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n562, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n602,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1127, new_n1128;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G113), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(G2105), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n466), .A2(G2105), .B1(G101), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g043(.A(KEYINPUT3), .B1(KEYINPUT64), .B2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(KEYINPUT64), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n472), .A2(KEYINPUT65), .A3(G137), .A4(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n475));
  AND3_X1   g050(.A1(KEYINPUT64), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n473), .B1(new_n476), .B2(new_n469), .ZN(new_n477));
  INV_X1    g052(.A(G137), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n468), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  AOI21_X1  g057(.A(new_n473), .B1(new_n470), .B2(new_n471), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n473), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n477), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(G136), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT66), .ZN(G162));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n461), .B2(new_n462), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT67), .B(KEYINPUT4), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT68), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n473), .C1(new_n476), .C2(new_n469), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT67), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT3), .B(G2104), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n502), .A2(new_n503), .A3(new_n504), .A4(new_n492), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n495), .A2(new_n497), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n507));
  INV_X1    g082(.A(G114), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(G2105), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n509), .B1(new_n483), .B2(G126), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n521), .B1(new_n519), .B2(KEYINPUT69), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n523), .A2(KEYINPUT6), .A3(G651), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n522), .A2(new_n524), .B1(new_n515), .B2(new_n516), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n514), .B1(new_n522), .B2(new_n524), .ZN(new_n526));
  AOI22_X1  g101(.A1(G88), .A2(new_n525), .B1(new_n526), .B2(G50), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n520), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(G166));
  NAND2_X1  g104(.A1(new_n525), .A2(G89), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n532), .A2(new_n533), .B1(new_n517), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n526), .A2(G51), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n530), .A2(new_n535), .A3(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  AOI22_X1  g113(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n519), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n526), .A2(G52), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n525), .A2(G90), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(G171));
  AOI22_X1  g118(.A1(G81), .A2(new_n525), .B1(new_n526), .B2(G43), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT70), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n519), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT71), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(new_n526), .A2(G53), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n525), .A2(G91), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n517), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n559));
  OAI211_X1 g134(.A(new_n557), .B(new_n558), .C1(new_n519), .C2(new_n559), .ZN(G299));
  INV_X1    g135(.A(G171), .ZN(G301));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n528), .B(new_n562), .ZN(G303));
  NAND2_X1  g138(.A1(new_n525), .A2(G87), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n526), .A2(G49), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(G288));
  AOI21_X1  g142(.A(KEYINPUT73), .B1(new_n525), .B2(G86), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n525), .A2(KEYINPUT73), .A3(G86), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n516), .ZN(new_n572));
  NOR2_X1   g147(.A1(KEYINPUT5), .A2(G543), .ZN(new_n573));
  OAI21_X1  g148(.A(G61), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(G73), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n514), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(G48), .B2(new_n526), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n571), .A2(new_n577), .ZN(G305));
  AOI22_X1  g153(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n519), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT74), .ZN(new_n581));
  AOI22_X1  g156(.A1(G85), .A2(new_n525), .B1(new_n526), .B2(G47), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n580), .A2(KEYINPUT74), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G290));
  INV_X1    g161(.A(G868), .ZN(new_n587));
  OR3_X1    g162(.A1(G171), .A2(KEYINPUT75), .A3(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT75), .B1(G171), .B2(new_n587), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n525), .A2(G92), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT10), .Z(new_n591));
  NAND2_X1  g166(.A1(new_n517), .A2(G66), .ZN(new_n592));
  INV_X1    g167(.A(G79), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(new_n514), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(G54), .B2(new_n526), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  OAI211_X1 g172(.A(new_n588), .B(new_n589), .C1(G868), .C2(new_n597), .ZN(G284));
  OAI211_X1 g173(.A(new_n588), .B(new_n589), .C1(G868), .C2(new_n597), .ZN(G321));
  NAND2_X1  g174(.A1(G299), .A2(new_n587), .ZN(new_n600));
  OR3_X1    g175(.A1(G168), .A2(KEYINPUT76), .A3(new_n587), .ZN(new_n601));
  OAI21_X1  g176(.A(KEYINPUT76), .B1(G168), .B2(new_n587), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(G297));
  NAND3_X1  g178(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n597), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND2_X1  g181(.A1(new_n597), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n503), .A2(new_n467), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT77), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(KEYINPUT13), .B(G2100), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n488), .A2(G135), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n483), .A2(G123), .ZN(new_n617));
  OR2_X1    g192(.A1(G99), .A2(G2105), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n618), .B(G2104), .C1(G111), .C2(new_n473), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n620), .A2(G2096), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(G2096), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n615), .A2(new_n621), .A3(new_n622), .ZN(G156));
  XOR2_X1   g198(.A(G2451), .B(G2454), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT16), .ZN(new_n625));
  XNOR2_X1  g200(.A(G1341), .B(G1348), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT14), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n631), .B2(new_n630), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n627), .B(new_n633), .Z(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(G14), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n638), .B1(new_n637), .B2(new_n635), .ZN(G401));
  XNOR2_X1  g214(.A(KEYINPUT79), .B(KEYINPUT18), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2084), .B(G2090), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT78), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT17), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n642), .A2(new_n643), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n640), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2096), .B(G2100), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n644), .ZN(new_n650));
  NOR2_X1   g225(.A1(G2072), .A2(G2078), .ZN(new_n651));
  OAI22_X1  g226(.A1(new_n650), .A2(new_n640), .B1(new_n444), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT80), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n649), .B(new_n653), .ZN(G227));
  XOR2_X1   g229(.A(G1971), .B(G1976), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT19), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1956), .B(G2474), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1961), .B(G1966), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n656), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n656), .A2(new_n659), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT20), .Z(new_n663));
  AOI211_X1 g238(.A(new_n661), .B(new_n663), .C1(new_n656), .C2(new_n660), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1991), .B(G1996), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT81), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1981), .B(G1986), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G229));
  NOR2_X1   g246(.A1(G16), .A2(G24), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n585), .B2(G16), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT84), .B(G1986), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT85), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n673), .B(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(G29), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G25), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n488), .A2(G131), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n483), .A2(G119), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n473), .A2(G107), .ZN(new_n681));
  OAI21_X1  g256(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n679), .B(new_n680), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT82), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n678), .B1(new_n685), .B2(new_n677), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT35), .B(G1991), .Z(new_n687));
  XOR2_X1   g262(.A(new_n686), .B(new_n687), .Z(new_n688));
  MUX2_X1   g263(.A(G6), .B(G305), .S(G16), .Z(new_n689));
  XOR2_X1   g264(.A(KEYINPUT32), .B(G1981), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G22), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G166), .B2(new_n692), .ZN(new_n694));
  INV_X1    g269(.A(G1971), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n692), .A2(G23), .ZN(new_n697));
  INV_X1    g272(.A(G288), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(new_n692), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT33), .B(G1976), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n691), .A2(new_n696), .A3(new_n701), .ZN(new_n702));
  OAI22_X1  g277(.A1(new_n688), .A2(KEYINPUT83), .B1(KEYINPUT34), .B2(new_n702), .ZN(new_n703));
  AOI211_X1 g278(.A(new_n676), .B(new_n703), .C1(KEYINPUT83), .C2(new_n688), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(KEYINPUT34), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT86), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT87), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(KEYINPUT36), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n707), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n692), .A2(G4), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n597), .B2(new_n692), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1348), .ZN(new_n713));
  NOR2_X1   g288(.A1(G5), .A2(G16), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT94), .Z(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G301), .B2(new_n692), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G1961), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n692), .A2(G21), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G168), .B2(new_n692), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(G1966), .Z(new_n720));
  INV_X1    g295(.A(KEYINPUT24), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n677), .B1(new_n721), .B2(G34), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n722), .A2(KEYINPUT89), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(G34), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n722), .B2(KEYINPUT89), .ZN(new_n725));
  OAI22_X1  g300(.A1(new_n481), .A2(new_n677), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G2084), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n677), .A2(G33), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT25), .Z(new_n731));
  INV_X1    g306(.A(G139), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(new_n477), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n503), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(new_n473), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n729), .B1(new_n736), .B2(new_n677), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(new_n442), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n717), .A2(new_n720), .A3(new_n728), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT27), .B(G1996), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n677), .A2(G32), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT90), .B(KEYINPUT26), .ZN(new_n742));
  AND3_X1   g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n744), .A2(new_n745), .B1(G105), .B2(new_n467), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n488), .A2(G141), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n483), .A2(G129), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT91), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n741), .B1(new_n750), .B2(new_n677), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT92), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n713), .B(new_n739), .C1(new_n740), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n692), .A2(G20), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT95), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT23), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G299), .B2(G16), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT96), .ZN(new_n758));
  INV_X1    g333(.A(G1956), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n753), .B(new_n760), .C1(new_n740), .C2(new_n752), .ZN(new_n761));
  NOR2_X1   g336(.A1(G29), .A2(G35), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G162), .B2(G29), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT29), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(G2090), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n677), .A2(G26), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT28), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n488), .A2(G140), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n483), .A2(G128), .ZN(new_n769));
  OR2_X1    g344(.A1(G104), .A2(G2105), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n770), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n767), .B1(new_n772), .B2(G29), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT88), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2067), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n692), .A2(G19), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n549), .B2(new_n692), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(G1341), .Z(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT30), .B(G28), .ZN(new_n779));
  OR2_X1    g354(.A1(KEYINPUT31), .A2(G11), .ZN(new_n780));
  NAND2_X1  g355(.A1(KEYINPUT31), .A2(G11), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n779), .A2(new_n677), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n620), .B2(new_n677), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT93), .Z(new_n784));
  NOR2_X1   g359(.A1(G164), .A2(new_n677), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G27), .B2(new_n677), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(new_n443), .ZN(new_n787));
  AOI211_X1 g362(.A(new_n784), .B(new_n787), .C1(new_n727), .C2(new_n726), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n765), .A2(new_n775), .A3(new_n778), .A4(new_n788), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n710), .A2(new_n761), .A3(new_n789), .ZN(G311));
  INV_X1    g365(.A(G311), .ZN(G150));
  NAND2_X1  g366(.A1(new_n597), .A2(G559), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT38), .ZN(new_n793));
  AOI22_X1  g368(.A1(G93), .A2(new_n525), .B1(new_n526), .B2(G55), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT97), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n519), .B2(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(new_n548), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n793), .B(new_n798), .Z(new_n799));
  AND2_X1   g374(.A1(new_n799), .A2(KEYINPUT39), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(KEYINPUT39), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n800), .A2(new_n801), .A3(G860), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n797), .A2(G860), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT98), .B(KEYINPUT37), .Z(new_n804));
  XOR2_X1   g379(.A(new_n803), .B(new_n804), .Z(new_n805));
  OR2_X1    g380(.A1(new_n802), .A2(new_n805), .ZN(G145));
  XNOR2_X1  g381(.A(G162), .B(new_n620), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(new_n481), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n810));
  INV_X1    g385(.A(G118), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(G2105), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n483), .A2(G130), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT101), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  AOI211_X1 g390(.A(new_n812), .B(new_n815), .C1(G142), .C2(new_n488), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(new_n684), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(new_n613), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT100), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n736), .B1(new_n749), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n819), .B2(new_n749), .ZN(new_n821));
  INV_X1    g396(.A(new_n736), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n750), .B2(new_n822), .ZN(new_n823));
  AND3_X1   g398(.A1(new_n506), .A2(KEYINPUT99), .A3(new_n510), .ZN(new_n824));
  AOI21_X1  g399(.A(KEYINPUT99), .B1(new_n506), .B2(new_n510), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n772), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n823), .B(new_n827), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n818), .A2(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n818), .A2(new_n828), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT102), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AND3_X1   g407(.A1(new_n818), .A2(new_n831), .A3(new_n828), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n809), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT103), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n829), .A2(new_n809), .ZN(new_n837));
  AOI21_X1  g412(.A(G37), .B1(new_n837), .B2(new_n830), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g415(.A1(new_n797), .A2(new_n587), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n585), .B(G288), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n843), .A2(KEYINPUT105), .ZN(new_n844));
  XNOR2_X1  g419(.A(G305), .B(new_n528), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(new_n843), .B2(KEYINPUT105), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n844), .B(new_n846), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT42), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n798), .B(new_n607), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n596), .B(G299), .Z(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n850), .B(KEYINPUT41), .Z(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  OAI211_X1 g428(.A(KEYINPUT104), .B(new_n851), .C1(new_n853), .C2(new_n849), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(KEYINPUT104), .B2(new_n851), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n848), .B(new_n855), .Z(new_n856));
  OAI21_X1  g431(.A(new_n841), .B1(new_n856), .B2(new_n587), .ZN(G295));
  OAI21_X1  g432(.A(new_n841), .B1(new_n856), .B2(new_n587), .ZN(G331));
  INV_X1    g433(.A(G37), .ZN(new_n859));
  AOI21_X1  g434(.A(G286), .B1(G171), .B2(KEYINPUT106), .ZN(new_n860));
  NOR2_X1   g435(.A1(G171), .A2(KEYINPUT106), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n860), .B(new_n861), .Z(new_n862));
  OR2_X1    g437(.A1(new_n862), .A2(new_n798), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT107), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n798), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(new_n864), .B2(new_n865), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(new_n850), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n863), .A2(new_n865), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n853), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n847), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n859), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n868), .A2(KEYINPUT108), .A3(new_n870), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT108), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n847), .B1(new_n871), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n873), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n877), .A2(KEYINPUT43), .ZN(new_n878));
  INV_X1    g453(.A(new_n873), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n869), .A2(new_n850), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(KEYINPUT109), .Z(new_n881));
  NOR2_X1   g456(.A1(new_n867), .A2(new_n853), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n872), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n879), .A2(new_n883), .A3(KEYINPUT43), .ZN(new_n884));
  OAI21_X1  g459(.A(KEYINPUT44), .B1(new_n878), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n879), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(new_n877), .B2(new_n886), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n885), .A2(new_n890), .ZN(G397));
  NAND2_X1  g466(.A1(G303), .A2(G8), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT55), .ZN(new_n893));
  INV_X1    g468(.A(G1384), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n511), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT50), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n468), .A2(new_n480), .A3(G40), .ZN(new_n897));
  AOI21_X1  g472(.A(G1384), .B1(new_n506), .B2(new_n510), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT50), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n901), .A2(G2090), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT99), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n511), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n506), .A2(KEYINPUT99), .A3(new_n510), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT45), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n906), .A2(G1384), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT110), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT110), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n904), .A2(new_n910), .A3(new_n905), .A4(new_n907), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n897), .B1(new_n898), .B2(KEYINPUT45), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n902), .B1(new_n915), .B2(new_n695), .ZN(new_n916));
  INV_X1    g491(.A(G8), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n893), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n913), .B1(new_n909), .B2(new_n911), .ZN(new_n919));
  OAI22_X1  g494(.A1(new_n919), .A2(G1971), .B1(G2090), .B2(new_n901), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT55), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n892), .B(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n922), .A3(G8), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT111), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n897), .A2(new_n898), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n924), .B1(new_n925), .B2(G8), .ZN(new_n926));
  AOI211_X1 g501(.A(KEYINPUT111), .B(new_n917), .C1(new_n897), .C2(new_n898), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(G1976), .ZN(new_n929));
  NOR2_X1   g504(.A1(G288), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT52), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(KEYINPUT113), .A2(KEYINPUT49), .ZN(new_n932));
  INV_X1    g507(.A(G1981), .ZN(new_n933));
  INV_X1    g508(.A(new_n570), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n577), .B(new_n933), .C1(new_n934), .C2(new_n568), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT112), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n571), .A2(KEYINPUT112), .A3(new_n933), .A4(new_n577), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n525), .A2(G86), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n933), .B1(new_n577), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n932), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n932), .ZN(new_n944));
  AOI211_X1 g519(.A(new_n941), .B(new_n944), .C1(new_n937), .C2(new_n938), .ZN(new_n945));
  OAI22_X1  g520(.A1(new_n943), .A2(new_n945), .B1(new_n927), .B2(new_n926), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT52), .B1(G288), .B2(new_n929), .ZN(new_n947));
  OAI221_X1 g522(.A(new_n947), .B1(new_n929), .B2(G288), .C1(new_n926), .C2(new_n927), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n931), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n918), .A2(new_n923), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT53), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(G2078), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n897), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n904), .A2(new_n894), .A3(new_n905), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n953), .B1(new_n954), .B2(new_n906), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n912), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G1961), .ZN(new_n957));
  INV_X1    g532(.A(new_n900), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT122), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT122), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n901), .A2(new_n962), .A3(new_n957), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n956), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT53), .B1(new_n919), .B2(new_n443), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n964), .A2(new_n965), .A3(G171), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT123), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT54), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT114), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n511), .A2(new_n969), .A3(new_n907), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(new_n511), .B2(new_n907), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n913), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n952), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n960), .ZN(new_n974));
  OAI21_X1  g549(.A(G171), .B1(new_n965), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n910), .B1(new_n826), .B2(new_n907), .ZN(new_n976));
  INV_X1    g551(.A(new_n911), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n443), .B(new_n914), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n951), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n912), .A2(new_n955), .B1(new_n960), .B2(KEYINPUT122), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n963), .A3(new_n980), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n975), .B(KEYINPUT123), .C1(new_n981), .C2(G171), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n950), .B1(new_n968), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT120), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n970), .A2(new_n971), .ZN(new_n985));
  AOI21_X1  g560(.A(G1966), .B1(new_n985), .B2(new_n914), .ZN(new_n986));
  XNOR2_X1  g561(.A(KEYINPUT115), .B(G2084), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n901), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n984), .B(G8), .C1(new_n986), .C2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(G168), .A2(new_n917), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(KEYINPUT51), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  OAI22_X1  g567(.A1(new_n972), .A2(G1966), .B1(new_n901), .B2(new_n987), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n984), .B1(new_n993), .B2(G8), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT121), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(G8), .B1(new_n986), .B2(new_n988), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT120), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT121), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n997), .A2(new_n998), .A3(new_n989), .A4(new_n991), .ZN(new_n999));
  INV_X1    g574(.A(new_n996), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT51), .B1(new_n1000), .B2(new_n990), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n995), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n993), .A2(new_n990), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n972), .A2(new_n952), .B1(new_n957), .B2(new_n901), .ZN(new_n1005));
  AOI211_X1 g580(.A(G2078), .B(new_n913), .C1(new_n909), .C2(new_n911), .ZN(new_n1006));
  OAI211_X1 g581(.A(G301), .B(new_n1005), .C1(new_n1006), .C2(KEYINPUT53), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT124), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n979), .A2(KEYINPUT124), .A3(G301), .A4(new_n1005), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(new_n981), .B2(G171), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1011), .A2(KEYINPUT125), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT125), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n983), .B(new_n1004), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT59), .ZN(new_n1018));
  AOI211_X1 g593(.A(G1996), .B(new_n913), .C1(new_n909), .C2(new_n911), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n897), .A2(KEYINPUT116), .A3(new_n898), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT116), .B1(new_n897), .B2(new_n898), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT58), .B(G1341), .Z(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1018), .B(new_n549), .C1(new_n1019), .C2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT118), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n1027));
  INV_X1    g602(.A(G1996), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1028), .B(new_n914), .C1(new_n976), .C2(new_n977), .ZN(new_n1029));
  OR3_X1    g604(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n548), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1027), .B1(new_n1031), .B2(new_n1018), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n1033), .A3(new_n1018), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1024), .B1(new_n919), .B2(new_n1028), .ZN(new_n1035));
  OAI211_X1 g610(.A(KEYINPUT117), .B(KEYINPUT59), .C1(new_n1035), .C2(new_n548), .ZN(new_n1036));
  AND4_X1   g611(.A1(new_n1026), .A2(new_n1032), .A3(new_n1034), .A4(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT61), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT56), .B(G2072), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  AOI211_X1 g615(.A(new_n913), .B(new_n1040), .C1(new_n909), .C2(new_n911), .ZN(new_n1041));
  XNOR2_X1  g616(.A(G299), .B(KEYINPUT57), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n901), .A2(new_n759), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1042), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n912), .A2(new_n914), .A3(new_n1039), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1046), .B1(new_n1047), .B2(new_n1043), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1038), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1042), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1047), .A2(new_n1046), .A3(new_n1043), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n1051), .A3(KEYINPUT61), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1017), .B1(new_n1037), .B2(new_n1053), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1026), .A2(new_n1032), .A3(new_n1034), .A4(new_n1036), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(KEYINPUT119), .A3(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n958), .A2(new_n959), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n1058), .A2(G1348), .ZN(new_n1059));
  INV_X1    g634(.A(G2067), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1063), .A2(KEYINPUT60), .A3(new_n596), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT60), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n597), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1064), .A2(new_n1066), .B1(new_n1065), .B2(new_n1062), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1054), .A2(new_n1057), .A3(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1063), .A2(new_n596), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1051), .B1(new_n1070), .B2(new_n1048), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1016), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1000), .A2(G168), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n950), .A2(new_n1073), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n1074), .A2(KEYINPUT63), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(KEYINPUT63), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n946), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n698), .A2(new_n929), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n939), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n927), .B2(new_n926), .ZN(new_n1081));
  INV_X1    g656(.A(new_n923), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n949), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1077), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT126), .B1(new_n1072), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT126), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1084), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1071), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1067), .B1(new_n1091), .B2(new_n1017), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1090), .B1(new_n1092), .B2(new_n1057), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1088), .B(new_n1089), .C1(new_n1093), .C2(new_n1016), .ZN(new_n1094));
  AOI211_X1 g669(.A(new_n950), .B(new_n975), .C1(new_n1004), .C2(KEYINPUT62), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(KEYINPUT62), .B2(new_n1004), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1087), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n750), .A2(new_n1028), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n772), .B(new_n1060), .ZN(new_n1099));
  INV_X1    g674(.A(new_n749), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1098), .B(new_n1099), .C1(new_n1028), .C2(new_n1100), .ZN(new_n1101));
  XOR2_X1   g676(.A(new_n684), .B(new_n687), .Z(new_n1102));
  NOR2_X1   g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n585), .B(G1986), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT45), .B1(new_n826), .B2(new_n894), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n897), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1097), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n897), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(new_n1100), .B2(new_n1099), .ZN(new_n1110));
  OR3_X1    g685(.A1(new_n1109), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT46), .B1(new_n1109), .B2(G1996), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  XOR2_X1   g688(.A(new_n1113), .B(KEYINPUT47), .Z(new_n1114));
  NAND2_X1  g689(.A1(new_n685), .A2(new_n687), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1101), .A2(new_n1115), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n772), .A2(G2067), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1103), .A2(new_n1109), .ZN(new_n1119));
  XOR2_X1   g694(.A(new_n1119), .B(KEYINPUT127), .Z(new_n1120));
  NOR3_X1   g695(.A1(new_n1109), .A2(G1986), .A3(G290), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT48), .ZN(new_n1122));
  OAI221_X1 g697(.A(new_n1114), .B1(new_n1109), .B2(new_n1118), .C1(new_n1120), .C2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1108), .A2(new_n1124), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g700(.A(G319), .ZN(new_n1127));
  NOR4_X1   g701(.A1(G229), .A2(new_n1127), .A3(G401), .A4(G227), .ZN(new_n1128));
  NAND3_X1  g702(.A1(new_n888), .A2(new_n839), .A3(new_n1128), .ZN(G225));
  INV_X1    g703(.A(G225), .ZN(G308));
endmodule


