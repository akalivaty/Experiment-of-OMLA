//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1207,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT65), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n215), .A2(new_n216), .B1(G77), .B2(G244), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G50), .A2(G226), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G68), .A2(G238), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  AND2_X1   g0021(.A1(G116), .A2(G270), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT66), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n223), .B1(new_n224), .B2(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(G50), .B1(G58), .B2(G68), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT64), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n209), .B(new_n227), .C1(new_n230), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  AND2_X1   g0049(.A1(G1), .A2(G13), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G238), .ZN(new_n257));
  INV_X1    g0057(.A(G274), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT67), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT67), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G41), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  AOI211_X1 g0064(.A(G1), .B(new_n258), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n235), .A2(G1698), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G226), .B2(G1698), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G97), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT72), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n252), .A2(KEYINPUT68), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT68), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n279), .B1(new_n250), .B2(new_n251), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n257), .B(new_n266), .C1(new_n277), .C2(new_n281), .ZN(new_n282));
  OR2_X1    g0082(.A1(new_n282), .A2(KEYINPUT13), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(KEYINPUT13), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(KEYINPUT73), .A3(new_n284), .ZN(new_n285));
  OR3_X1    g0085(.A1(new_n282), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(G169), .A3(new_n286), .ZN(new_n287));
  OR2_X1    g0087(.A1(new_n287), .A2(KEYINPUT14), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n283), .A2(KEYINPUT74), .A3(new_n284), .ZN(new_n289));
  OR3_X1    g0089(.A1(new_n282), .A2(KEYINPUT74), .A3(KEYINPUT13), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G179), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n287), .A2(KEYINPUT14), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n288), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G20), .A2(G33), .ZN(new_n295));
  INV_X1    g0095(.A(G68), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n295), .A2(G50), .B1(G20), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G77), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n229), .A2(G33), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n228), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT11), .ZN(new_n304));
  INV_X1    g0104(.A(G13), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(G1), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(G20), .A3(new_n296), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT12), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n302), .B1(new_n253), .B2(G20), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n304), .B(new_n308), .C1(new_n296), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n294), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n311), .B1(new_n291), .B2(G190), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n285), .A2(G200), .A3(new_n286), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n252), .B(KEYINPUT68), .ZN(new_n316));
  INV_X1    g0116(.A(new_n273), .ZN(new_n317));
  NOR2_X1   g0117(.A1(G232), .A2(G1698), .ZN(new_n318));
  INV_X1    g0118(.A(G1698), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(G238), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n317), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n316), .B(new_n321), .C1(G107), .C2(new_n317), .ZN(new_n322));
  INV_X1    g0122(.A(G244), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n322), .B(new_n266), .C1(new_n323), .C2(new_n255), .ZN(new_n324));
  INV_X1    g0124(.A(G169), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n309), .A2(G77), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT70), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT8), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(G58), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(G58), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n295), .ZN(new_n334));
  OAI22_X1  g0134(.A1(new_n333), .A2(new_n334), .B1(new_n229), .B2(new_n298), .ZN(new_n335));
  XOR2_X1   g0135(.A(KEYINPUT15), .B(G87), .Z(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(new_n299), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n302), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n305), .A2(new_n229), .A3(G1), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n328), .B(new_n339), .C1(G77), .C2(new_n341), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n326), .B(new_n342), .C1(G179), .C2(new_n324), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n324), .A2(G200), .ZN(new_n344));
  INV_X1    g0144(.A(G190), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n344), .B1(new_n345), .B2(new_n324), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n346), .A2(new_n342), .ZN(new_n347));
  AND4_X1   g0147(.A1(new_n312), .A2(new_n315), .A3(new_n343), .A4(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT9), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT69), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n332), .B1(new_n330), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n350), .B2(new_n332), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n352), .A2(new_n229), .A3(G33), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n203), .A2(G20), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n295), .A2(G150), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n356), .A2(new_n302), .B1(new_n202), .B2(new_n340), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n309), .A2(G50), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n349), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n357), .A2(new_n349), .A3(new_n358), .ZN(new_n361));
  NOR2_X1   g0161(.A1(G222), .A2(G1698), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n319), .A2(G223), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n317), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n316), .B(new_n364), .C1(G77), .C2(new_n317), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n256), .A2(G226), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(new_n266), .A3(new_n366), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n360), .A2(new_n361), .B1(G200), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT71), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT10), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n367), .A2(new_n345), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n368), .A2(new_n369), .A3(new_n370), .A4(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n367), .A2(G200), .ZN(new_n374));
  INV_X1    g0174(.A(new_n361), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n369), .B(new_n374), .C1(new_n375), .C2(new_n359), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT10), .B1(new_n376), .B2(new_n371), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n357), .A2(new_n358), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n367), .A2(G179), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n367), .A2(new_n325), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n271), .A2(KEYINPUT75), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT75), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G33), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n269), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT7), .B1(new_n390), .B2(G20), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n392), .B(new_n229), .C1(new_n388), .C2(new_n389), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(G68), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g0194(.A(G58), .B(G68), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n395), .A2(G20), .B1(G159), .B2(new_n295), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n394), .A2(KEYINPUT16), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT76), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT7), .B1(new_n273), .B2(new_n229), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n385), .A2(new_n387), .A3(new_n269), .ZN(new_n400));
  AOI21_X1  g0200(.A(G20), .B1(new_n400), .B2(new_n272), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n399), .B1(new_n401), .B2(KEYINPUT7), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n396), .B1(new_n402), .B2(new_n296), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT16), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT76), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n394), .A2(new_n406), .A3(KEYINPUT16), .A4(new_n396), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n398), .A2(new_n302), .A3(new_n405), .A4(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n310), .A2(new_n352), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n340), .B2(new_n352), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n385), .A2(new_n387), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT3), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n270), .ZN(new_n414));
  NOR2_X1   g0214(.A1(G223), .A2(G1698), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n319), .A2(G226), .ZN(new_n416));
  NOR3_X1   g0216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n271), .A2(new_n211), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n316), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n256), .A2(G232), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n266), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G169), .ZN(new_n422));
  INV_X1    g0222(.A(G179), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n423), .B2(new_n421), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n411), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n411), .A2(new_n424), .A3(KEYINPUT18), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n421), .A2(new_n345), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n421), .A2(G200), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n408), .A2(new_n430), .A3(new_n410), .A4(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT17), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n432), .B(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n348), .A2(new_n384), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  AND2_X1   g0237(.A1(G264), .A2(G1698), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n413), .A2(new_n270), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT85), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  XOR2_X1   g0241(.A(KEYINPUT86), .B(G303), .Z(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n273), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n438), .A2(KEYINPUT85), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n214), .B2(G1698), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n390), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n441), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n316), .ZN(new_n448));
  NOR2_X1   g0248(.A1(KEYINPUT80), .A2(G41), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT5), .B1(new_n449), .B2(KEYINPUT67), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n262), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n253), .A2(G45), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(KEYINPUT5), .B2(new_n449), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n451), .A2(new_n453), .B1(new_n250), .B2(new_n251), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G270), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n451), .A2(new_n453), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G274), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n448), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G190), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G283), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n460), .B(new_n229), .C1(G33), .C2(new_n213), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n461), .B(new_n302), .C1(new_n229), .C2(G116), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT87), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT20), .ZN(new_n464));
  XNOR2_X1  g0264(.A(new_n462), .B(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT20), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n465), .B1(KEYINPUT87), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G116), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n306), .A2(G20), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n253), .A2(G33), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n341), .A2(new_n470), .A3(new_n228), .A4(new_n301), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n469), .B1(new_n471), .B2(new_n468), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G200), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n459), .B(new_n473), .C1(new_n474), .C2(new_n458), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n473), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n448), .A2(new_n455), .A3(new_n457), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n477), .A2(G169), .A3(new_n478), .ZN(new_n479));
  XNOR2_X1  g0279(.A(KEYINPUT89), .B(KEYINPUT21), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n390), .B1(G250), .B2(G1698), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(new_n214), .B2(G1698), .ZN(new_n483));
  INV_X1    g0283(.A(G294), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n412), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n316), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n454), .A2(G264), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n486), .A2(new_n457), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n423), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT22), .ZN(new_n491));
  NOR4_X1   g0291(.A1(new_n388), .A2(new_n491), .A3(new_n211), .A4(new_n389), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n412), .A2(new_n468), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n229), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n317), .A2(new_n229), .A3(G87), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n491), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n229), .A2(G107), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n497), .B(KEYINPUT23), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT24), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n494), .A2(KEYINPUT24), .A3(new_n496), .A4(new_n498), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n302), .A3(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n471), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G107), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n306), .A2(new_n497), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n506), .B(KEYINPUT25), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n503), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n488), .A2(new_n325), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n490), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n478), .A2(KEYINPUT21), .A3(G169), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n448), .A2(G179), .A3(new_n455), .A4(new_n457), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT88), .B1(new_n514), .B2(new_n477), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT88), .ZN(new_n516));
  AOI211_X1 g0316(.A(new_n516), .B(new_n473), .C1(new_n512), .C2(new_n513), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n481), .B(new_n511), .C1(new_n515), .C2(new_n517), .ZN(new_n518));
  AOI22_X1  g0318(.A1(G257), .A2(new_n454), .B1(new_n456), .B2(G274), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n323), .A2(G1698), .ZN(new_n520));
  XNOR2_X1  g0320(.A(KEYINPUT75), .B(G33), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n270), .B(new_n520), .C1(new_n521), .C2(new_n269), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT4), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n319), .A2(G244), .ZN(new_n525));
  OAI22_X1  g0325(.A1(new_n525), .A2(new_n523), .B1(new_n212), .B2(new_n319), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n317), .A2(new_n526), .B1(G33), .B2(G283), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n281), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(KEYINPUT79), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT79), .ZN(new_n530));
  AOI211_X1 g0330(.A(new_n530), .B(new_n281), .C1(new_n524), .C2(new_n527), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n423), .B(new_n519), .C1(new_n529), .C2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n528), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n519), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n325), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n341), .A2(G97), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(new_n504), .B2(G97), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT77), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT6), .ZN(new_n541));
  AND2_X1   g0341(.A1(G97), .A2(G107), .ZN(new_n542));
  NOR2_X1   g0342(.A1(G97), .A2(G107), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(G107), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n545), .A2(KEYINPUT6), .A3(G97), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n229), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n334), .A2(new_n298), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n540), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n548), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n545), .A2(KEYINPUT6), .A3(G97), .ZN(new_n551));
  XNOR2_X1  g0351(.A(G97), .B(G107), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n551), .B1(new_n552), .B2(new_n541), .ZN(new_n553));
  OAI211_X1 g0353(.A(KEYINPUT77), .B(new_n550), .C1(new_n553), .C2(new_n229), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT78), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n402), .B2(new_n545), .ZN(new_n557));
  AOI211_X1 g0357(.A(new_n392), .B(G20), .C1(new_n400), .C2(new_n272), .ZN(new_n558));
  OAI211_X1 g0358(.A(KEYINPUT78), .B(G107), .C1(new_n558), .C2(new_n399), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n555), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n539), .B1(new_n560), .B2(new_n302), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n536), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n519), .B1(new_n529), .B2(new_n531), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G200), .ZN(new_n564));
  INV_X1    g0364(.A(new_n534), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G190), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n561), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT81), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT81), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n564), .A2(new_n561), .A3(new_n566), .A4(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n562), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n341), .A2(new_n336), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n471), .A2(new_n211), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n413), .A2(new_n229), .A3(G68), .A4(new_n270), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT19), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n275), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(G20), .B1(new_n276), .B2(KEYINPUT19), .ZN(new_n577));
  NOR3_X1   g0377(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n574), .B(new_n576), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  AOI211_X1 g0379(.A(new_n572), .B(new_n573), .C1(new_n579), .C2(new_n302), .ZN(new_n580));
  AND2_X1   g0380(.A1(G33), .A2(G41), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n452), .B(G250), .C1(new_n581), .C2(new_n228), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n258), .B2(new_n452), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT82), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n582), .B(KEYINPUT82), .C1(new_n258), .C2(new_n452), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n323), .A2(G1698), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(G238), .B2(G1698), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n388), .A2(new_n589), .A3(new_n389), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n316), .B1(new_n590), .B2(new_n493), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n587), .A2(new_n591), .A3(G190), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT84), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n587), .A2(new_n591), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G200), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT84), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n587), .A2(new_n591), .A3(new_n596), .A4(G190), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n580), .A2(new_n593), .A3(new_n595), .A4(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n572), .B1(new_n579), .B2(new_n302), .ZN(new_n599));
  XNOR2_X1  g0399(.A(new_n336), .B(KEYINPUT83), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n504), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n587), .A2(new_n591), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n423), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n594), .A2(new_n325), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n602), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n598), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n489), .A2(G190), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n503), .A2(new_n508), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n488), .A2(G200), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n505), .A4(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n571), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  NOR4_X1   g0412(.A1(new_n437), .A2(new_n476), .A3(new_n518), .A4(new_n612), .ZN(G372));
  NAND2_X1  g0413(.A1(new_n312), .A2(new_n343), .ZN(new_n614));
  XNOR2_X1  g0414(.A(new_n432), .B(KEYINPUT17), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(new_n315), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n427), .A2(new_n428), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n383), .B1(new_n618), .B2(new_n378), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n479), .A2(new_n480), .B1(new_n514), .B2(new_n477), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n612), .B1(new_n511), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT93), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT90), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n536), .B2(new_n561), .ZN(new_n624));
  AOI21_X1  g0424(.A(G169), .B1(new_n533), .B2(new_n519), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n454), .A2(G257), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n457), .ZN(new_n627));
  AND2_X1   g0427(.A1(G250), .A2(G1698), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n520), .B2(KEYINPUT4), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n460), .B1(new_n629), .B2(new_n273), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(new_n523), .B2(new_n522), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n530), .B1(new_n631), .B2(new_n281), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n528), .A2(KEYINPUT79), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n627), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n625), .B1(new_n634), .B2(new_n423), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n560), .A2(new_n302), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n538), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n635), .A2(new_n637), .A3(KEYINPUT90), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n624), .A2(new_n638), .A3(new_n607), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT91), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n640), .B1(new_n639), .B2(new_n641), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT92), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n635), .A2(new_n637), .A3(new_n606), .A4(new_n598), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(new_n641), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n607), .A2(new_n562), .A3(KEYINPUT92), .A4(KEYINPUT26), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n642), .A2(new_n643), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n606), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n622), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n624), .A2(new_n638), .A3(new_n607), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT91), .B1(new_n652), .B2(KEYINPUT26), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n646), .A2(new_n647), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n656), .A2(KEYINPUT93), .A3(new_n606), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n621), .B1(new_n651), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n619), .B1(new_n437), .B2(new_n658), .ZN(G369));
  OAI21_X1  g0459(.A(new_n481), .B1(new_n515), .B2(new_n517), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n306), .A2(new_n229), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT94), .ZN(new_n662));
  OR3_X1    g0462(.A1(new_n661), .A2(new_n662), .A3(KEYINPUT27), .ZN(new_n663));
  INV_X1    g0463(.A(G213), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(new_n661), .B2(KEYINPUT27), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n662), .B1(new_n661), .B2(KEYINPUT27), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n660), .B1(new_n473), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n473), .A2(new_n670), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n476), .B1(new_n620), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  INV_X1    g0476(.A(new_n511), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n509), .A2(new_n669), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n677), .B1(new_n611), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n511), .A2(new_n669), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n680), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n660), .A2(new_n670), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n684), .A2(new_n685), .A3(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n263), .ZN(new_n690));
  INV_X1    g0490(.A(new_n207), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n578), .A2(new_n468), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n692), .A2(new_n253), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT95), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n692), .A2(new_n232), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n694), .A2(new_n695), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT28), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n571), .A2(new_n607), .A3(new_n611), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n518), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n606), .B1(new_n645), .B2(KEYINPUT26), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(KEYINPUT26), .B2(new_n639), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n669), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT29), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n658), .A2(new_n669), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n709), .B1(new_n710), .B2(KEYINPUT29), .ZN(new_n711));
  INV_X1    g0511(.A(new_n518), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n701), .A2(new_n712), .A3(new_n475), .A4(new_n670), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT96), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n513), .A2(new_n714), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n486), .A2(new_n487), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(new_n716), .A3(new_n603), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT30), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n565), .B1(new_n513), .B2(new_n714), .ZN(new_n719));
  OR3_X1    g0519(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n718), .B1(new_n717), .B2(new_n719), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n458), .A2(G179), .A3(new_n603), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(new_n488), .A3(new_n563), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n720), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n669), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n725), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n725), .A2(KEYINPUT31), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n728), .A2(G330), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n711), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n700), .B1(new_n732), .B2(G1), .ZN(G364));
  NOR2_X1   g0533(.A1(new_n305), .A2(G20), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n253), .B1(new_n734), .B2(G45), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n692), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G330), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n674), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n676), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT97), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n674), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n228), .B1(G20), .B2(new_n325), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n229), .A2(G179), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G190), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n751), .B(KEYINPUT100), .Z(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n474), .A2(G190), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n753), .A2(G329), .B1(G283), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT101), .Z(new_n758));
  NOR3_X1   g0558(.A1(new_n345), .A2(G179), .A3(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n229), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n345), .A2(new_n474), .ZN(new_n761));
  NAND2_X1  g0561(.A1(G20), .A2(G179), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G326), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n760), .A2(new_n484), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n758), .A2(new_n317), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n761), .A2(new_n749), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G303), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n763), .A2(new_n750), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT98), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n771), .A2(new_n772), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G311), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n762), .A2(new_n474), .A3(G190), .ZN(new_n778));
  XNOR2_X1  g0578(.A(KEYINPUT33), .B(G317), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n762), .A2(new_n345), .A3(G200), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n778), .A2(new_n779), .B1(new_n780), .B2(G322), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n767), .A2(new_n770), .A3(new_n777), .A4(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n776), .A2(G77), .B1(G58), .B2(new_n780), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n769), .A2(G87), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n756), .A2(G107), .ZN(new_n785));
  AND3_X1   g0585(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n273), .B1(G68), .B2(new_n778), .ZN(new_n787));
  INV_X1    g0587(.A(new_n760), .ZN(new_n788));
  INV_X1    g0588(.A(new_n764), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n788), .A2(G97), .B1(new_n789), .B2(G50), .ZN(new_n790));
  INV_X1    g0590(.A(G159), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n751), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(KEYINPUT99), .B(KEYINPUT32), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n786), .A2(new_n787), .A3(new_n790), .A4(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n748), .B1(new_n782), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n745), .A2(new_n747), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n232), .A2(new_n264), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n390), .A2(new_n691), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n798), .B(new_n799), .C1(new_n248), .C2(new_n264), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n317), .A2(G355), .A3(new_n207), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n800), .B(new_n801), .C1(G116), .C2(new_n207), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n796), .B1(new_n797), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n746), .A2(new_n737), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n742), .A2(new_n804), .ZN(G396));
  INV_X1    g0605(.A(new_n621), .ZN(new_n806));
  AND3_X1   g0606(.A1(new_n656), .A2(KEYINPUT93), .A3(new_n606), .ZN(new_n807));
  AOI21_X1  g0607(.A(KEYINPUT93), .B1(new_n656), .B2(new_n606), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n670), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n343), .A2(new_n670), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n811), .A2(KEYINPUT103), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n342), .A2(new_n669), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n347), .A2(new_n343), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n811), .A2(KEYINPUT103), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n810), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n809), .A2(new_n670), .A3(new_n816), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(new_n729), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n738), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n755), .A2(new_n211), .ZN(new_n823));
  INV_X1    g0623(.A(new_n776), .ZN(new_n824));
  INV_X1    g0624(.A(G311), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n824), .A2(new_n468), .B1(new_n752), .B2(new_n825), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n823), .B(new_n826), .C1(G294), .C2(new_n780), .ZN(new_n827));
  XNOR2_X1  g0627(.A(KEYINPUT102), .B(G283), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n778), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n317), .B1(new_n769), .B2(G107), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n788), .A2(G97), .B1(new_n789), .B2(G303), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n827), .A2(new_n829), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n768), .A2(new_n202), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G143), .A2(new_n780), .B1(new_n778), .B2(G150), .ZN(new_n834));
  INV_X1    g0634(.A(G137), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n834), .B1(new_n835), .B2(new_n764), .C1(new_n824), .C2(new_n791), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT34), .Z(new_n837));
  AOI211_X1 g0637(.A(new_n833), .B(new_n837), .C1(G132), .C2(new_n753), .ZN(new_n838));
  INV_X1    g0638(.A(G58), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n838), .B1(new_n839), .B2(new_n760), .C1(new_n296), .C2(new_n755), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n832), .B1(new_n840), .B2(new_n414), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n747), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n817), .A2(new_n743), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n747), .A2(new_n743), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n298), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n842), .A2(new_n737), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n822), .A2(new_n846), .ZN(G384));
  NAND2_X1  g0647(.A1(new_n728), .A2(new_n436), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT106), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n311), .A2(new_n669), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n312), .A2(new_n315), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n294), .A2(new_n311), .A3(new_n669), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n817), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n726), .A2(new_n727), .A3(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT40), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT38), .ZN(new_n856));
  INV_X1    g0656(.A(new_n667), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n411), .B1(new_n424), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n432), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n411), .A2(new_n857), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n615), .B2(new_n617), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n856), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n394), .A2(new_n396), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n404), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n398), .A2(new_n866), .A3(new_n302), .A4(new_n407), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n410), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n857), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n429), .B2(new_n434), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n868), .A2(new_n424), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(new_n869), .A3(new_n432), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n858), .A2(new_n860), .A3(new_n432), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n871), .A2(new_n876), .A3(KEYINPUT38), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n855), .B1(new_n864), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n854), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n726), .A2(new_n727), .A3(new_n853), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n874), .A2(new_n875), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n869), .B1(new_n615), .B2(new_n617), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n881), .A2(new_n882), .A3(new_n856), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT38), .B1(new_n871), .B2(new_n876), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n855), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n879), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n849), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(G330), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n885), .A2(KEYINPUT39), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n864), .A2(new_n877), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT39), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n312), .A2(new_n669), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  OAI22_X1  g0696(.A1(new_n894), .A2(new_n896), .B1(new_n617), .B2(new_n857), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n851), .A2(new_n852), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n343), .A2(new_n669), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n899), .B1(new_n819), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n856), .B1(new_n881), .B2(new_n882), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n877), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n898), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n889), .B(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n619), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n708), .B1(new_n810), .B2(new_n707), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n908), .B1(new_n909), .B2(new_n436), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT105), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n907), .B(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n253), .B2(new_n734), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n232), .B(G77), .C1(new_n839), .C2(new_n296), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(G50), .B2(new_n296), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n915), .A2(G1), .A3(new_n305), .ZN(new_n916));
  INV_X1    g0716(.A(new_n553), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n468), .B1(new_n917), .B2(KEYINPUT35), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n918), .B(new_n230), .C1(KEYINPUT35), .C2(new_n917), .ZN(new_n919));
  XOR2_X1   g0719(.A(KEYINPUT104), .B(KEYINPUT36), .Z(new_n920));
  XNOR2_X1  g0720(.A(new_n919), .B(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n913), .A2(new_n916), .A3(new_n921), .ZN(G367));
  INV_X1    g0722(.A(new_n778), .ZN(new_n923));
  INV_X1    g0723(.A(G317), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n923), .A2(new_n484), .B1(new_n751), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n768), .A2(new_n468), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n926), .A2(KEYINPUT46), .B1(new_n213), .B2(new_n755), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n925), .B(new_n927), .C1(KEYINPUT46), .C2(new_n926), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n776), .A2(new_n828), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n789), .A2(G311), .B1(new_n442), .B2(new_n780), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n390), .B1(G107), .B2(new_n788), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n928), .A2(new_n929), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n755), .A2(new_n298), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n760), .A2(new_n296), .ZN(new_n934));
  INV_X1    g0734(.A(new_n780), .ZN(new_n935));
  INV_X1    g0735(.A(G150), .ZN(new_n936));
  INV_X1    g0736(.A(G143), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n935), .A2(new_n936), .B1(new_n764), .B2(new_n937), .ZN(new_n938));
  AOI211_X1 g0738(.A(new_n934), .B(new_n938), .C1(G58), .C2(new_n769), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n273), .B1(new_n776), .B2(G50), .ZN(new_n940));
  INV_X1    g0740(.A(new_n751), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n941), .A2(G137), .B1(G159), .B2(new_n778), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n939), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n932), .B1(new_n933), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT47), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n747), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n607), .B1(new_n580), .B2(new_n670), .ZN(new_n947));
  OR3_X1    g0747(.A1(new_n606), .A2(new_n580), .A3(new_n670), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(new_n745), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n799), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n797), .B1(new_n207), .B2(new_n337), .C1(new_n950), .C2(new_n241), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n946), .A2(new_n737), .A3(new_n949), .A4(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n681), .B(new_n687), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n683), .B1(new_n953), .B2(new_n676), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n731), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n571), .B1(new_n561), .B2(new_n670), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n562), .A2(new_n669), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n688), .B2(new_n685), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT44), .Z(new_n961));
  NAND3_X1  g0761(.A1(new_n688), .A2(new_n685), .A3(new_n959), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT45), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n956), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n732), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n692), .B(KEYINPUT41), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n736), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n681), .A2(new_n571), .A3(new_n687), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n969), .A2(KEYINPUT42), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n957), .A2(new_n511), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n670), .B1(new_n971), .B2(new_n562), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n969), .A2(KEYINPUT42), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n947), .A2(new_n948), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n977), .A2(new_n978), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n683), .A2(new_n959), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n982), .B(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n952), .B1(new_n968), .B2(new_n984), .ZN(G387));
  INV_X1    g0785(.A(new_n692), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(new_n731), .B2(new_n955), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n731), .B2(new_n955), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n789), .A2(G322), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n989), .B1(new_n825), .B2(new_n923), .C1(new_n924), .C2(new_n935), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(new_n442), .B2(new_n776), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT48), .Z(new_n992));
  INV_X1    g0792(.A(new_n828), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n992), .B1(new_n484), .B2(new_n768), .C1(new_n760), .C2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT110), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT49), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n414), .B1(new_n468), .B2(new_n755), .C1(new_n765), .C2(new_n751), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT111), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n776), .A2(G68), .B1(new_n352), .B2(new_n778), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT109), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n600), .A2(new_n788), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n764), .A2(new_n791), .B1(new_n768), .B2(new_n298), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n935), .A2(new_n202), .B1(new_n755), .B2(new_n213), .ZN(new_n1004));
  NOR4_X1   g0804(.A1(new_n1002), .A2(new_n414), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1001), .B(new_n1005), .C1(new_n936), .C2(new_n751), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n748), .B1(new_n999), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n333), .A2(new_n1008), .A3(G50), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1009), .A2(new_n693), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1008), .B1(new_n333), .B2(G50), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1010), .A2(new_n264), .A3(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n296), .A2(new_n298), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n799), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT108), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n238), .A2(new_n264), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1015), .A2(new_n1016), .B1(new_n545), .B2(new_n691), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n317), .A2(new_n693), .A3(new_n207), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n738), .B(new_n1007), .C1(new_n797), .C2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n682), .A2(new_n745), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1020), .A2(new_n1021), .B1(new_n736), .B2(new_n954), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n988), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT112), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n988), .A2(KEYINPUT112), .A3(new_n1022), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(G393));
  XNOR2_X1  g0827(.A(new_n964), .B(new_n684), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n692), .B(new_n965), .C1(new_n1028), .C2(new_n956), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n736), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n957), .A2(new_n745), .A3(new_n958), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n797), .B1(new_n213), .B2(new_n207), .C1(new_n950), .C2(new_n245), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n789), .A2(G317), .B1(G311), .B2(new_n780), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT52), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n442), .B2(new_n778), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n941), .A2(G322), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n776), .A2(G294), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n785), .B1(new_n768), .B2(new_n993), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n317), .B(new_n1038), .C1(G116), .C2(new_n788), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n789), .A2(G150), .B1(G159), .B2(new_n780), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT51), .Z(new_n1042));
  AOI22_X1  g0842(.A1(new_n941), .A2(G143), .B1(G50), .B2(new_n778), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n823), .B1(G77), .B2(new_n788), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n414), .B1(G68), .B2(new_n769), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n824), .A2(new_n333), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1040), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n747), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1031), .A2(new_n737), .A3(new_n1032), .A4(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1029), .A2(new_n1030), .A3(new_n1050), .ZN(G390));
  NAND4_X1  g0851(.A1(new_n726), .A2(new_n853), .A3(new_n727), .A4(G330), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n894), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n899), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n658), .A2(new_n669), .A3(new_n817), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1055), .B1(new_n1056), .B2(new_n900), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1054), .B1(new_n1057), .B2(new_n896), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n900), .B1(new_n705), .B2(new_n816), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n896), .B(new_n891), .C1(new_n1059), .C2(new_n899), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1053), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n894), .B1(new_n902), .B2(new_n895), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1063), .A2(new_n1060), .A3(new_n1052), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n736), .A3(new_n1064), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n776), .A2(G97), .B1(G107), .B2(new_n778), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT113), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n784), .B1(new_n468), .B2(new_n935), .C1(new_n298), .C2(new_n760), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G68), .B2(new_n756), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n753), .A2(G294), .B1(G283), .B2(new_n789), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1067), .A2(new_n273), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  NOR3_X1   g0871(.A1(new_n768), .A2(KEYINPUT53), .A3(new_n936), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT53), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n769), .B2(G150), .ZN(new_n1074));
  INV_X1    g0874(.A(G128), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n764), .A2(new_n1075), .B1(new_n755), .B2(new_n202), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1074), .B(new_n1076), .C1(new_n753), .C2(G125), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n788), .A2(G159), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G132), .A2(new_n780), .B1(new_n778), .B2(G137), .ZN(new_n1079));
  XOR2_X1   g0879(.A(KEYINPUT54), .B(G143), .Z(new_n1080));
  AOI21_X1  g0880(.A(new_n273), .B1(new_n776), .B2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .A4(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1071), .B1(new_n1072), .B2(new_n1082), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT114), .Z(new_n1084));
  AOI22_X1  g0884(.A1(new_n894), .A2(new_n743), .B1(new_n747), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n844), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1085), .B(new_n737), .C1(new_n352), .C2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(KEYINPUT115), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1065), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n726), .A2(new_n727), .A3(G330), .A4(new_n816), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n899), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1091), .A2(new_n1059), .A3(new_n1052), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1056), .A2(new_n900), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1053), .B1(new_n899), .B2(new_n1090), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1092), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n728), .A2(G330), .A3(new_n436), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1095), .A2(new_n910), .A3(new_n1096), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n1063), .A2(new_n1060), .A3(new_n1052), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1052), .B1(new_n1063), .B2(new_n1060), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n819), .A2(new_n901), .B1(new_n1091), .B2(new_n1052), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1092), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n619), .B(new_n1096), .C1(new_n711), .C2(new_n437), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1062), .A2(new_n1064), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1100), .A2(new_n692), .A3(new_n1106), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n1087), .A2(KEYINPUT115), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1089), .A2(new_n1107), .A3(new_n1108), .ZN(G378));
  NAND2_X1  g0909(.A1(new_n380), .A2(new_n857), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n383), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1110), .B1(new_n378), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n378), .A2(new_n1111), .A3(new_n1110), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1115), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1110), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n383), .B(new_n1118), .C1(new_n373), .C2(new_n377), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1117), .B1(new_n1112), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1116), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n904), .A2(new_n726), .A3(new_n727), .A4(new_n853), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1122), .A2(new_n855), .B1(new_n854), .B2(new_n878), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1121), .B1(new_n1123), .B2(G330), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT118), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1116), .A2(new_n1120), .A3(KEYINPUT118), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AND4_X1   g0928(.A1(G330), .A2(new_n879), .A3(new_n1128), .A4(new_n886), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n905), .B(new_n898), .C1(new_n1124), .C2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1121), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n887), .B2(new_n739), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1123), .A2(G330), .A3(new_n1128), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n885), .B(new_n899), .C1(new_n819), .C2(new_n901), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1132), .B(new_n1133), .C1(new_n1134), .C2(new_n897), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1130), .A2(new_n1135), .A3(new_n736), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1126), .A2(new_n743), .A3(new_n1127), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n844), .A2(new_n202), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n768), .A2(new_n298), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n935), .A2(new_n545), .B1(new_n755), .B2(new_n839), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1139), .B(new_n1140), .C1(G116), .C2(new_n789), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n753), .A2(G283), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n414), .A2(new_n263), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n776), .B2(new_n600), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n934), .B1(G97), .B2(new_n778), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1141), .A2(new_n1142), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT58), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1143), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(G159), .A2(new_n756), .B1(new_n941), .B2(G124), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1149), .A2(new_n271), .A3(new_n259), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n776), .A2(G137), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n780), .A2(G128), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n789), .A2(G125), .B1(new_n769), .B2(new_n1080), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n788), .A2(G150), .B1(new_n778), .B2(G132), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  XOR2_X1   g0955(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n1156));
  XNOR2_X1  g0956(.A(new_n1155), .B(new_n1156), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1147), .B(new_n1148), .C1(new_n1150), .C2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT117), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n747), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1137), .A2(new_n737), .A3(new_n1138), .A4(new_n1160), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1136), .A2(KEYINPUT119), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(KEYINPUT119), .B1(new_n1136), .B2(new_n1161), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1104), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1106), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1130), .A2(new_n1135), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT57), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n1130), .A2(new_n1135), .A3(KEYINPUT57), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n986), .B1(new_n1166), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1164), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT120), .ZN(G375));
  NAND2_X1  g0975(.A1(new_n899), .A2(new_n743), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n317), .B1(G283), .B2(new_n780), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n298), .B2(new_n755), .C1(new_n468), .C2(new_n923), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1002), .B1(G294), .B2(new_n789), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n753), .A2(G303), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(new_n213), .C2(new_n768), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1178), .B(new_n1181), .C1(G107), .C2(new_n776), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n390), .B1(new_n835), .B2(new_n935), .C1(new_n824), .C2(new_n936), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n760), .A2(new_n202), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n752), .A2(new_n1075), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n769), .A2(G159), .B1(new_n789), .B2(G132), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n756), .A2(G58), .B1(new_n1080), .B2(new_n778), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NOR4_X1   g0988(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .A4(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n747), .B1(new_n1182), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n844), .A2(new_n296), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1176), .A2(new_n737), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n1103), .B2(new_n735), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n967), .B1(new_n1165), .B2(new_n1095), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1194), .B1(new_n1195), .B2(new_n1105), .ZN(G381));
  NOR2_X1   g0996(.A1(G375), .A2(G378), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(G387), .A2(G390), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(G381), .A2(G384), .ZN(new_n1199));
  INV_X1    g0999(.A(G396), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1025), .A2(new_n1200), .A3(new_n1026), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1198), .A2(new_n1199), .A3(new_n1202), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1203), .A2(KEYINPUT121), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(KEYINPUT121), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1197), .A2(new_n1204), .A3(new_n1205), .ZN(G407));
  AOI21_X1  g1006(.A(new_n664), .B1(new_n1197), .B2(new_n668), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(G407), .ZN(G409));
  INV_X1    g1008(.A(KEYINPUT123), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1136), .A2(new_n1161), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1167), .B1(new_n1106), .B2(new_n1165), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n1211), .B2(new_n967), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1209), .B1(new_n1212), .B2(G378), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1166), .A2(new_n967), .A3(new_n1168), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1210), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1065), .A2(new_n1108), .A3(new_n1088), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n1106), .A2(new_n692), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1217), .B1(new_n1218), .B2(new_n1100), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1216), .A2(new_n1219), .A3(KEYINPUT123), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1213), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT122), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n1174), .B2(G378), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n1098), .A2(new_n1099), .A3(new_n1097), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1172), .B1(new_n1224), .B2(new_n1104), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1225), .B(new_n692), .C1(KEYINPUT57), .C2(new_n1211), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1227));
  AND4_X1   g1027(.A1(new_n1222), .A2(new_n1226), .A3(G378), .A4(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1221), .B1(new_n1223), .B2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1103), .A2(new_n1104), .A3(KEYINPUT60), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1230), .A2(new_n692), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT60), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(new_n1105), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT124), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1231), .A2(new_n1233), .A3(KEYINPUT124), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(G384), .B1(new_n1238), .B2(new_n1194), .ZN(new_n1239));
  INV_X1    g1039(.A(G384), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1240), .B(new_n1193), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n664), .A2(G343), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1229), .A2(new_n1242), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(KEYINPUT62), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(G387), .B(G390), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT126), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(G393), .A2(G396), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1249), .B1(new_n1250), .B2(new_n1201), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(new_n1249), .A3(new_n1201), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1248), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1253), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1247), .B1(new_n1255), .B2(new_n1251), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT127), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1257), .A2(KEYINPUT61), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1254), .A2(new_n1256), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(KEYINPUT61), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT62), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1229), .A2(new_n1242), .A3(new_n1262), .A4(new_n1244), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1246), .A2(new_n1261), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT125), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  OAI211_X1 g1067(.A(G2897), .B(new_n1243), .C1(new_n1239), .C2(new_n1241), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1238), .A2(new_n1194), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1240), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1238), .A2(G384), .A3(new_n1194), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1243), .A2(G2897), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1268), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1213), .A2(new_n1220), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1174), .A2(G378), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(KEYINPUT122), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1174), .A2(new_n1222), .A3(G378), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1275), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1274), .B1(new_n1279), .B2(new_n1243), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1245), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT125), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1274), .B(new_n1283), .C1(new_n1279), .C2(new_n1243), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1229), .A2(new_n1242), .A3(KEYINPUT63), .A4(new_n1244), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1282), .A2(new_n1284), .A3(new_n1285), .A4(new_n1286), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1267), .A2(new_n1280), .B1(new_n1265), .B2(new_n1287), .ZN(G405));
  NAND2_X1  g1088(.A1(G375), .A2(new_n1219), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1242), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1289), .B(new_n1290), .C1(new_n1239), .C2(new_n1241), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1265), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1294), .B(new_n1295), .ZN(G402));
endmodule


