//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n206));
  INV_X1    g0006(.A(G68), .ZN(new_n207));
  INV_X1    g0007(.A(G238), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n212));
  INV_X1    g0012(.A(G77), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  INV_X1    g0014(.A(G107), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n205), .B1(new_n211), .B2(new_n217), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT64), .Z(new_n219));
  INV_X1    g0019(.A(KEYINPUT1), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT65), .Z(new_n222));
  NAND2_X1  g0022(.A1(new_n202), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  AND2_X1   g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n205), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT0), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n229), .B(new_n232), .C1(new_n219), .C2(new_n220), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n222), .A2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  OAI21_X1  g0050(.A(KEYINPUT68), .B1(new_n205), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT68), .ZN(new_n252));
  NAND4_X1  g0052(.A1(new_n252), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G13), .A3(G20), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n251), .A2(new_n226), .A3(new_n253), .A4(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(G20), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G50), .ZN(new_n258));
  OAI22_X1  g0058(.A1(new_n256), .A2(new_n258), .B1(G50), .B2(new_n255), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n259), .B(KEYINPUT69), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n226), .A2(new_n253), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n251), .ZN(new_n262));
  INV_X1    g0062(.A(G50), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n227), .B1(new_n201), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT8), .B(G58), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n227), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(G150), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  OAI22_X1  g0069(.A1(new_n265), .A2(new_n266), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n262), .B1(new_n264), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n260), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n272), .B(KEYINPUT9), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(G222), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(G1698), .ZN(new_n277));
  INV_X1    g0077(.A(G223), .ZN(new_n278));
  OAI221_X1 g0078(.A(new_n276), .B1(new_n213), .B2(new_n274), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n225), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(new_n281), .B(KEYINPUT67), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G41), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT66), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT66), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G41), .ZN(new_n287));
  INV_X1    g0087(.A(G45), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G274), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(new_n225), .B2(new_n280), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(new_n291), .A3(new_n254), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n284), .A2(new_n288), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n254), .A2(new_n293), .B1(new_n225), .B2(new_n280), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G226), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n283), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(G200), .B2(new_n296), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n273), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT10), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n274), .A2(G232), .A3(G1698), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n274), .A2(G226), .A3(new_n275), .ZN(new_n303));
  INV_X1    g0103(.A(G97), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n302), .B(new_n303), .C1(new_n250), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n282), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT71), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n208), .B1(new_n294), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(new_n307), .B2(new_n294), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(new_n292), .A3(new_n309), .ZN(new_n310));
  OR2_X1    g0110(.A1(new_n310), .A2(KEYINPUT13), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(KEYINPUT13), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G169), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT14), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n312), .A2(KEYINPUT72), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n312), .A2(KEYINPUT72), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n316), .A2(G179), .A3(new_n317), .A4(new_n311), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT14), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n313), .A2(new_n319), .A3(G169), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n315), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n255), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n207), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n323), .B(KEYINPUT12), .ZN(new_n324));
  INV_X1    g0124(.A(new_n256), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(G68), .A3(new_n257), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n327), .A2(KEYINPUT74), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n268), .A2(G50), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT73), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n266), .A2(new_n213), .B1(new_n227), .B2(G68), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n262), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT11), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n327), .A2(KEYINPUT74), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n328), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n321), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n335), .B1(new_n313), .B2(G200), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n316), .A2(G190), .A3(new_n317), .A4(new_n311), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G179), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n274), .A2(G232), .A3(new_n275), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT3), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G33), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G107), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n341), .B(new_n346), .C1(new_n277), .C2(new_n208), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n282), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n294), .A2(G244), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n349), .A2(new_n292), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n348), .A2(KEYINPUT70), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT70), .B1(new_n348), .B2(new_n350), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n340), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n348), .A2(new_n350), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT70), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G169), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n357), .A2(new_n358), .A3(new_n351), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT15), .B(G87), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(new_n266), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n265), .A2(new_n269), .B1(new_n227), .B2(new_n213), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n262), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n325), .A2(G77), .A3(new_n257), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n322), .A2(new_n213), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n354), .A2(new_n359), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(G190), .B1(new_n352), .B2(new_n353), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n357), .A2(G200), .A3(new_n351), .ZN(new_n369));
  INV_X1    g0169(.A(new_n366), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n296), .A2(new_n358), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n372), .B(new_n272), .C1(G179), .C2(new_n296), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n367), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n301), .A2(new_n336), .A3(new_n339), .A4(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G58), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n376), .A2(new_n207), .ZN(new_n377));
  OAI21_X1  g0177(.A(G20), .B1(new_n377), .B2(new_n201), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n268), .A2(G159), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT7), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(new_n274), .B2(G20), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT75), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n343), .A2(G33), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n386));
  OAI211_X1 g0186(.A(KEYINPUT7), .B(new_n227), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  AND3_X1   g0187(.A1(new_n383), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  OAI211_X1 g0188(.A(KEYINPUT75), .B(new_n382), .C1(new_n274), .C2(G20), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G68), .ZN(new_n390));
  OAI211_X1 g0190(.A(KEYINPUT16), .B(new_n381), .C1(new_n388), .C2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT16), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n207), .B1(new_n383), .B2(new_n387), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n392), .B1(new_n393), .B2(new_n380), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n391), .A2(new_n262), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n265), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n257), .ZN(new_n397));
  OAI22_X1  g0197(.A1(new_n397), .A2(new_n256), .B1(new_n396), .B2(new_n255), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT76), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI221_X1 g0200(.A(KEYINPUT76), .B1(new_n396), .B2(new_n255), .C1(new_n397), .C2(new_n256), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n342), .A2(new_n344), .A3(G226), .A4(G1698), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n342), .A2(new_n344), .A3(G223), .A4(new_n275), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n404), .B(new_n405), .C1(new_n250), .C2(new_n209), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n282), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n293), .A2(new_n254), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(G232), .A3(new_n281), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n292), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n407), .A2(new_n410), .A3(new_n297), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n292), .A2(new_n409), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n282), .B2(new_n406), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n411), .B1(new_n413), .B2(G200), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n395), .A2(new_n403), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT17), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(KEYINPUT79), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT79), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n415), .B2(KEYINPUT17), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT78), .ZN(new_n423));
  INV_X1    g0223(.A(new_n262), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT7), .B1(new_n345), .B2(new_n227), .ZN(new_n425));
  AOI211_X1 g0225(.A(new_n382), .B(G20), .C1(new_n342), .C2(new_n344), .ZN(new_n426));
  OAI21_X1  g0226(.A(G68), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n381), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n424), .B1(new_n428), .B2(new_n392), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n402), .B1(new_n429), .B2(new_n391), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n423), .B1(new_n430), .B2(new_n414), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n395), .A2(new_n403), .A3(new_n414), .A4(new_n423), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT17), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n422), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n395), .A2(new_n403), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT77), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n430), .A2(KEYINPUT77), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n413), .A2(new_n358), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n441), .B1(G179), .B2(new_n413), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n439), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT18), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n439), .A2(new_n440), .A3(new_n443), .A4(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n436), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n375), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n274), .A2(new_n227), .A3(G68), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT19), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n266), .B2(new_n304), .ZN(new_n452));
  NAND3_X1  g0252(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n227), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT82), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n209), .A2(new_n304), .A3(new_n215), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n454), .A2(KEYINPUT82), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n450), .B(new_n452), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n262), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n254), .A2(G33), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n261), .A2(new_n251), .A3(new_n255), .A4(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT83), .B1(new_n462), .B2(new_n360), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT83), .ZN(new_n464));
  INV_X1    g0264(.A(new_n360), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n325), .A2(new_n464), .A3(new_n465), .A4(new_n461), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n360), .A2(new_n322), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n460), .A2(new_n463), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n254), .A2(new_n290), .A3(G45), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n210), .B1(new_n288), .B2(G1), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n281), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT67), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n281), .B(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G116), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(G238), .A2(G1698), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n214), .B2(G1698), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n475), .B1(new_n477), .B2(new_n274), .ZN(new_n478));
  OAI211_X1 g0278(.A(G179), .B(new_n471), .C1(new_n473), .C2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n471), .ZN(new_n480));
  INV_X1    g0280(.A(new_n478), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n480), .B1(new_n481), .B2(new_n282), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n479), .B1(new_n482), .B2(new_n358), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n468), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n459), .A2(new_n262), .B1(new_n322), .B2(new_n360), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n471), .B1(new_n473), .B2(new_n478), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G200), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n256), .B1(new_n254), .B2(G33), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G87), .ZN(new_n489));
  OAI211_X1 g0289(.A(G190), .B(new_n471), .C1(new_n473), .C2(new_n478), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n485), .A2(new_n487), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n484), .A2(KEYINPUT84), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT84), .B1(new_n484), .B2(new_n491), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n274), .A2(G257), .A3(G1698), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G294), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n342), .A2(new_n344), .A3(G250), .A4(new_n275), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT86), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n282), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT5), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n254), .B(G45), .C1(new_n501), .C2(G41), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n285), .A2(new_n287), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(new_n501), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n291), .ZN(new_n505));
  XNOR2_X1  g0305(.A(KEYINPUT66), .B(G41), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n507));
  OAI211_X1 g0307(.A(G264), .B(new_n281), .C1(new_n507), .C2(new_n502), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n500), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n499), .B1(new_n498), .B2(new_n282), .ZN(new_n510));
  OAI21_X1  g0310(.A(G169), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n498), .A2(new_n282), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(new_n505), .A3(new_n508), .ZN(new_n513));
  OR2_X1    g0313(.A1(new_n513), .A2(new_n340), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n274), .A2(new_n227), .A3(G87), .ZN(new_n516));
  XNOR2_X1  g0316(.A(KEYINPUT85), .B(KEYINPUT22), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n274), .A2(new_n517), .A3(new_n227), .A4(G87), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT24), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT23), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n227), .B2(G107), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n215), .A2(KEYINPUT23), .A3(G20), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n524), .A2(new_n525), .B1(new_n475), .B2(new_n227), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n521), .A2(new_n522), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n522), .B1(new_n521), .B2(new_n526), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n262), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n322), .A2(new_n215), .ZN(new_n530));
  XNOR2_X1  g0330(.A(new_n530), .B(KEYINPUT25), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(G107), .B2(new_n488), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n515), .A2(new_n533), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n509), .A2(G190), .A3(new_n510), .ZN(new_n535));
  INV_X1    g0335(.A(G200), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n513), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n529), .B(new_n532), .C1(new_n535), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n494), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n488), .A2(G116), .ZN(new_n541));
  INV_X1    g0341(.A(G116), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n322), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(G20), .B1(G33), .B2(G283), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n250), .A2(G97), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n544), .A2(new_n545), .B1(G20), .B2(new_n542), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n262), .A2(KEYINPUT20), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT20), .B1(new_n262), .B2(new_n546), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n541), .B(new_n543), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(G270), .B(new_n281), .C1(new_n507), .C2(new_n502), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n550), .A2(new_n505), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n274), .A2(G257), .A3(new_n275), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n345), .A2(G303), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n552), .B(new_n553), .C1(new_n277), .C2(new_n216), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n282), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n549), .A2(new_n556), .A3(KEYINPUT21), .A4(G169), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n549), .A2(G179), .A3(new_n555), .A4(new_n551), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n549), .A2(new_n556), .A3(G169), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT21), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n556), .A2(G200), .ZN(new_n563));
  INV_X1    g0363(.A(new_n549), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n563), .B(new_n564), .C1(new_n297), .C2(new_n556), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n559), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n268), .A2(G77), .ZN(new_n567));
  XNOR2_X1  g0367(.A(G97), .B(G107), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT80), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n568), .B1(new_n569), .B2(KEYINPUT6), .ZN(new_n570));
  MUX2_X1   g0370(.A(new_n569), .B(G97), .S(KEYINPUT6), .Z(new_n571));
  OAI21_X1  g0371(.A(new_n570), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n567), .B1(new_n572), .B2(new_n227), .ZN(new_n573));
  OAI21_X1  g0373(.A(G107), .B1(new_n425), .B2(new_n426), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n262), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n488), .A2(G97), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n255), .A2(G97), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n274), .A2(G244), .A3(new_n275), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT4), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(G33), .A2(G283), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n274), .A2(KEYINPUT4), .A3(G244), .A4(new_n275), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n274), .A2(G250), .A3(G1698), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n583), .A2(new_n584), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n282), .ZN(new_n588));
  OAI211_X1 g0388(.A(G257), .B(new_n281), .C1(new_n507), .C2(new_n502), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n589), .A2(new_n505), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n358), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n588), .A2(new_n590), .A3(new_n340), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n580), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n591), .A2(G200), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n574), .B(new_n567), .C1(new_n227), .C2(new_n572), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n578), .B1(new_n596), .B2(new_n262), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n588), .A2(new_n590), .A3(G190), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n595), .A2(new_n597), .A3(new_n577), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT81), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n594), .A2(new_n599), .A3(KEYINPUT81), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AND4_X1   g0404(.A1(new_n449), .A2(new_n540), .A3(new_n566), .A4(new_n604), .ZN(G372));
  XOR2_X1   g0405(.A(new_n300), .B(KEYINPUT10), .Z(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT87), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT87), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n301), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n442), .A2(new_n430), .ZN(new_n611));
  XNOR2_X1  g0411(.A(new_n611), .B(new_n446), .ZN(new_n612));
  INV_X1    g0412(.A(new_n339), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n336), .B1(new_n613), .B2(new_n367), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n612), .B1(new_n614), .B2(new_n436), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n373), .B1(new_n610), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n449), .ZN(new_n618));
  INV_X1    g0418(.A(new_n594), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n484), .A2(new_n491), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n600), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n623), .A2(new_n491), .A3(new_n538), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n559), .A2(new_n534), .A3(new_n562), .ZN(new_n625));
  OAI221_X1 g0425(.A(new_n484), .B1(KEYINPUT26), .B2(new_n622), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  INV_X1    g0427(.A(new_n494), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n627), .B1(new_n628), .B2(new_n619), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n617), .B1(new_n618), .B2(new_n630), .ZN(G369));
  NAND3_X1  g0431(.A1(new_n254), .A2(new_n227), .A3(G13), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(G213), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(G343), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n549), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n566), .A2(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n559), .A2(new_n562), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n639), .B1(new_n640), .B2(new_n638), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n641), .A2(G330), .ZN(new_n642));
  INV_X1    g0442(.A(new_n539), .ZN(new_n643));
  INV_X1    g0443(.A(new_n533), .ZN(new_n644));
  INV_X1    g0444(.A(new_n637), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n534), .B2(new_n645), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n534), .A2(new_n637), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n640), .A2(new_n637), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n650), .B1(new_n651), .B2(new_n643), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n649), .A2(new_n652), .ZN(G399));
  OR2_X1    g0453(.A1(new_n456), .A2(G116), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n654), .B(KEYINPUT88), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n506), .A2(new_n230), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(G1), .ZN(new_n657));
  OAI22_X1  g0457(.A1(new_n655), .A2(new_n657), .B1(new_n223), .B2(new_n656), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT28), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT29), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n660), .B(new_n645), .C1(new_n626), .C2(new_n629), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n622), .A2(KEYINPUT26), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n484), .B(new_n662), .C1(new_n624), .C2(new_n625), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n628), .A2(new_n627), .A3(new_n619), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n637), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n661), .B1(new_n666), .B2(new_n660), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT92), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n512), .A2(new_n508), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT90), .B1(new_n669), .B2(new_n486), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT90), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n482), .A2(new_n671), .A3(new_n512), .A4(new_n508), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n591), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n555), .A2(G179), .A3(new_n505), .A4(new_n550), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT91), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT91), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n551), .A2(new_n676), .A3(G179), .A4(new_n555), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n668), .B1(new_n673), .B2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT30), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n673), .A2(new_n678), .A3(new_n668), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n673), .A2(new_n678), .A3(KEYINPUT30), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n482), .A2(G179), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n591), .A2(new_n556), .A3(new_n513), .A4(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n683), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g0487(.A(KEYINPUT89), .B(KEYINPUT31), .Z(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n687), .A2(new_n637), .A3(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n604), .A2(new_n540), .A3(new_n566), .A4(new_n645), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n556), .A2(new_n685), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT93), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n692), .A2(new_n693), .A3(new_n513), .A4(new_n591), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n686), .A2(KEYINPUT93), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n696), .A2(new_n684), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n645), .B1(new_n697), .B2(new_n683), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n690), .B(new_n691), .C1(KEYINPUT31), .C2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n667), .B1(G330), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n659), .B1(new_n700), .B2(G1), .ZN(G364));
  NAND3_X1  g0501(.A1(new_n227), .A2(G13), .A3(G45), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT94), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(KEYINPUT94), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G1), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n656), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n642), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(G330), .B2(new_n641), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n274), .A2(new_n230), .ZN(new_n711));
  INV_X1    g0511(.A(G355), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n711), .A2(new_n712), .B1(G116), .B2(new_n230), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n245), .A2(new_n288), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n345), .A2(new_n230), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(new_n288), .B2(new_n224), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n713), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n226), .B1(G20), .B2(new_n358), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n718), .A2(KEYINPUT95), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(KEYINPUT95), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G13), .A2(G33), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G20), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n717), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n707), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n227), .A2(G179), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(G190), .A3(G200), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n209), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n227), .A2(new_n340), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G190), .A2(G200), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n732), .A2(G190), .A3(new_n536), .ZN(new_n735));
  OAI221_X1 g0535(.A(new_n274), .B1(new_n734), .B2(new_n213), .C1(new_n376), .C2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n732), .A2(G200), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n297), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n731), .B(new_n736), .C1(G50), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n737), .A2(G190), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n729), .A2(new_n297), .A3(G200), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n741), .A2(new_n207), .B1(new_n742), .B2(new_n215), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n297), .A2(G179), .A3(G200), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n227), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n743), .B1(G97), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n729), .A2(new_n733), .ZN(new_n748));
  INV_X1    g0548(.A(G159), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT32), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n739), .A2(new_n747), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT96), .ZN(new_n753));
  INV_X1    g0553(.A(G311), .ZN(new_n754));
  INV_X1    g0554(.A(G322), .ZN(new_n755));
  OAI221_X1 g0555(.A(new_n345), .B1(new_n734), .B2(new_n754), .C1(new_n755), .C2(new_n735), .ZN(new_n756));
  XOR2_X1   g0556(.A(KEYINPUT33), .B(G317), .Z(new_n757));
  NOR2_X1   g0557(.A1(new_n741), .A2(new_n757), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n756), .B(new_n758), .C1(G326), .C2(new_n738), .ZN(new_n759));
  INV_X1    g0559(.A(G294), .ZN(new_n760));
  INV_X1    g0560(.A(G303), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n745), .A2(new_n760), .B1(new_n730), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n742), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n762), .B1(G283), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n748), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT97), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(KEYINPUT97), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G329), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n759), .A2(new_n764), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n753), .A2(new_n771), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n772), .A2(KEYINPUT98), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n721), .B1(new_n772), .B2(KEYINPUT98), .ZN(new_n774));
  INV_X1    g0574(.A(new_n724), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n728), .B1(new_n773), .B2(new_n774), .C1(new_n641), .C2(new_n775), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n710), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(G396));
  NOR2_X1   g0578(.A1(new_n630), .A2(new_n637), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT101), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n366), .A2(new_n637), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n367), .A2(new_n371), .A3(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT99), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n367), .A2(new_n371), .A3(KEYINPUT99), .A4(new_n781), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n354), .A2(new_n359), .A3(new_n366), .A4(new_n637), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT100), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n780), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n786), .A2(new_n780), .A3(new_n788), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n779), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n699), .A2(G330), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n708), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n794), .B2(new_n793), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n721), .A2(new_n722), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n708), .B1(new_n798), .B2(G77), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n769), .A2(G311), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n209), .A2(new_n742), .B1(new_n730), .B2(new_n215), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(G283), .B2(new_n740), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n345), .B1(new_n734), .B2(new_n542), .ZN(new_n803));
  INV_X1    g0603(.A(new_n735), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n803), .B1(G294), .B2(new_n804), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G97), .A2(new_n746), .B1(new_n738), .B2(G303), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n800), .A2(new_n802), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n734), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n804), .A2(G143), .B1(new_n808), .B2(G159), .ZN(new_n809));
  INV_X1    g0609(.A(new_n738), .ZN(new_n810));
  INV_X1    g0610(.A(G137), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n809), .B1(new_n810), .B2(new_n811), .C1(new_n267), .C2(new_n741), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT34), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n263), .A2(new_n730), .B1(new_n742), .B2(new_n207), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n345), .B(new_n815), .C1(G58), .C2(new_n746), .ZN(new_n816));
  INV_X1    g0616(.A(G132), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n814), .B(new_n816), .C1(new_n817), .C2(new_n768), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n812), .A2(new_n813), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n807), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n799), .B1(new_n820), .B2(new_n721), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n792), .B2(new_n723), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n796), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G384));
  INV_X1    g0624(.A(KEYINPUT35), .ZN(new_n825));
  OAI211_X1 g0625(.A(G116), .B(new_n228), .C1(new_n572), .C2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n825), .B2(new_n572), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT36), .ZN(new_n828));
  OR3_X1    g0628(.A1(new_n223), .A2(new_n213), .A3(new_n377), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n263), .A2(G68), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n254), .B(G13), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n391), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n384), .A2(KEYINPUT7), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n207), .B1(new_n425), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n383), .A2(new_n384), .A3(new_n387), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n380), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n262), .B1(new_n837), .B2(KEYINPUT16), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT102), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n833), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI211_X1 g0640(.A(KEYINPUT102), .B(new_n262), .C1(new_n837), .C2(KEYINPUT16), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n398), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(new_n635), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n415), .A2(KEYINPUT78), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n432), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n845), .A2(new_n417), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(new_n421), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n445), .A2(new_n447), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n843), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(KEYINPUT38), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT37), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n844), .B(new_n432), .C1(new_n842), .C2(new_n442), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n843), .B1(new_n852), .B2(KEYINPUT103), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n836), .A2(G68), .A3(new_n389), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT16), .B1(new_n854), .B2(new_n381), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n839), .B1(new_n855), .B2(new_n424), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n856), .A2(new_n391), .A3(new_n841), .ZN(new_n857));
  INV_X1    g0657(.A(new_n398), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n443), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT103), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n860), .A2(new_n861), .A3(new_n434), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n851), .B1(new_n853), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n635), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n439), .A2(new_n440), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n444), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n844), .A2(new_n851), .A3(new_n432), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT104), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n442), .B1(new_n857), .B2(new_n858), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT103), .B1(new_n870), .B2(new_n845), .ZN(new_n871));
  INV_X1    g0671(.A(new_n843), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n862), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT104), .ZN(new_n875));
  INV_X1    g0675(.A(new_n868), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n850), .B1(new_n869), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n865), .B1(new_n611), .B2(new_n416), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n422), .A2(new_n435), .A3(KEYINPUT106), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n612), .A2(new_n865), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n847), .A2(KEYINPUT106), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n881), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n880), .B1(new_n886), .B2(KEYINPUT37), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n878), .A2(new_n887), .A3(KEYINPUT39), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n850), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n875), .B1(new_n874), .B2(new_n876), .ZN(new_n891));
  AOI211_X1 g0691(.A(KEYINPUT104), .B(new_n868), .C1(new_n873), .C2(KEYINPUT37), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(KEYINPUT105), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT105), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n895), .B(new_n890), .C1(new_n891), .C2(new_n892), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n849), .B1(new_n891), .B2(new_n892), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n894), .A2(new_n896), .B1(new_n879), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT39), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n889), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n336), .A2(new_n637), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n897), .A2(new_n879), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n878), .A2(new_n895), .ZN(new_n904));
  AOI211_X1 g0704(.A(KEYINPUT105), .B(new_n850), .C1(new_n869), .C2(new_n877), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n367), .A2(new_n637), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n779), .B2(new_n792), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n335), .A2(new_n637), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n336), .A2(new_n339), .A3(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n335), .B(new_n637), .C1(new_n613), .C2(new_n321), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n908), .A2(new_n913), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n906), .A2(new_n914), .B1(new_n612), .B2(new_n635), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n902), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n616), .B1(new_n449), .B2(new_n667), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n916), .B(new_n917), .Z(new_n918));
  INV_X1    g0718(.A(G330), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n673), .A2(new_n678), .A3(new_n668), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n920), .A2(new_n679), .A3(KEYINPUT30), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n696), .A2(new_n684), .ZN(new_n922));
  OAI211_X1 g0722(.A(KEYINPUT31), .B(new_n637), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n691), .B(new_n923), .C1(new_n698), .C2(new_n689), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT107), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n637), .B1(new_n921), .B2(new_n922), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n688), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT107), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n927), .A2(new_n928), .A3(new_n691), .A4(new_n923), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n786), .A2(new_n780), .A3(new_n788), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n931), .A2(new_n789), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n913), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n930), .B(new_n933), .C1(new_n878), .C2(new_n887), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(KEYINPUT40), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT40), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n933), .A2(new_n930), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n935), .B1(new_n898), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n618), .B1(new_n929), .B2(new_n925), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n919), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n939), .B2(new_n938), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n918), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(KEYINPUT108), .ZN(new_n943));
  INV_X1    g0743(.A(G13), .ZN(new_n944));
  OAI21_X1  g0744(.A(G1), .B1(new_n944), .B2(G20), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n943), .B(new_n945), .C1(new_n918), .C2(new_n941), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n942), .A2(KEYINPUT108), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n832), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT109), .ZN(G367));
  OAI21_X1  g0749(.A(new_n725), .B1(new_n230), .B2(new_n360), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n241), .A2(new_n715), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n952), .A2(new_n707), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n741), .A2(new_n749), .B1(new_n730), .B2(new_n376), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(G68), .B2(new_n746), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n735), .A2(new_n267), .B1(new_n748), .B2(new_n811), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n345), .B(new_n956), .C1(G50), .C2(new_n808), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n738), .A2(G143), .B1(new_n763), .B2(G77), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n955), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n730), .A2(new_n542), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT46), .ZN(new_n961));
  AOI22_X1  g0761(.A1(G107), .A2(new_n746), .B1(new_n738), .B2(G311), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n274), .B1(new_n804), .B2(G303), .ZN(new_n963));
  AOI22_X1  g0763(.A1(G283), .A2(new_n808), .B1(new_n765), .B2(G317), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n740), .A2(G294), .B1(new_n763), .B2(G97), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n962), .A2(new_n963), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n959), .B1(new_n961), .B2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT47), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n721), .B1(new_n967), .B2(new_n968), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n485), .A2(new_n489), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n637), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n621), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT110), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n621), .A2(KEYINPUT110), .A3(new_n972), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n975), .B(new_n976), .C1(new_n484), .C2(new_n972), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n953), .B1(new_n969), .B2(new_n970), .C1(new_n977), .C2(new_n775), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n580), .A2(new_n637), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n623), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n619), .A2(new_n637), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n652), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT45), .Z(new_n984));
  NOR2_X1   g0784(.A1(new_n652), .A2(new_n982), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT44), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(new_n648), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n651), .A2(new_n643), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n647), .B2(new_n651), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(new_n642), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n700), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n700), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n656), .B(KEYINPUT41), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n705), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n648), .A2(new_n982), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT112), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT111), .Z(new_n1001));
  XNOR2_X1  g0801(.A(new_n999), .B(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n989), .B1(new_n980), .B2(new_n981), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1004), .A2(KEYINPUT42), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n594), .B1(new_n980), .B2(new_n534), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n1004), .A2(KEYINPUT42), .B1(new_n645), .B2(new_n1006), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n1005), .A2(new_n1007), .B1(KEYINPUT43), .B2(new_n977), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1002), .B(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n978), .B1(new_n997), .B2(new_n1009), .ZN(G387));
  OR2_X1    g0810(.A1(new_n647), .A2(new_n775), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n655), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n1012), .A2(new_n711), .B1(G107), .B2(new_n230), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1012), .A2(KEYINPUT113), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(KEYINPUT113), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n396), .A2(new_n263), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1016), .A2(KEYINPUT50), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n288), .B1(new_n207), .B2(new_n213), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n1016), .B2(KEYINPUT50), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .A4(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n715), .B1(new_n238), .B2(G45), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1013), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n708), .B1(new_n1022), .B2(new_n726), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n734), .A2(new_n207), .B1(new_n748), .B2(new_n267), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n345), .B(new_n1024), .C1(G50), .C2(new_n804), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n730), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(G77), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n465), .A2(new_n746), .B1(new_n740), .B2(new_n396), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n738), .A2(G159), .B1(new_n763), .B2(G97), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1025), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n274), .B1(new_n765), .B2(G326), .ZN(new_n1031));
  INV_X1    g0831(.A(G283), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n745), .A2(new_n1032), .B1(new_n730), .B2(new_n760), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n804), .A2(G317), .B1(new_n808), .B2(G303), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n810), .B2(new_n755), .C1(new_n754), .C2(new_n741), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT48), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1033), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n1036), .B2(new_n1035), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT49), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1031), .B1(new_n542), .B2(new_n742), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1030), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1023), .B1(new_n1042), .B2(new_n721), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n991), .A2(new_n705), .B1(new_n1011), .B2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n656), .B(KEYINPUT114), .Z(new_n1045));
  NAND2_X1  g0845(.A1(new_n992), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n700), .A2(new_n991), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(G393));
  OAI21_X1  g0848(.A(new_n725), .B1(new_n304), .B2(new_n230), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n248), .A2(new_n715), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n708), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n345), .B1(new_n765), .B2(G143), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n207), .B2(new_n730), .C1(new_n209), .C2(new_n742), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT115), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n745), .A2(new_n213), .B1(new_n734), .B2(new_n265), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G150), .A2(new_n738), .B1(new_n804), .B2(G159), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT51), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1055), .B(new_n1057), .C1(G50), .C2(new_n740), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n745), .A2(new_n542), .B1(new_n734), .B2(new_n760), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G317), .A2(new_n738), .B1(new_n804), .B2(G311), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT52), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1059), .B(new_n1061), .C1(G303), .C2(new_n740), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n345), .B1(new_n748), .B2(new_n755), .C1(new_n215), .C2(new_n742), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G283), .B2(new_n1026), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT116), .Z(new_n1065));
  AOI22_X1  g0865(.A1(new_n1054), .A2(new_n1058), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1066), .A2(KEYINPUT117), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n721), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n1066), .B2(KEYINPUT117), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1051), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n982), .B2(new_n775), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n993), .A2(new_n1045), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n988), .A2(new_n992), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1071), .B1(new_n706), .B2(new_n988), .C1(new_n1072), .C2(new_n1074), .ZN(G390));
  AOI21_X1  g0875(.A(new_n919), .B1(new_n925), .B2(new_n929), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n933), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n913), .B1(new_n794), .B2(new_n932), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n908), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n907), .B1(new_n666), .B2(new_n792), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n792), .A2(new_n699), .A3(G330), .A4(new_n912), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n912), .B1(new_n1076), .B2(new_n792), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT119), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n919), .B(new_n932), .C1(new_n925), .C2(new_n929), .ZN(new_n1086));
  OAI21_X1  g0886(.A(KEYINPUT119), .B1(new_n1086), .B2(new_n912), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1079), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1076), .A2(new_n449), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n917), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n901), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n908), .B2(new_n913), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n889), .B(new_n1093), .C1(new_n898), .C2(new_n899), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1092), .B1(new_n1080), .B2(new_n913), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n878), .A2(new_n887), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1077), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT118), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1081), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n1094), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1077), .A2(new_n1100), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1091), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1079), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n930), .A2(G330), .A3(new_n792), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1107), .A2(new_n1084), .A3(new_n913), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1082), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1106), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1090), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1094), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n888), .B1(new_n906), .B2(KEYINPUT39), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1097), .B1(new_n1116), .B2(new_n1093), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1114), .B(new_n1115), .C1(new_n1117), .C2(new_n1103), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1105), .A2(new_n1045), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1115), .B1(new_n1117), .B2(new_n1103), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1116), .A2(new_n722), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n708), .B1(new_n798), .B2(new_n396), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n745), .A2(new_n749), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n741), .A2(new_n811), .B1(new_n742), .B2(new_n263), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1123), .B(new_n1124), .C1(G128), .C2(new_n738), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n730), .A2(new_n267), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT53), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n769), .A2(G125), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT54), .B(G143), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n274), .B1(new_n734), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G132), .B2(new_n804), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1125), .A2(new_n1127), .A3(new_n1128), .A4(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n738), .A2(G283), .B1(new_n808), .B2(G97), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n215), .B2(new_n741), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT120), .Z(new_n1135));
  AOI211_X1 g0935(.A(new_n274), .B(new_n731), .C1(G116), .C2(new_n804), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n746), .A2(G77), .B1(new_n763), .B2(G68), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1136), .B(new_n1137), .C1(new_n760), .C2(new_n768), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1132), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1122), .B1(new_n1139), .B2(new_n721), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1120), .A2(new_n705), .B1(new_n1121), .B2(new_n1140), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1119), .A2(KEYINPUT121), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(KEYINPUT121), .B1(new_n1119), .B2(new_n1141), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1142), .A2(new_n1143), .ZN(G378));
  INV_X1    g0944(.A(new_n937), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n906), .A2(new_n1145), .B1(KEYINPUT40), .B2(new_n934), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n607), .A2(new_n373), .A3(new_n609), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n272), .A2(new_n864), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1147), .B(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1150), .B(new_n1151), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1146), .A2(new_n1152), .A3(new_n919), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1151), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1150), .B(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n938), .B2(G330), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n916), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1152), .B1(new_n1146), .B2(new_n919), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n938), .A2(new_n1155), .A3(G330), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1158), .A2(new_n902), .A3(new_n1159), .A4(new_n915), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT123), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1157), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n916), .B(KEYINPUT123), .C1(new_n1153), .C2(new_n1156), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n705), .A3(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n503), .A2(new_n274), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n360), .B2(new_n734), .C1(new_n207), .C2(new_n745), .ZN(new_n1166));
  OAI21_X1  g0966(.A(KEYINPUT122), .B1(new_n735), .B2(new_n215), .ZN(new_n1167));
  OR3_X1    g0967(.A1(new_n735), .A2(KEYINPUT122), .A3(new_n215), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1166), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n810), .A2(new_n542), .B1(new_n742), .B2(new_n376), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1027), .B1(new_n741), .B2(new_n304), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1169), .B(new_n1172), .C1(new_n1032), .C2(new_n768), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT58), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n263), .B1(G33), .B2(G41), .C1(new_n503), .C2(new_n274), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n738), .A2(G125), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n741), .B2(new_n817), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n804), .A2(G128), .B1(new_n808), .B2(G137), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n730), .B2(new_n1129), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1179), .B(new_n1181), .C1(G150), .C2(new_n746), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n763), .A2(G159), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G33), .B(G41), .C1(new_n765), .C2(G124), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1177), .B1(new_n1174), .B2(new_n1173), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n721), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n707), .B1(new_n797), .B2(new_n263), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(new_n1155), .C2(new_n723), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1164), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1105), .A2(new_n1113), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1162), .A2(new_n1194), .A3(new_n1163), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT57), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1045), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1196), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1198), .B1(new_n1199), .B2(new_n1194), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1193), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(G375));
  NAND2_X1  g1002(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1114), .A2(new_n1203), .A3(new_n996), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT124), .Z(new_n1205));
  OAI22_X1  g1005(.A1(new_n810), .A2(new_n760), .B1(new_n730), .B2(new_n304), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G116), .B2(new_n740), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n769), .A2(G303), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n345), .B1(new_n734), .B2(new_n215), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G283), .B2(new_n804), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n746), .A2(new_n465), .B1(new_n763), .B2(G77), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1207), .A2(new_n1208), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n810), .A2(new_n817), .B1(new_n730), .B2(new_n749), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G50), .B2(new_n746), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n769), .A2(G128), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n274), .B1(new_n734), .B2(new_n267), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G137), .B2(new_n804), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1129), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n740), .A2(new_n1218), .B1(new_n763), .B2(G58), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1214), .A2(new_n1215), .A3(new_n1217), .A4(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1068), .B1(new_n1212), .B2(new_n1220), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n707), .B(new_n1221), .C1(new_n207), .C2(new_n797), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n912), .B2(new_n723), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n1088), .B2(new_n706), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1205), .A2(new_n1225), .ZN(G381));
  NAND2_X1  g1026(.A1(new_n1119), .A2(new_n1141), .ZN(new_n1227));
  INV_X1    g1027(.A(G390), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n823), .ZN(new_n1229));
  OR4_X1    g1029(.A1(G396), .A2(new_n1229), .A3(G387), .A4(G393), .ZN(new_n1230));
  OR4_X1    g1030(.A1(new_n1227), .A2(new_n1230), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1031(.A(new_n1227), .ZN(new_n1232));
  INV_X1    g1032(.A(G213), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1233), .A2(G343), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1201), .A2(new_n1232), .A3(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(G407), .A2(G213), .A3(new_n1235), .ZN(G409));
  XNOR2_X1  g1036(.A(G387), .B(G390), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(G393), .B(new_n777), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1237), .B(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1193), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1240), .A2(G378), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n705), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1192), .B(new_n1244), .C1(new_n1195), .C2(new_n995), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1232), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1242), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1234), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1045), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT60), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1087), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1252), .A2(KEYINPUT60), .A3(new_n1106), .A4(new_n1090), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT125), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1088), .A2(KEYINPUT125), .A3(KEYINPUT60), .A4(new_n1090), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT126), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1251), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1258), .B1(new_n1251), .B2(new_n1257), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1225), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n823), .ZN(new_n1262));
  OAI211_X1 g1062(.A(G384), .B(new_n1225), .C1(new_n1259), .C2(new_n1260), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1247), .A2(new_n1248), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT62), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT62), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1247), .A2(new_n1267), .A3(new_n1248), .A4(new_n1264), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT61), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1264), .A2(KEYINPUT127), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1201), .A2(G378), .B1(new_n1232), .B2(new_n1245), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1271), .B1(new_n1272), .B2(new_n1234), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1234), .A2(G2897), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT127), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1274), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1274), .ZN(new_n1278));
  AOI211_X1 g1078(.A(KEYINPUT127), .B(new_n1278), .C1(new_n1262), .C2(new_n1263), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1270), .B1(new_n1273), .B2(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1239), .B1(new_n1269), .B2(new_n1281), .ZN(new_n1282));
  OAI221_X1 g1082(.A(new_n1271), .B1(new_n1272), .B2(new_n1234), .C1(new_n1277), .C2(new_n1279), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT63), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1239), .B1(new_n1265), .B2(new_n1284), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1247), .A2(KEYINPUT63), .A3(new_n1248), .A4(new_n1264), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1283), .A2(new_n1285), .A3(new_n1270), .A4(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1282), .A2(new_n1287), .ZN(G405));
  INV_X1    g1088(.A(new_n1242), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1201), .A2(new_n1227), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1264), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1242), .B(new_n1275), .C1(new_n1227), .C2(new_n1201), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(new_n1293), .B(new_n1239), .ZN(G402));
endmodule


