//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964;
  XOR2_X1   g000(.A(G113gat), .B(G120gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT1), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT68), .ZN(new_n204));
  XNOR2_X1  g003(.A(G127gat), .B(G134gat), .ZN(new_n205));
  OAI211_X1 g004(.A(new_n202), .B(new_n203), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G127gat), .B(G134gat), .Z(new_n207));
  NAND2_X1  g006(.A1(new_n204), .A2(new_n203), .ZN(new_n208));
  XNOR2_X1  g007(.A(G113gat), .B(G120gat), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n207), .B(new_n208), .C1(KEYINPUT1), .C2(new_n209), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT66), .ZN(new_n212));
  NOR3_X1   g011(.A1(new_n212), .A2(G169gat), .A3(G176gat), .ZN(new_n213));
  INV_X1    g012(.A(G169gat), .ZN(new_n214));
  INV_X1    g013(.A(G176gat), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT66), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT23), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n220), .B(new_n221), .C1(G183gat), .C2(G190gat), .ZN(new_n222));
  AND2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n214), .A2(new_n215), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n217), .A2(new_n222), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT25), .ZN(new_n228));
  INV_X1    g027(.A(new_n218), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT27), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G183gat), .ZN(new_n231));
  INV_X1    g030(.A(G183gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT27), .ZN(new_n233));
  INV_X1    g032(.A(G190gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n229), .B1(new_n235), .B2(KEYINPUT28), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n231), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n230), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n233), .A4(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n212), .ZN(new_n242));
  NOR2_X1   g041(.A1(G169gat), .A2(G176gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT66), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT26), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n224), .A2(KEYINPUT26), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(new_n214), .B2(new_n215), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n236), .B(new_n241), .C1(new_n245), .C2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n249), .A2(new_n221), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n251));
  OR3_X1    g050(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT64), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n218), .A2(new_n253), .A3(new_n219), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n250), .A2(new_n251), .A3(new_n252), .A4(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n224), .A2(new_n225), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n243), .A2(KEYINPUT23), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT25), .B1(G169gat), .B2(G176gat), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  AND4_X1   g059(.A1(new_n211), .A2(new_n228), .A3(new_n248), .A4(new_n260), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n227), .A2(KEYINPUT25), .B1(new_n255), .B2(new_n259), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n211), .B1(new_n262), .B2(new_n248), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G227gat), .A2(G233gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(G15gat), .B(G43gat), .Z(new_n267));
  XOR2_X1   g066(.A(G71gat), .B(G99gat), .Z(new_n268));
  XOR2_X1   g067(.A(new_n267), .B(new_n268), .Z(new_n269));
  NAND3_X1  g068(.A1(new_n228), .A2(new_n248), .A3(new_n260), .ZN(new_n270));
  INV_X1    g069(.A(new_n211), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n262), .A2(new_n211), .A3(new_n248), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n265), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT33), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(KEYINPUT32), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n269), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT69), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n279), .B(new_n269), .C1(new_n274), .C2(new_n276), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n265), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(new_n261), .B2(new_n263), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n269), .A2(KEYINPUT33), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n283), .A2(KEYINPUT32), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n266), .B1(new_n281), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n266), .ZN(new_n288));
  AOI211_X1 g087(.A(new_n288), .B(new_n285), .C1(new_n278), .C2(new_n280), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NOR3_X1   g090(.A1(new_n287), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n276), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n283), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n279), .B1(new_n294), .B2(new_n269), .ZN(new_n295));
  INV_X1    g094(.A(new_n269), .ZN(new_n296));
  AOI211_X1 g095(.A(KEYINPUT69), .B(new_n296), .C1(new_n283), .C2(new_n293), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n286), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n288), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n281), .A2(new_n266), .A3(new_n286), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n290), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(G197gat), .B(G204gat), .Z(new_n303));
  XOR2_X1   g102(.A(KEYINPUT73), .B(G211gat), .Z(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G218gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT22), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G211gat), .B(G218gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT29), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT3), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G148gat), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT76), .B1(new_n314), .B2(G141gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT76), .ZN(new_n316));
  INV_X1    g115(.A(G141gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n317), .A3(G148gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n314), .A2(G141gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n315), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT2), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT77), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(new_n327), .A3(new_n321), .ZN(new_n328));
  INV_X1    g127(.A(new_n321), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT77), .B1(new_n329), .B2(new_n325), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n324), .A2(KEYINPUT78), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT78), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n328), .A2(new_n330), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n333), .B1(new_n334), .B2(new_n323), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n317), .A2(G148gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n319), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n338), .A2(KEYINPUT75), .B1(KEYINPUT2), .B2(new_n321), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(KEYINPUT75), .B2(new_n338), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n325), .B1(new_n329), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n321), .A2(KEYINPUT74), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n336), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n313), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n336), .A2(new_n312), .A3(new_n345), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n309), .B1(new_n348), .B2(new_n310), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G22gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n332), .A2(new_n335), .B1(new_n340), .B2(new_n344), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n353), .B1(new_n311), .B2(new_n312), .ZN(new_n354));
  OAI21_X1  g153(.A(G22gat), .B1(new_n354), .B2(new_n349), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT81), .ZN(new_n357));
  OAI211_X1 g156(.A(G228gat), .B(G233gat), .C1(new_n354), .C2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n352), .A2(new_n358), .A3(new_n355), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G78gat), .B(G106gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT31), .B(G50gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(KEYINPUT82), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT82), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n360), .A2(new_n368), .A3(new_n365), .A4(new_n361), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n302), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT4), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n336), .A2(new_n372), .A3(new_n345), .A4(new_n211), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n353), .A2(KEYINPUT79), .A3(new_n372), .A4(new_n211), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n336), .A2(new_n345), .A3(new_n211), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT4), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G225gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n211), .B1(new_n353), .B2(new_n312), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n346), .A2(KEYINPUT3), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n346), .A2(new_n271), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n377), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n387), .B1(new_n389), .B2(new_n381), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n373), .A2(new_n378), .B1(new_n382), .B2(new_n383), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n386), .A2(new_n381), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT85), .ZN(new_n396));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397));
  INV_X1    g196(.A(G85gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n397), .B(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT0), .B(G57gat), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n399), .B(new_n400), .Z(new_n401));
  NAND3_X1  g200(.A1(new_n395), .A2(new_n396), .A3(new_n401), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n385), .A2(new_n390), .B1(new_n392), .B2(new_n393), .ZN(new_n403));
  INV_X1    g202(.A(new_n401), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT85), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT6), .B1(new_n403), .B2(new_n404), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT6), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n403), .A2(new_n409), .A3(new_n404), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g211(.A1(G226gat), .A2(G233gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n270), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT29), .B1(new_n262), .B2(new_n248), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n414), .B1(new_n415), .B2(new_n413), .ZN(new_n416));
  INV_X1    g215(.A(new_n309), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n414), .B(new_n309), .C1(new_n415), .C2(new_n413), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G8gat), .B(G36gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(G64gat), .B(G92gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n423), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n425), .B1(new_n418), .B2(new_n419), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT30), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n420), .A2(KEYINPUT30), .A3(new_n423), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n430), .A2(KEYINPUT35), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n371), .A2(new_n412), .A3(new_n431), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n367), .A2(new_n369), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n291), .B1(new_n287), .B2(new_n289), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n299), .A2(new_n300), .A3(new_n290), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n437), .A2(KEYINPUT88), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(KEYINPUT88), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n407), .B1(new_n404), .B2(new_n403), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n411), .ZN(new_n441));
  INV_X1    g240(.A(new_n430), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n438), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT35), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n432), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT83), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n370), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n367), .A2(new_n369), .A3(KEYINPUT83), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n443), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT37), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n451), .B1(new_n420), .B2(KEYINPUT86), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT86), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n418), .A2(new_n419), .A3(new_n453), .A4(KEYINPUT37), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n425), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT38), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n424), .B1(new_n455), .B2(new_n456), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n391), .A2(new_n404), .A3(new_n394), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n409), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n405), .B2(new_n402), .ZN(new_n462));
  NOR3_X1   g261(.A1(new_n459), .A2(new_n462), .A3(new_n410), .ZN(new_n463));
  INV_X1    g262(.A(new_n373), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n372), .B1(new_n353), .B2(new_n211), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n348), .A2(new_n271), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n353), .A2(new_n312), .ZN(new_n467));
  OAI22_X1  g266(.A1(new_n464), .A2(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT39), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n469), .A3(new_n381), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n404), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT39), .B1(new_n389), .B2(new_n381), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n472), .B1(new_n381), .B2(new_n468), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT84), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT40), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT40), .ZN(new_n476));
  OAI211_X1 g275(.A(KEYINPUT84), .B(new_n476), .C1(new_n471), .C2(new_n473), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n406), .A2(new_n475), .A3(new_n430), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n433), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT87), .B1(new_n463), .B2(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n408), .A2(new_n411), .A3(new_n457), .A4(new_n458), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT87), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n481), .A2(new_n482), .A3(new_n433), .A4(new_n478), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n450), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT36), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n434), .A2(new_n435), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT72), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT72), .A4(new_n485), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT71), .B1(new_n436), .B2(KEYINPUT36), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT71), .ZN(new_n492));
  AOI211_X1 g291(.A(new_n492), .B(new_n485), .C1(new_n434), .C2(new_n435), .ZN(new_n493));
  OAI22_X1  g292(.A1(new_n488), .A2(new_n490), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n484), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n446), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G15gat), .B(G22gat), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT16), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(G1gat), .B1(new_n497), .B2(KEYINPUT89), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n497), .A2(KEYINPUT89), .A3(G1gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G8gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT21), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(KEYINPUT92), .ZN(new_n508));
  INV_X1    g307(.A(G57gat), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n509), .A2(KEYINPUT91), .A3(G64gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(G71gat), .B(G78gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(G57gat), .B(G64gat), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT91), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n508), .A2(new_n510), .A3(new_n511), .A4(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n511), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT9), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n516), .B1(new_n517), .B2(new_n512), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n505), .B1(new_n506), .B2(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n519), .B(KEYINPUT21), .Z(new_n521));
  AOI21_X1  g320(.A(new_n520), .B1(new_n505), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n523));
  XNOR2_X1  g322(.A(G183gat), .B(G211gat), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n523), .B(new_n524), .Z(new_n525));
  XNOR2_X1  g324(.A(new_n522), .B(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(G231gat), .A2(G233gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(KEYINPUT93), .ZN(new_n528));
  XNOR2_X1  g327(.A(G127gat), .B(G155gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n526), .B(new_n530), .Z(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT14), .ZN(new_n533));
  INV_X1    g332(.A(G29gat), .ZN(new_n534));
  INV_X1    g333(.A(G36gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n536), .A2(new_n537), .B1(G29gat), .B2(G36gat), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n538), .A2(KEYINPUT15), .ZN(new_n539));
  XNOR2_X1  g338(.A(G43gat), .B(G50gat), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n538), .A2(KEYINPUT15), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n540), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n544), .A2(KEYINPUT17), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(KEYINPUT17), .ZN(new_n546));
  INV_X1    g345(.A(G99gat), .ZN(new_n547));
  INV_X1    g346(.A(G106gat), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT95), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT95), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n550), .A2(G99gat), .A3(G106gat), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n549), .A2(KEYINPUT8), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G85gat), .A2(G92gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT7), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n553), .B1(new_n554), .B2(KEYINPUT94), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT94), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n556), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n555), .B(new_n557), .C1(G85gat), .C2(G92gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(G99gat), .B(G106gat), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  OR4_X1    g359(.A1(KEYINPUT96), .A2(new_n552), .A3(new_n558), .A4(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n552), .A2(new_n558), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n559), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n560), .B1(new_n558), .B2(new_n552), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(KEYINPUT96), .A3(new_n564), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n545), .A2(new_n546), .A3(new_n561), .A4(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(G190gat), .B(G218gat), .Z(new_n567));
  INV_X1    g366(.A(KEYINPUT41), .ZN(new_n568));
  NAND2_X1  g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569));
  OAI22_X1  g368(.A1(new_n567), .A2(KEYINPUT97), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n544), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n565), .A2(new_n561), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G134gat), .B(G162gat), .Z(new_n575));
  OR2_X1    g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n575), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n567), .A2(KEYINPUT97), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n579), .B(KEYINPUT98), .Z(new_n580));
  NAND2_X1  g379(.A1(new_n569), .A2(new_n568), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n580), .B(new_n581), .Z(new_n582));
  OR2_X1    g381(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n576), .A2(new_n582), .A3(new_n577), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n532), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n545), .A2(new_n505), .A3(new_n546), .ZN(new_n588));
  OR2_X1    g387(.A1(new_n588), .A2(KEYINPUT90), .ZN(new_n589));
  NAND2_X1  g388(.A1(G229gat), .A2(G233gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n505), .A2(new_n544), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n591), .B1(new_n588), .B2(KEYINPUT90), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT18), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n505), .B(new_n544), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n590), .B(KEYINPUT13), .Z(new_n596));
  AOI22_X1  g395(.A1(new_n593), .A2(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n589), .A2(new_n592), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(KEYINPUT18), .A3(new_n590), .ZN(new_n599));
  XNOR2_X1  g398(.A(G113gat), .B(G141gat), .ZN(new_n600));
  INV_X1    g399(.A(G197gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(KEYINPUT11), .B(G169gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT12), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n597), .A2(new_n599), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n605), .B1(new_n597), .B2(new_n599), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G230gat), .A2(G233gat), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n572), .A2(new_n519), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n563), .A2(KEYINPUT99), .A3(new_n564), .ZN(new_n613));
  OR3_X1    g412(.A1(new_n562), .A2(KEYINPUT99), .A3(new_n559), .ZN(new_n614));
  INV_X1    g413(.A(new_n519), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(KEYINPUT10), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n572), .A2(KEYINPUT10), .A3(new_n615), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n611), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n612), .A2(new_n611), .A3(new_n616), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n626), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n621), .A2(new_n622), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n587), .A2(new_n609), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n496), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n441), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g437(.A1(new_n634), .A2(new_n442), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT42), .B1(new_n639), .B2(new_n504), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT100), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G8gat), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  MUX2_X1   g442(.A(KEYINPUT42), .B(new_n640), .S(new_n643), .Z(G1325gat));
  NAND2_X1  g443(.A1(new_n494), .A2(KEYINPUT102), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT36), .B1(new_n292), .B2(new_n301), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n492), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n436), .A2(KEYINPUT71), .A3(KEYINPUT36), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n486), .A2(new_n487), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n489), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n645), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n635), .A2(G15gat), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT101), .ZN(new_n657));
  INV_X1    g456(.A(G15gat), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(new_n634), .B2(new_n302), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n656), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n660), .B1(new_n657), .B2(new_n659), .ZN(G1326gat));
  NAND2_X1  g460(.A1(new_n448), .A2(new_n449), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n634), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT43), .B(G22gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1327gat));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666));
  INV_X1    g465(.A(new_n432), .ZN(new_n667));
  OR3_X1    g466(.A1(new_n438), .A2(new_n439), .A3(new_n443), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n667), .B1(new_n668), .B2(KEYINPUT35), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n650), .B1(new_n649), .B2(new_n652), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n484), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT103), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n484), .B(new_n674), .C1(new_n670), .C2(new_n671), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n669), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n666), .B1(new_n676), .B2(new_n585), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n608), .A2(new_n531), .A3(new_n630), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n585), .B1(new_n446), .B2(new_n495), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT44), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(G29gat), .B1(new_n682), .B2(new_n441), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n679), .A2(new_n678), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(new_n534), .A3(new_n636), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT45), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n686), .ZN(G1328gat));
  OAI21_X1  g486(.A(G36gat), .B1(new_n682), .B2(new_n442), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n684), .A2(new_n535), .A3(new_n430), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT46), .Z(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(G1329gat));
  NAND3_X1  g490(.A1(new_n681), .A2(G43gat), .A3(new_n655), .ZN(new_n692));
  INV_X1    g491(.A(new_n684), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(new_n302), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(G43gat), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n697));
  OR3_X1    g496(.A1(new_n693), .A2(G50gat), .A3(new_n662), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n677), .A2(new_n370), .A3(new_n678), .A4(new_n680), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT104), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(G50gat), .B1(new_n699), .B2(KEYINPUT104), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n698), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT48), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT48), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n698), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n662), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n681), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n706), .B1(new_n708), .B2(G50gat), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n697), .B1(new_n704), .B2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n680), .ZN(new_n712));
  INV_X1    g511(.A(new_n675), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n674), .B1(new_n654), .B2(new_n484), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n446), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n586), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n712), .B1(new_n716), .B2(new_n666), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n717), .A2(new_n718), .A3(new_n370), .A4(new_n678), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n719), .A2(new_n700), .A3(G50gat), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n705), .B1(new_n720), .B2(new_n698), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n721), .A2(KEYINPUT105), .A3(new_n709), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n711), .A2(new_n722), .ZN(G1331gat));
  INV_X1    g522(.A(new_n587), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n724), .A2(new_n609), .A3(new_n631), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n715), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n636), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g527(.A(new_n726), .B(KEYINPUT106), .ZN(new_n729));
  XOR2_X1   g528(.A(new_n430), .B(KEYINPUT107), .Z(new_n730));
  AOI21_X1  g529(.A(new_n730), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT108), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n729), .A2(new_n734), .A3(new_n731), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1333gat));
  NAND3_X1  g537(.A1(new_n729), .A2(G71gat), .A3(new_n655), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n726), .A2(new_n436), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(G71gat), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g541(.A1(new_n729), .A2(new_n707), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g543(.A1(new_n609), .A2(new_n531), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n715), .A2(new_n586), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n747), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n631), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(G85gat), .B1(new_n751), .B2(new_n636), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n753));
  INV_X1    g552(.A(new_n745), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n631), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n717), .A2(new_n755), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n756), .A2(new_n398), .A3(new_n441), .ZN(new_n757));
  OR3_X1    g556(.A1(new_n752), .A2(new_n753), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n753), .B1(new_n752), .B2(new_n757), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(G1336gat));
  NAND2_X1  g559(.A1(new_n749), .A2(new_n750), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n730), .A2(G92gat), .A3(new_n631), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT52), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n756), .ZN(new_n764));
  INV_X1    g563(.A(new_n730), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n764), .A2(KEYINPUT112), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G92gat), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT112), .B1(new_n764), .B2(new_n765), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n763), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(G92gat), .B1(new_n756), .B2(new_n442), .ZN(new_n770));
  INV_X1    g569(.A(new_n762), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n747), .A2(KEYINPUT110), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n746), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n746), .A2(new_n772), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n770), .B1(new_n775), .B2(KEYINPUT111), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n775), .A2(KEYINPUT111), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT52), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n769), .A2(new_n778), .ZN(G1337gat));
  NOR3_X1   g578(.A1(new_n756), .A2(new_n547), .A3(new_n654), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n751), .A2(new_n436), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n780), .B1(new_n781), .B2(new_n547), .ZN(G1338gat));
  NOR2_X1   g581(.A1(new_n433), .A2(G106gat), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n630), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n784), .B1(new_n773), .B2(new_n774), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n677), .A2(new_n707), .A3(new_n680), .A4(new_n755), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n786), .A2(G106gat), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT53), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n677), .A2(new_n370), .A3(new_n680), .A4(new_n755), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n790));
  OAI21_X1  g589(.A(G106gat), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n791), .B1(new_n790), .B2(new_n789), .ZN(new_n792));
  INV_X1    g591(.A(new_n750), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n630), .B(new_n783), .C1(new_n793), .C2(new_n748), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n788), .B1(new_n792), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n788), .B(KEYINPUT114), .C1(new_n792), .C2(new_n796), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(G1339gat));
  NOR3_X1   g600(.A1(new_n724), .A2(new_n609), .A3(new_n630), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n618), .A2(new_n611), .A3(new_n619), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n621), .A2(KEYINPUT54), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n628), .B1(new_n620), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n805), .A2(KEYINPUT55), .A3(new_n807), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(new_n629), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n598), .A2(new_n590), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n595), .A2(new_n596), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n604), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n597), .A2(new_n599), .A3(new_n605), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n812), .A2(new_n585), .A3(new_n817), .ZN(new_n818));
  OAI22_X1  g617(.A1(new_n608), .A2(new_n812), .B1(new_n631), .B2(new_n817), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n818), .B1(new_n819), .B2(new_n585), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n532), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI211_X1 g621(.A(KEYINPUT115), .B(new_n818), .C1(new_n585), .C2(new_n819), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n803), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(new_n441), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n730), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n707), .A2(new_n302), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(G113gat), .B1(new_n831), .B2(new_n608), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n438), .A2(new_n439), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n827), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(G113gat), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(new_n836), .A3(new_n609), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n832), .A2(new_n837), .ZN(G1340gat));
  OAI21_X1  g637(.A(G120gat), .B1(new_n831), .B2(new_n631), .ZN(new_n839));
  INV_X1    g638(.A(G120gat), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n835), .A2(new_n840), .A3(new_n630), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(G1341gat));
  AOI21_X1  g641(.A(G127gat), .B1(new_n835), .B2(new_n531), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n531), .A2(G127gat), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n843), .B1(new_n830), .B2(new_n844), .ZN(G1342gat));
  INV_X1    g644(.A(G134gat), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n585), .A2(new_n430), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n826), .A2(new_n846), .A3(new_n833), .A4(new_n847), .ZN(new_n848));
  XOR2_X1   g647(.A(new_n848), .B(KEYINPUT116), .Z(new_n849));
  OR2_X1    g648(.A1(new_n849), .A2(KEYINPUT56), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(KEYINPUT56), .ZN(new_n851));
  OAI21_X1  g650(.A(G134gat), .B1(new_n831), .B2(new_n585), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(G1343gat));
  NAND2_X1  g652(.A1(new_n824), .A2(new_n370), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT117), .B1(new_n855), .B2(KEYINPUT57), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n854), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n820), .A2(new_n531), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n707), .B1(new_n860), .B2(new_n802), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(new_n858), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n856), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n655), .A2(new_n441), .A3(new_n765), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n609), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(G141gat), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n655), .A2(new_n441), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n855), .A2(KEYINPUT119), .A3(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n869));
  INV_X1    g668(.A(new_n867), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n854), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n765), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n608), .A2(G141gat), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT58), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n866), .A2(new_n874), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n855), .A2(new_n864), .A3(new_n873), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n863), .A2(new_n877), .A3(new_n864), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n877), .B1(new_n863), .B2(new_n864), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n609), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n876), .B1(new_n881), .B2(G141gat), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT58), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n875), .B1(new_n882), .B2(new_n883), .ZN(G1344gat));
  NAND3_X1  g683(.A1(new_n872), .A2(new_n314), .A3(new_n630), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(G148gat), .ZN(new_n887));
  INV_X1    g686(.A(new_n880), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n878), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n887), .B1(new_n889), .B2(new_n630), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n824), .A2(KEYINPUT57), .A3(new_n370), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n861), .A2(new_n858), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n631), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n864), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n886), .B1(new_n895), .B2(G148gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n885), .B1(new_n890), .B2(new_n896), .ZN(G1345gat));
  AOI21_X1  g696(.A(G155gat), .B1(new_n872), .B2(new_n531), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n531), .A2(G155gat), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n889), .B2(new_n899), .ZN(G1346gat));
  NAND2_X1  g699(.A1(new_n868), .A2(new_n871), .ZN(new_n901));
  INV_X1    g700(.A(G162gat), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(new_n902), .A3(new_n847), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n585), .B1(new_n888), .B2(new_n878), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(new_n902), .ZN(G1347gat));
  NOR4_X1   g704(.A1(new_n825), .A2(new_n636), .A3(new_n834), .A4(new_n730), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n214), .A3(new_n609), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n824), .A2(new_n441), .A3(new_n430), .A4(new_n828), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n908), .B(KEYINPUT120), .Z(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(G169gat), .B1(new_n910), .B2(new_n608), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n911), .A2(KEYINPUT121), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n911), .A2(KEYINPUT121), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n907), .B1(new_n912), .B2(new_n913), .ZN(G1348gat));
  AOI21_X1  g713(.A(G176gat), .B1(new_n906), .B2(new_n630), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n631), .A2(new_n215), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n909), .B2(new_n916), .ZN(G1349gat));
  OAI21_X1  g716(.A(G183gat), .B1(new_n910), .B2(new_n532), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n906), .A2(new_n231), .A3(new_n233), .A4(new_n531), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n234), .A3(new_n586), .ZN(new_n922));
  OAI21_X1  g721(.A(G190gat), .B1(new_n910), .B2(new_n585), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n923), .A2(KEYINPUT61), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n923), .A2(KEYINPUT61), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(G1351gat));
  NOR4_X1   g725(.A1(new_n854), .A2(new_n636), .A3(new_n655), .A4(new_n730), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n601), .A3(new_n609), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n654), .A2(new_n441), .A3(new_n430), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n929), .A2(KEYINPUT122), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n929), .A2(KEYINPUT122), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n932));
  OR3_X1    g731(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n930), .B2(new_n931), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n893), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n935), .A2(new_n609), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n928), .B1(new_n936), .B2(new_n601), .ZN(G1352gat));
  INV_X1    g736(.A(G204gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n927), .A2(new_n938), .A3(new_n630), .ZN(new_n939));
  XOR2_X1   g738(.A(new_n939), .B(KEYINPUT62), .Z(new_n940));
  AOI211_X1 g739(.A(new_n631), .B(new_n893), .C1(new_n933), .C2(new_n934), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(new_n938), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT124), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n940), .B(KEYINPUT124), .C1(new_n938), .C2(new_n941), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1353gat));
  NOR2_X1   g745(.A1(new_n532), .A2(new_n304), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n927), .A2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(G211gat), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n532), .B1(new_n891), .B2(new_n892), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n950), .B1(new_n930), .B2(new_n931), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n949), .B1(new_n951), .B2(KEYINPUT125), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT125), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n950), .B(new_n953), .C1(new_n931), .C2(new_n930), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n952), .A2(KEYINPUT63), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT63), .B1(new_n952), .B2(new_n954), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n948), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI211_X1 g758(.A(KEYINPUT126), .B(new_n948), .C1(new_n955), .C2(new_n956), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1354gat));
  AOI21_X1  g760(.A(G218gat), .B1(new_n927), .B2(new_n586), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n586), .A2(G218gat), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT127), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n962), .B1(new_n935), .B2(new_n964), .ZN(G1355gat));
endmodule


