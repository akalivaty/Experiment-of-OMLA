

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U557 ( .A1(n727), .A2(n726), .ZN(n728) );
  BUF_X1 U558 ( .A(n621), .Z(n622) );
  BUF_X1 U559 ( .A(n617), .Z(n618) );
  INV_X1 U560 ( .A(KEYINPUT104), .ZN(n714) );
  XOR2_X1 U561 ( .A(n717), .B(KEYINPUT27), .Z(n524) );
  XNOR2_X1 U562 ( .A(n719), .B(KEYINPUT100), .ZN(n723) );
  AND2_X1 U563 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U564 ( .A1(n773), .A2(n772), .ZN(n748) );
  INV_X1 U565 ( .A(KEYINPUT17), .ZN(n525) );
  NOR2_X1 U566 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U567 ( .A(n525), .B(KEYINPUT66), .ZN(n526) );
  NOR2_X1 U568 ( .A1(G651), .A2(n646), .ZN(n658) );
  NOR2_X1 U569 ( .A1(n537), .A2(n536), .ZN(G164) );
  NOR2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  XNOR2_X2 U571 ( .A(n527), .B(n526), .ZN(n898) );
  NAND2_X1 U572 ( .A1(G138), .A2(n898), .ZN(n529) );
  INV_X1 U573 ( .A(G2105), .ZN(n530) );
  XOR2_X1 U574 ( .A(G2104), .B(KEYINPUT65), .Z(n531) );
  AND2_X1 U575 ( .A1(n530), .A2(n531), .ZN(n617) );
  NAND2_X1 U576 ( .A1(n617), .A2(G102), .ZN(n528) );
  NAND2_X1 U577 ( .A1(n529), .A2(n528), .ZN(n537) );
  INV_X1 U578 ( .A(KEYINPUT91), .ZN(n535) );
  AND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n901) );
  NAND2_X1 U580 ( .A1(G114), .A2(n901), .ZN(n533) );
  NOR2_X1 U581 ( .A1(n531), .A2(n530), .ZN(n621) );
  NAND2_X1 U582 ( .A1(G126), .A2(n621), .ZN(n532) );
  NAND2_X1 U583 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U584 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U585 ( .A(G543), .B(KEYINPUT0), .Z(n646) );
  XNOR2_X1 U586 ( .A(G651), .B(KEYINPUT67), .ZN(n541) );
  NOR2_X1 U587 ( .A1(n646), .A2(n541), .ZN(n663) );
  NAND2_X1 U588 ( .A1(n663), .A2(G75), .ZN(n540) );
  NOR2_X1 U589 ( .A1(G543), .A2(G651), .ZN(n538) );
  XNOR2_X1 U590 ( .A(n538), .B(KEYINPUT64), .ZN(n662) );
  NAND2_X1 U591 ( .A1(G88), .A2(n662), .ZN(n539) );
  NAND2_X1 U592 ( .A1(n540), .A2(n539), .ZN(n547) );
  NOR2_X1 U593 ( .A1(n541), .A2(G543), .ZN(n542) );
  XOR2_X2 U594 ( .A(KEYINPUT1), .B(n542), .Z(n657) );
  NAND2_X1 U595 ( .A1(G62), .A2(n657), .ZN(n544) );
  NAND2_X1 U596 ( .A1(G50), .A2(n658), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U598 ( .A(KEYINPUT85), .B(n545), .Z(n546) );
  NOR2_X1 U599 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U600 ( .A(KEYINPUT86), .B(n548), .ZN(G166) );
  INV_X1 U601 ( .A(G166), .ZN(G303) );
  NAND2_X1 U602 ( .A1(n663), .A2(G78), .ZN(n550) );
  NAND2_X1 U603 ( .A1(G91), .A2(n662), .ZN(n549) );
  NAND2_X1 U604 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U605 ( .A1(G65), .A2(n657), .ZN(n552) );
  NAND2_X1 U606 ( .A1(G53), .A2(n658), .ZN(n551) );
  NAND2_X1 U607 ( .A1(n552), .A2(n551), .ZN(n553) );
  OR2_X1 U608 ( .A1(n554), .A2(n553), .ZN(G299) );
  NAND2_X1 U609 ( .A1(n657), .A2(G64), .ZN(n555) );
  XOR2_X1 U610 ( .A(KEYINPUT69), .B(n555), .Z(n557) );
  NAND2_X1 U611 ( .A1(n658), .A2(G52), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U613 ( .A(KEYINPUT70), .B(n558), .ZN(n564) );
  NAND2_X1 U614 ( .A1(n663), .A2(G77), .ZN(n560) );
  NAND2_X1 U615 ( .A1(G90), .A2(n662), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U617 ( .A(KEYINPUT9), .B(n561), .ZN(n562) );
  XNOR2_X1 U618 ( .A(KEYINPUT71), .B(n562), .ZN(n563) );
  NOR2_X1 U619 ( .A1(n564), .A2(n563), .ZN(G171) );
  AND2_X1 U620 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U621 ( .A1(G113), .A2(n901), .ZN(n566) );
  NAND2_X1 U622 ( .A1(G137), .A2(n898), .ZN(n565) );
  NAND2_X1 U623 ( .A1(n566), .A2(n565), .ZN(n571) );
  NAND2_X1 U624 ( .A1(n617), .A2(G101), .ZN(n567) );
  XOR2_X1 U625 ( .A(KEYINPUT23), .B(n567), .Z(n569) );
  NAND2_X1 U626 ( .A1(n621), .A2(G125), .ZN(n568) );
  NAND2_X1 U627 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U628 ( .A1(n571), .A2(n570), .ZN(n695) );
  BUF_X1 U629 ( .A(n695), .Z(G160) );
  INV_X1 U630 ( .A(G132), .ZN(G219) );
  INV_X1 U631 ( .A(G82), .ZN(G220) );
  INV_X1 U632 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U633 ( .A(KEYINPUT6), .B(KEYINPUT76), .ZN(n575) );
  NAND2_X1 U634 ( .A1(G63), .A2(n657), .ZN(n573) );
  NAND2_X1 U635 ( .A1(G51), .A2(n658), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U637 ( .A(n575), .B(n574), .ZN(n582) );
  NAND2_X1 U638 ( .A1(n663), .A2(G76), .ZN(n576) );
  XNOR2_X1 U639 ( .A(KEYINPUT75), .B(n576), .ZN(n579) );
  NAND2_X1 U640 ( .A1(G89), .A2(n662), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT4), .B(n577), .Z(n578) );
  NOR2_X1 U642 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U643 ( .A(n580), .B(KEYINPUT5), .ZN(n581) );
  NOR2_X1 U644 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U645 ( .A(n583), .B(KEYINPUT7), .ZN(n584) );
  XNOR2_X1 U646 ( .A(n584), .B(KEYINPUT77), .ZN(G168) );
  XOR2_X1 U647 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U648 ( .A1(G7), .A2(G661), .ZN(n585) );
  XNOR2_X1 U649 ( .A(n585), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U650 ( .A(G223), .ZN(n853) );
  NAND2_X1 U651 ( .A1(n853), .A2(G567), .ZN(n586) );
  XOR2_X1 U652 ( .A(KEYINPUT11), .B(n586), .Z(G234) );
  NAND2_X1 U653 ( .A1(n657), .A2(G56), .ZN(n587) );
  XOR2_X1 U654 ( .A(KEYINPUT14), .B(n587), .Z(n593) );
  NAND2_X1 U655 ( .A1(G81), .A2(n662), .ZN(n588) );
  XNOR2_X1 U656 ( .A(n588), .B(KEYINPUT12), .ZN(n590) );
  NAND2_X1 U657 ( .A1(G68), .A2(n663), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U659 ( .A(KEYINPUT13), .B(n591), .Z(n592) );
  XNOR2_X1 U660 ( .A(KEYINPUT72), .B(n594), .ZN(n596) );
  NAND2_X1 U661 ( .A1(G43), .A2(n658), .ZN(n595) );
  NAND2_X1 U662 ( .A1(n596), .A2(n595), .ZN(n614) );
  INV_X2 U663 ( .A(n614), .ZN(n1006) );
  NAND2_X1 U664 ( .A1(n1006), .A2(G860), .ZN(G153) );
  NAND2_X1 U665 ( .A1(G171), .A2(G868), .ZN(n606) );
  NAND2_X1 U666 ( .A1(G54), .A2(n658), .ZN(n598) );
  NAND2_X1 U667 ( .A1(G79), .A2(n663), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n603) );
  NAND2_X1 U669 ( .A1(G66), .A2(n657), .ZN(n600) );
  NAND2_X1 U670 ( .A1(G92), .A2(n662), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U672 ( .A(KEYINPUT73), .B(n601), .Z(n602) );
  NOR2_X1 U673 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U674 ( .A(KEYINPUT15), .B(n604), .Z(n989) );
  INV_X1 U675 ( .A(G868), .ZN(n676) );
  NAND2_X1 U676 ( .A1(n989), .A2(n676), .ZN(n605) );
  NAND2_X1 U677 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U678 ( .A(KEYINPUT74), .B(n607), .Z(G284) );
  NOR2_X1 U679 ( .A1(G868), .A2(G299), .ZN(n608) );
  XNOR2_X1 U680 ( .A(n608), .B(KEYINPUT78), .ZN(n610) );
  NOR2_X1 U681 ( .A1(n676), .A2(G286), .ZN(n609) );
  NOR2_X1 U682 ( .A1(n610), .A2(n609), .ZN(G297) );
  INV_X1 U683 ( .A(G860), .ZN(n633) );
  NAND2_X1 U684 ( .A1(n633), .A2(G559), .ZN(n611) );
  NAND2_X1 U685 ( .A1(n611), .A2(n989), .ZN(n612) );
  XNOR2_X1 U686 ( .A(n612), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U687 ( .A1(n989), .A2(G868), .ZN(n613) );
  NOR2_X1 U688 ( .A1(G559), .A2(n613), .ZN(n616) );
  NOR2_X1 U689 ( .A1(G868), .A2(n614), .ZN(n615) );
  NOR2_X1 U690 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U691 ( .A1(G111), .A2(n901), .ZN(n620) );
  NAND2_X1 U692 ( .A1(G99), .A2(n618), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n628) );
  NAND2_X1 U694 ( .A1(n622), .A2(G123), .ZN(n623) );
  XNOR2_X1 U695 ( .A(n623), .B(KEYINPUT18), .ZN(n625) );
  NAND2_X1 U696 ( .A1(G135), .A2(n898), .ZN(n624) );
  NAND2_X1 U697 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U698 ( .A(KEYINPUT79), .B(n626), .Z(n627) );
  NOR2_X1 U699 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U700 ( .A(KEYINPUT80), .B(n629), .ZN(n980) );
  XOR2_X1 U701 ( .A(G2096), .B(n980), .Z(n630) );
  NOR2_X1 U702 ( .A1(G2100), .A2(n630), .ZN(n631) );
  XNOR2_X1 U703 ( .A(KEYINPUT81), .B(n631), .ZN(G156) );
  NAND2_X1 U704 ( .A1(G559), .A2(n989), .ZN(n632) );
  XNOR2_X1 U705 ( .A(n632), .B(n1006), .ZN(n674) );
  NAND2_X1 U706 ( .A1(n633), .A2(n674), .ZN(n641) );
  NAND2_X1 U707 ( .A1(G67), .A2(n657), .ZN(n635) );
  NAND2_X1 U708 ( .A1(G80), .A2(n663), .ZN(n634) );
  NAND2_X1 U709 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U710 ( .A1(n662), .A2(G93), .ZN(n636) );
  XOR2_X1 U711 ( .A(KEYINPUT82), .B(n636), .Z(n637) );
  NOR2_X1 U712 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n658), .A2(G55), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n640), .A2(n639), .ZN(n677) );
  XNOR2_X1 U715 ( .A(n641), .B(n677), .ZN(G145) );
  NAND2_X1 U716 ( .A1(G49), .A2(n658), .ZN(n643) );
  NAND2_X1 U717 ( .A1(G74), .A2(G651), .ZN(n642) );
  NAND2_X1 U718 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U719 ( .A(KEYINPUT83), .B(n644), .Z(n645) );
  NOR2_X1 U720 ( .A1(n657), .A2(n645), .ZN(n648) );
  NAND2_X1 U721 ( .A1(n646), .A2(G87), .ZN(n647) );
  NAND2_X1 U722 ( .A1(n648), .A2(n647), .ZN(G288) );
  NAND2_X1 U723 ( .A1(G48), .A2(n658), .ZN(n649) );
  XNOR2_X1 U724 ( .A(n649), .B(KEYINPUT84), .ZN(n656) );
  NAND2_X1 U725 ( .A1(G61), .A2(n657), .ZN(n651) );
  NAND2_X1 U726 ( .A1(G86), .A2(n662), .ZN(n650) );
  NAND2_X1 U727 ( .A1(n651), .A2(n650), .ZN(n654) );
  NAND2_X1 U728 ( .A1(n663), .A2(G73), .ZN(n652) );
  XOR2_X1 U729 ( .A(KEYINPUT2), .B(n652), .Z(n653) );
  NOR2_X1 U730 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U731 ( .A1(n656), .A2(n655), .ZN(G305) );
  NAND2_X1 U732 ( .A1(G60), .A2(n657), .ZN(n660) );
  NAND2_X1 U733 ( .A1(G47), .A2(n658), .ZN(n659) );
  NAND2_X1 U734 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U735 ( .A(KEYINPUT68), .B(n661), .Z(n667) );
  NAND2_X1 U736 ( .A1(n662), .A2(G85), .ZN(n665) );
  NAND2_X1 U737 ( .A1(n663), .A2(G72), .ZN(n664) );
  AND2_X1 U738 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U739 ( .A1(n667), .A2(n666), .ZN(G290) );
  XNOR2_X1 U740 ( .A(KEYINPUT87), .B(G288), .ZN(n668) );
  XNOR2_X1 U741 ( .A(n668), .B(G299), .ZN(n671) );
  XNOR2_X1 U742 ( .A(G303), .B(G305), .ZN(n669) );
  XNOR2_X1 U743 ( .A(n669), .B(n677), .ZN(n670) );
  XNOR2_X1 U744 ( .A(n671), .B(n670), .ZN(n673) );
  XNOR2_X1 U745 ( .A(G290), .B(KEYINPUT19), .ZN(n672) );
  XNOR2_X1 U746 ( .A(n673), .B(n672), .ZN(n917) );
  XOR2_X1 U747 ( .A(n917), .B(n674), .Z(n675) );
  NOR2_X1 U748 ( .A1(n676), .A2(n675), .ZN(n679) );
  NOR2_X1 U749 ( .A1(G868), .A2(n677), .ZN(n678) );
  NOR2_X1 U750 ( .A1(n679), .A2(n678), .ZN(G295) );
  NAND2_X1 U751 ( .A1(G2084), .A2(G2078), .ZN(n680) );
  XOR2_X1 U752 ( .A(KEYINPUT20), .B(n680), .Z(n681) );
  NAND2_X1 U753 ( .A1(n681), .A2(G2090), .ZN(n682) );
  XNOR2_X1 U754 ( .A(n682), .B(KEYINPUT88), .ZN(n683) );
  XNOR2_X1 U755 ( .A(KEYINPUT21), .B(n683), .ZN(n684) );
  NAND2_X1 U756 ( .A1(n684), .A2(G2072), .ZN(n685) );
  XOR2_X1 U757 ( .A(KEYINPUT89), .B(n685), .Z(G158) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U759 ( .A1(G120), .A2(G69), .ZN(n686) );
  NOR2_X1 U760 ( .A1(G237), .A2(n686), .ZN(n687) );
  XNOR2_X1 U761 ( .A(KEYINPUT90), .B(n687), .ZN(n688) );
  NAND2_X1 U762 ( .A1(n688), .A2(G108), .ZN(n857) );
  NAND2_X1 U763 ( .A1(n857), .A2(G567), .ZN(n693) );
  NOR2_X1 U764 ( .A1(G220), .A2(G219), .ZN(n689) );
  XOR2_X1 U765 ( .A(KEYINPUT22), .B(n689), .Z(n690) );
  NOR2_X1 U766 ( .A1(G218), .A2(n690), .ZN(n691) );
  NAND2_X1 U767 ( .A1(G96), .A2(n691), .ZN(n858) );
  NAND2_X1 U768 ( .A1(n858), .A2(G2106), .ZN(n692) );
  NAND2_X1 U769 ( .A1(n693), .A2(n692), .ZN(n859) );
  NAND2_X1 U770 ( .A1(G483), .A2(G661), .ZN(n694) );
  NOR2_X1 U771 ( .A1(n859), .A2(n694), .ZN(n856) );
  NAND2_X1 U772 ( .A1(n856), .A2(G36), .ZN(G176) );
  AND2_X1 U773 ( .A1(n695), .A2(G40), .ZN(n773) );
  NOR2_X1 U774 ( .A1(G164), .A2(G1384), .ZN(n772) );
  INV_X1 U775 ( .A(n748), .ZN(n696) );
  NAND2_X1 U776 ( .A1(G1996), .A2(n696), .ZN(n697) );
  XNOR2_X1 U777 ( .A(n697), .B(KEYINPUT26), .ZN(n698) );
  NAND2_X1 U778 ( .A1(n748), .A2(G1341), .ZN(n701) );
  NAND2_X1 U779 ( .A1(n698), .A2(n701), .ZN(n699) );
  NAND2_X1 U780 ( .A1(n699), .A2(KEYINPUT102), .ZN(n700) );
  NAND2_X1 U781 ( .A1(n700), .A2(n1006), .ZN(n705) );
  INV_X1 U782 ( .A(KEYINPUT26), .ZN(n702) );
  NOR2_X1 U783 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U784 ( .A1(KEYINPUT102), .A2(n703), .ZN(n704) );
  NOR2_X2 U785 ( .A1(n705), .A2(n704), .ZN(n707) );
  NOR2_X1 U786 ( .A1(n707), .A2(n989), .ZN(n706) );
  XNOR2_X1 U787 ( .A(n706), .B(KEYINPUT103), .ZN(n713) );
  NAND2_X1 U788 ( .A1(n707), .A2(n989), .ZN(n711) );
  XOR2_X1 U789 ( .A(n696), .B(KEYINPUT98), .Z(n716) );
  INV_X1 U790 ( .A(n716), .ZN(n730) );
  NAND2_X1 U791 ( .A1(G2067), .A2(n730), .ZN(n709) );
  NAND2_X1 U792 ( .A1(G1348), .A2(n748), .ZN(n708) );
  NAND2_X1 U793 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U794 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U795 ( .A1(n713), .A2(n712), .ZN(n715) );
  XNOR2_X1 U796 ( .A(n715), .B(n714), .ZN(n721) );
  NAND2_X1 U797 ( .A1(G1956), .A2(n716), .ZN(n718) );
  NAND2_X1 U798 ( .A1(G2072), .A2(n730), .ZN(n717) );
  NAND2_X1 U799 ( .A1(n718), .A2(n524), .ZN(n719) );
  NOR2_X1 U800 ( .A1(n723), .A2(G299), .ZN(n720) );
  NOR2_X1 U801 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U802 ( .A(KEYINPUT105), .B(n722), .Z(n727) );
  NAND2_X1 U803 ( .A1(G299), .A2(n723), .ZN(n724) );
  XNOR2_X1 U804 ( .A(n724), .B(KEYINPUT28), .ZN(n725) );
  XNOR2_X1 U805 ( .A(KEYINPUT101), .B(n725), .ZN(n726) );
  XNOR2_X1 U806 ( .A(n728), .B(KEYINPUT29), .ZN(n734) );
  XOR2_X1 U807 ( .A(G2078), .B(KEYINPUT99), .Z(n729) );
  XNOR2_X1 U808 ( .A(KEYINPUT25), .B(n729), .ZN(n937) );
  NAND2_X1 U809 ( .A1(n730), .A2(n937), .ZN(n732) );
  INV_X1 U810 ( .A(G1961), .ZN(n1014) );
  NAND2_X1 U811 ( .A1(n1014), .A2(n748), .ZN(n731) );
  NAND2_X1 U812 ( .A1(n732), .A2(n731), .ZN(n740) );
  NAND2_X1 U813 ( .A1(G171), .A2(n740), .ZN(n733) );
  NAND2_X1 U814 ( .A1(n734), .A2(n733), .ZN(n746) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n748), .ZN(n761) );
  NAND2_X1 U816 ( .A1(n748), .A2(G8), .ZN(n735) );
  XNOR2_X1 U817 ( .A(n735), .B(KEYINPUT95), .ZN(n827) );
  INV_X1 U818 ( .A(n827), .ZN(n821) );
  NOR2_X1 U819 ( .A1(G1966), .A2(n821), .ZN(n757) );
  NOR2_X1 U820 ( .A1(n761), .A2(n757), .ZN(n736) );
  NAND2_X1 U821 ( .A1(G8), .A2(n736), .ZN(n737) );
  XNOR2_X1 U822 ( .A(KEYINPUT106), .B(n737), .ZN(n738) );
  XNOR2_X1 U823 ( .A(KEYINPUT30), .B(n738), .ZN(n739) );
  NOR2_X1 U824 ( .A1(G168), .A2(n739), .ZN(n742) );
  NOR2_X1 U825 ( .A1(G171), .A2(n740), .ZN(n741) );
  NOR2_X1 U826 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U827 ( .A(KEYINPUT31), .B(n743), .ZN(n744) );
  XNOR2_X1 U828 ( .A(n744), .B(KEYINPUT107), .ZN(n745) );
  NAND2_X1 U829 ( .A1(n746), .A2(n745), .ZN(n759) );
  AND2_X1 U830 ( .A1(G286), .A2(G8), .ZN(n747) );
  NAND2_X1 U831 ( .A1(n759), .A2(n747), .ZN(n755) );
  INV_X1 U832 ( .A(G8), .ZN(n753) );
  NOR2_X1 U833 ( .A1(G1971), .A2(n821), .ZN(n750) );
  NOR2_X1 U834 ( .A1(G2090), .A2(n748), .ZN(n749) );
  NOR2_X1 U835 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U836 ( .A1(G303), .A2(n751), .ZN(n752) );
  OR2_X1 U837 ( .A1(n753), .A2(n752), .ZN(n754) );
  AND2_X1 U838 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U839 ( .A(n756), .B(KEYINPUT32), .ZN(n765) );
  INV_X1 U840 ( .A(n757), .ZN(n758) );
  XNOR2_X1 U841 ( .A(n760), .B(KEYINPUT108), .ZN(n763) );
  NAND2_X1 U842 ( .A1(n761), .A2(G8), .ZN(n762) );
  NAND2_X1 U843 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U844 ( .A1(n765), .A2(n764), .ZN(n819) );
  NOR2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n769) );
  NOR2_X1 U846 ( .A1(G303), .A2(G1971), .ZN(n766) );
  NOR2_X1 U847 ( .A1(n769), .A2(n766), .ZN(n1000) );
  NAND2_X1 U848 ( .A1(n819), .A2(n1000), .ZN(n767) );
  NAND2_X1 U849 ( .A1(G1976), .A2(G288), .ZN(n999) );
  NAND2_X1 U850 ( .A1(n767), .A2(n999), .ZN(n768) );
  XNOR2_X1 U851 ( .A(n768), .B(KEYINPUT109), .ZN(n808) );
  INV_X1 U852 ( .A(KEYINPUT33), .ZN(n811) );
  NAND2_X1 U853 ( .A1(n827), .A2(n769), .ZN(n770) );
  NOR2_X1 U854 ( .A1(n811), .A2(n770), .ZN(n771) );
  XOR2_X1 U855 ( .A(n771), .B(KEYINPUT110), .Z(n810) );
  AND2_X1 U856 ( .A1(n827), .A2(n810), .ZN(n806) );
  XNOR2_X1 U857 ( .A(G1981), .B(G305), .ZN(n997) );
  XNOR2_X1 U858 ( .A(G1986), .B(G290), .ZN(n995) );
  INV_X1 U859 ( .A(n773), .ZN(n774) );
  NOR2_X1 U860 ( .A1(n772), .A2(n774), .ZN(n839) );
  AND2_X1 U861 ( .A1(n995), .A2(n839), .ZN(n805) );
  XNOR2_X1 U862 ( .A(KEYINPUT34), .B(KEYINPUT92), .ZN(n778) );
  NAND2_X1 U863 ( .A1(G104), .A2(n618), .ZN(n776) );
  NAND2_X1 U864 ( .A1(G140), .A2(n898), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U866 ( .A(n778), .B(n777), .ZN(n783) );
  NAND2_X1 U867 ( .A1(G116), .A2(n901), .ZN(n780) );
  NAND2_X1 U868 ( .A1(G128), .A2(n622), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U870 ( .A(KEYINPUT35), .B(n781), .Z(n782) );
  NOR2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U872 ( .A(KEYINPUT36), .B(n784), .ZN(n908) );
  XNOR2_X1 U873 ( .A(KEYINPUT37), .B(G2067), .ZN(n829) );
  NOR2_X1 U874 ( .A1(n908), .A2(n829), .ZN(n962) );
  NAND2_X1 U875 ( .A1(n839), .A2(n962), .ZN(n837) );
  NAND2_X1 U876 ( .A1(G107), .A2(n901), .ZN(n786) );
  NAND2_X1 U877 ( .A1(G95), .A2(n618), .ZN(n785) );
  NAND2_X1 U878 ( .A1(n786), .A2(n785), .ZN(n790) );
  NAND2_X1 U879 ( .A1(G119), .A2(n622), .ZN(n788) );
  NAND2_X1 U880 ( .A1(G131), .A2(n898), .ZN(n787) );
  NAND2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U883 ( .A(KEYINPUT93), .B(n791), .ZN(n893) );
  AND2_X1 U884 ( .A1(n893), .A2(G1991), .ZN(n801) );
  NAND2_X1 U885 ( .A1(G105), .A2(n618), .ZN(n792) );
  XNOR2_X1 U886 ( .A(n792), .B(KEYINPUT38), .ZN(n799) );
  NAND2_X1 U887 ( .A1(G117), .A2(n901), .ZN(n794) );
  NAND2_X1 U888 ( .A1(G141), .A2(n898), .ZN(n793) );
  NAND2_X1 U889 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U890 ( .A1(n622), .A2(G129), .ZN(n795) );
  XOR2_X1 U891 ( .A(KEYINPUT94), .B(n795), .Z(n796) );
  NOR2_X1 U892 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n895) );
  AND2_X1 U894 ( .A1(n895), .A2(G1996), .ZN(n800) );
  NOR2_X1 U895 ( .A1(n801), .A2(n800), .ZN(n969) );
  INV_X1 U896 ( .A(n839), .ZN(n802) );
  NOR2_X1 U897 ( .A1(n969), .A2(n802), .ZN(n832) );
  INV_X1 U898 ( .A(n832), .ZN(n803) );
  NAND2_X1 U899 ( .A1(n837), .A2(n803), .ZN(n804) );
  OR2_X1 U900 ( .A1(n805), .A2(n804), .ZN(n845) );
  NOR2_X1 U901 ( .A1(n997), .A2(n845), .ZN(n809) );
  AND2_X1 U902 ( .A1(n806), .A2(n809), .ZN(n807) );
  AND2_X1 U903 ( .A1(n808), .A2(n807), .ZN(n816) );
  INV_X1 U904 ( .A(n809), .ZN(n814) );
  INV_X1 U905 ( .A(n810), .ZN(n812) );
  OR2_X1 U906 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U908 ( .A1(n816), .A2(n815), .ZN(n851) );
  NOR2_X1 U909 ( .A1(G2090), .A2(G303), .ZN(n817) );
  NAND2_X1 U910 ( .A1(G8), .A2(n817), .ZN(n818) );
  NAND2_X1 U911 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U912 ( .A1(n821), .A2(n820), .ZN(n823) );
  INV_X1 U913 ( .A(KEYINPUT111), .ZN(n822) );
  XNOR2_X1 U914 ( .A(n823), .B(n822), .ZN(n843) );
  XNOR2_X1 U915 ( .A(KEYINPUT24), .B(KEYINPUT97), .ZN(n826) );
  NOR2_X1 U916 ( .A1(G1981), .A2(G305), .ZN(n824) );
  XOR2_X1 U917 ( .A(n824), .B(KEYINPUT96), .Z(n825) );
  XNOR2_X1 U918 ( .A(n826), .B(n825), .ZN(n828) );
  NAND2_X1 U919 ( .A1(n828), .A2(n827), .ZN(n841) );
  NAND2_X1 U920 ( .A1(n908), .A2(n829), .ZN(n961) );
  XOR2_X1 U921 ( .A(KEYINPUT112), .B(KEYINPUT39), .Z(n835) );
  NOR2_X1 U922 ( .A1(G1996), .A2(n895), .ZN(n972) );
  NOR2_X1 U923 ( .A1(G1991), .A2(n893), .ZN(n979) );
  NOR2_X1 U924 ( .A1(G1986), .A2(G290), .ZN(n830) );
  NOR2_X1 U925 ( .A1(n979), .A2(n830), .ZN(n831) );
  NOR2_X1 U926 ( .A1(n832), .A2(n831), .ZN(n833) );
  NOR2_X1 U927 ( .A1(n972), .A2(n833), .ZN(n834) );
  XOR2_X1 U928 ( .A(n835), .B(n834), .Z(n836) );
  NAND2_X1 U929 ( .A1(n837), .A2(n836), .ZN(n838) );
  NAND2_X1 U930 ( .A1(n961), .A2(n838), .ZN(n840) );
  NAND2_X1 U931 ( .A1(n840), .A2(n839), .ZN(n844) );
  AND2_X1 U932 ( .A1(n841), .A2(n844), .ZN(n842) );
  NAND2_X1 U933 ( .A1(n843), .A2(n842), .ZN(n849) );
  INV_X1 U934 ( .A(n844), .ZN(n847) );
  INV_X1 U935 ( .A(n845), .ZN(n846) );
  OR2_X1 U936 ( .A1(n847), .A2(n846), .ZN(n848) );
  NAND2_X1 U937 ( .A1(n849), .A2(n848), .ZN(n850) );
  NAND2_X1 U938 ( .A1(n851), .A2(n850), .ZN(n852) );
  XNOR2_X1 U939 ( .A(n852), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U940 ( .A1(G2106), .A2(n853), .ZN(G217) );
  AND2_X1 U941 ( .A1(G15), .A2(G2), .ZN(n854) );
  NAND2_X1 U942 ( .A1(G661), .A2(n854), .ZN(G259) );
  NAND2_X1 U943 ( .A1(G3), .A2(G1), .ZN(n855) );
  NAND2_X1 U944 ( .A1(n856), .A2(n855), .ZN(G188) );
  INV_X1 U946 ( .A(G120), .ZN(G236) );
  INV_X1 U947 ( .A(G108), .ZN(G238) );
  INV_X1 U948 ( .A(G96), .ZN(G221) );
  INV_X1 U949 ( .A(G69), .ZN(G235) );
  NOR2_X1 U950 ( .A1(n858), .A2(n857), .ZN(G325) );
  INV_X1 U951 ( .A(G325), .ZN(G261) );
  INV_X1 U952 ( .A(n859), .ZN(G319) );
  XNOR2_X1 U953 ( .A(G1981), .B(KEYINPUT41), .ZN(n869) );
  XOR2_X1 U954 ( .A(G1956), .B(G1961), .Z(n861) );
  XNOR2_X1 U955 ( .A(G1986), .B(G1966), .ZN(n860) );
  XNOR2_X1 U956 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U957 ( .A(G1971), .B(G1976), .Z(n863) );
  XNOR2_X1 U958 ( .A(G1996), .B(G1991), .ZN(n862) );
  XNOR2_X1 U959 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U960 ( .A(n865), .B(n864), .Z(n867) );
  XNOR2_X1 U961 ( .A(KEYINPUT114), .B(G2474), .ZN(n866) );
  XNOR2_X1 U962 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U963 ( .A(n869), .B(n868), .ZN(G229) );
  XOR2_X1 U964 ( .A(KEYINPUT42), .B(G2090), .Z(n871) );
  XNOR2_X1 U965 ( .A(G2078), .B(G2072), .ZN(n870) );
  XNOR2_X1 U966 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U967 ( .A(n872), .B(G2100), .Z(n874) );
  XNOR2_X1 U968 ( .A(G2067), .B(G2084), .ZN(n873) );
  XNOR2_X1 U969 ( .A(n874), .B(n873), .ZN(n878) );
  XOR2_X1 U970 ( .A(G2096), .B(KEYINPUT43), .Z(n876) );
  XNOR2_X1 U971 ( .A(G2678), .B(KEYINPUT113), .ZN(n875) );
  XNOR2_X1 U972 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U973 ( .A(n878), .B(n877), .Z(G227) );
  NAND2_X1 U974 ( .A1(G124), .A2(n622), .ZN(n879) );
  XNOR2_X1 U975 ( .A(n879), .B(KEYINPUT44), .ZN(n881) );
  NAND2_X1 U976 ( .A1(n901), .A2(G112), .ZN(n880) );
  NAND2_X1 U977 ( .A1(n881), .A2(n880), .ZN(n885) );
  NAND2_X1 U978 ( .A1(G100), .A2(n618), .ZN(n883) );
  NAND2_X1 U979 ( .A1(G136), .A2(n898), .ZN(n882) );
  NAND2_X1 U980 ( .A1(n883), .A2(n882), .ZN(n884) );
  NOR2_X1 U981 ( .A1(n885), .A2(n884), .ZN(G162) );
  NAND2_X1 U982 ( .A1(G118), .A2(n901), .ZN(n887) );
  NAND2_X1 U983 ( .A1(G130), .A2(n622), .ZN(n886) );
  NAND2_X1 U984 ( .A1(n887), .A2(n886), .ZN(n892) );
  NAND2_X1 U985 ( .A1(G106), .A2(n618), .ZN(n889) );
  NAND2_X1 U986 ( .A1(G142), .A2(n898), .ZN(n888) );
  NAND2_X1 U987 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U988 ( .A(n890), .B(KEYINPUT45), .Z(n891) );
  NOR2_X1 U989 ( .A1(n892), .A2(n891), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n894), .B(n893), .ZN(n914) );
  XOR2_X1 U991 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n897) );
  XOR2_X1 U992 ( .A(G160), .B(n895), .Z(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n910) );
  NAND2_X1 U994 ( .A1(G103), .A2(n618), .ZN(n900) );
  NAND2_X1 U995 ( .A1(G139), .A2(n898), .ZN(n899) );
  NAND2_X1 U996 ( .A1(n900), .A2(n899), .ZN(n906) );
  NAND2_X1 U997 ( .A1(G115), .A2(n901), .ZN(n903) );
  NAND2_X1 U998 ( .A1(G127), .A2(n622), .ZN(n902) );
  NAND2_X1 U999 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1000 ( .A(KEYINPUT47), .B(n904), .Z(n905) );
  NOR2_X1 U1001 ( .A1(n906), .A2(n905), .ZN(n964) );
  XOR2_X1 U1002 ( .A(G164), .B(n964), .Z(n907) );
  XNOR2_X1 U1003 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(n910), .B(n909), .ZN(n912) );
  XNOR2_X1 U1005 ( .A(n980), .B(G162), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1007 ( .A(n914), .B(n913), .Z(n915) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n915), .ZN(n916) );
  XOR2_X1 U1009 ( .A(KEYINPUT115), .B(n916), .Z(G395) );
  XOR2_X1 U1010 ( .A(n917), .B(G286), .Z(n919) );
  XNOR2_X1 U1011 ( .A(G171), .B(n989), .ZN(n918) );
  XNOR2_X1 U1012 ( .A(n919), .B(n918), .ZN(n920) );
  XOR2_X1 U1013 ( .A(n1006), .B(n920), .Z(n921) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n921), .ZN(G397) );
  XOR2_X1 U1015 ( .A(G2451), .B(G2430), .Z(n923) );
  XNOR2_X1 U1016 ( .A(G2438), .B(G2443), .ZN(n922) );
  XNOR2_X1 U1017 ( .A(n923), .B(n922), .ZN(n929) );
  XOR2_X1 U1018 ( .A(G2435), .B(G2454), .Z(n925) );
  XNOR2_X1 U1019 ( .A(G1341), .B(G1348), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(n925), .B(n924), .ZN(n927) );
  XOR2_X1 U1021 ( .A(G2446), .B(G2427), .Z(n926) );
  XNOR2_X1 U1022 ( .A(n927), .B(n926), .ZN(n928) );
  XOR2_X1 U1023 ( .A(n929), .B(n928), .Z(n930) );
  NAND2_X1 U1024 ( .A1(G14), .A2(n930), .ZN(n936) );
  NAND2_X1 U1025 ( .A1(G319), .A2(n936), .ZN(n933) );
  NOR2_X1 U1026 ( .A1(G229), .A2(G227), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(KEYINPUT49), .B(n931), .ZN(n932) );
  NOR2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n935) );
  NOR2_X1 U1029 ( .A1(G395), .A2(G397), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(G225) );
  INV_X1 U1031 ( .A(G225), .ZN(G308) );
  INV_X1 U1032 ( .A(n936), .ZN(G401) );
  INV_X1 U1033 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U1034 ( .A(n937), .B(G27), .ZN(n939) );
  XOR2_X1 U1035 ( .A(G1996), .B(G32), .Z(n938) );
  NAND2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n946) );
  XNOR2_X1 U1037 ( .A(G2072), .B(KEYINPUT120), .ZN(n940) );
  XNOR2_X1 U1038 ( .A(n940), .B(G33), .ZN(n943) );
  XOR2_X1 U1039 ( .A(G2067), .B(G26), .Z(n941) );
  XNOR2_X1 U1040 ( .A(KEYINPUT119), .B(n941), .ZN(n942) );
  NOR2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1042 ( .A(n944), .B(KEYINPUT121), .ZN(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(KEYINPUT122), .B(n947), .ZN(n948) );
  NAND2_X1 U1045 ( .A1(n948), .A2(G28), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(G25), .B(G1991), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1048 ( .A(KEYINPUT53), .B(n951), .Z(n955) );
  XNOR2_X1 U1049 ( .A(KEYINPUT54), .B(G34), .ZN(n952) );
  XNOR2_X1 U1050 ( .A(n952), .B(KEYINPUT123), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(G2084), .B(n953), .ZN(n954) );
  NAND2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(G35), .B(G2090), .ZN(n956) );
  NOR2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1055 ( .A(n958), .B(KEYINPUT124), .ZN(n959) );
  NOR2_X1 U1056 ( .A1(G29), .A2(n959), .ZN(n960) );
  XNOR2_X1 U1057 ( .A(KEYINPUT55), .B(n960), .ZN(n1044) );
  INV_X1 U1058 ( .A(n961), .ZN(n963) );
  NOR2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n985) );
  XOR2_X1 U1060 ( .A(G2072), .B(n964), .Z(n966) );
  XOR2_X1 U1061 ( .A(G164), .B(G2078), .Z(n965) );
  NOR2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1063 ( .A(KEYINPUT118), .B(n967), .ZN(n968) );
  XNOR2_X1 U1064 ( .A(n968), .B(KEYINPUT50), .ZN(n978) );
  XNOR2_X1 U1065 ( .A(G160), .B(G2084), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(G2090), .B(G162), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(n971), .B(KEYINPUT117), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(KEYINPUT51), .B(n974), .ZN(n975) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n983) );
  NOR2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1074 ( .A(KEYINPUT116), .B(n981), .Z(n982) );
  NOR2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(KEYINPUT52), .B(n986), .ZN(n987) );
  NAND2_X1 U1078 ( .A1(n987), .A2(G29), .ZN(n988) );
  NAND2_X1 U1079 ( .A1(G11), .A2(n988), .ZN(n1042) );
  XNOR2_X1 U1080 ( .A(G16), .B(KEYINPUT56), .ZN(n1013) );
  XNOR2_X1 U1081 ( .A(n989), .B(G1348), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(G301), .B(G1961), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(G299), .B(G1956), .ZN(n990) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n1011) );
  XOR2_X1 U1087 ( .A(G1966), .B(G168), .Z(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1089 ( .A(KEYINPUT57), .B(n998), .Z(n1005) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  AND2_X1 U1091 ( .A1(G303), .A2(G1971), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1093 ( .A(KEYINPUT125), .B(n1003), .Z(n1004) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1009) );
  XOR2_X1 U1095 ( .A(G1341), .B(n1006), .Z(n1007) );
  XNOR2_X1 U1096 ( .A(KEYINPUT126), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1040) );
  INV_X1 U1100 ( .A(G16), .ZN(n1038) );
  XNOR2_X1 U1101 ( .A(G5), .B(n1014), .ZN(n1027) );
  INV_X1 U1102 ( .A(G1341), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(G19), .B(n1015), .ZN(n1019) );
  XNOR2_X1 U1104 ( .A(G1981), .B(G6), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(G20), .B(G1956), .ZN(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1022) );
  XOR2_X1 U1108 ( .A(KEYINPUT59), .B(G1348), .Z(n1020) );
  XNOR2_X1 U1109 ( .A(G4), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1111 ( .A(KEYINPUT60), .B(n1023), .Z(n1025) );
  XNOR2_X1 U1112 ( .A(G1966), .B(G21), .ZN(n1024) );
  NOR2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1035) );
  XNOR2_X1 U1115 ( .A(G1986), .B(G24), .ZN(n1029) );
  XNOR2_X1 U1116 ( .A(G22), .B(G1971), .ZN(n1028) );
  NOR2_X1 U1117 ( .A1(n1029), .A2(n1028), .ZN(n1032) );
  XNOR2_X1 U1118 ( .A(G1976), .B(KEYINPUT127), .ZN(n1030) );
  XNOR2_X1 U1119 ( .A(n1030), .B(G23), .ZN(n1031) );
  NAND2_X1 U1120 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1121 ( .A(KEYINPUT58), .B(n1033), .ZN(n1034) );
  NOR2_X1 U1122 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1123 ( .A(KEYINPUT61), .B(n1036), .ZN(n1037) );
  NAND2_X1 U1124 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NAND2_X1 U1125 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  NOR2_X1 U1126 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  NAND2_X1 U1127 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  XOR2_X1 U1128 ( .A(KEYINPUT62), .B(n1045), .Z(G311) );
  INV_X1 U1129 ( .A(G311), .ZN(G150) );
endmodule

