//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  AND2_X1   g001(.A1(KEYINPUT66), .A2(G128), .ZN(new_n188));
  NOR2_X1   g002(.A1(KEYINPUT66), .A2(G128), .ZN(new_n189));
  OAI211_X1 g003(.A(KEYINPUT23), .B(G119), .C1(new_n188), .C2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT72), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT66), .B(G128), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n193), .A2(KEYINPUT72), .A3(KEYINPUT23), .A4(G119), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  AOI21_X1  g009(.A(KEYINPUT23), .B1(new_n195), .B2(G119), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(G119), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n192), .A2(new_n194), .A3(new_n198), .ZN(new_n199));
  XOR2_X1   g013(.A(KEYINPUT77), .B(G110), .Z(new_n200));
  AOI21_X1  g014(.A(new_n197), .B1(new_n193), .B2(G119), .ZN(new_n201));
  XOR2_X1   g015(.A(KEYINPUT24), .B(G110), .Z(new_n202));
  OAI22_X1  g016(.A1(new_n199), .A2(new_n200), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  AND2_X1   g017(.A1(KEYINPUT74), .A2(G140), .ZN(new_n204));
  NOR2_X1   g018(.A1(KEYINPUT74), .A2(G140), .ZN(new_n205));
  OAI21_X1  g019(.A(G125), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT75), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G125), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n209), .A2(KEYINPUT76), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(KEYINPUT76), .ZN(new_n211));
  OAI21_X1  g025(.A(G140), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OAI211_X1 g026(.A(KEYINPUT75), .B(G125), .C1(new_n204), .C2(new_n205), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n208), .A2(KEYINPUT16), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  OR4_X1    g028(.A1(KEYINPUT16), .A2(new_n210), .A3(new_n211), .A4(G140), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(G146), .ZN(new_n216));
  XOR2_X1   g030(.A(G125), .B(G140), .Z(new_n217));
  OAI211_X1 g031(.A(new_n203), .B(new_n216), .C1(G146), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n201), .A2(new_n202), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n214), .A2(G146), .A3(new_n215), .ZN(new_n220));
  AOI21_X1  g034(.A(G146), .B1(new_n214), .B2(new_n215), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT73), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n199), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n192), .A2(new_n194), .A3(KEYINPUT73), .A4(new_n198), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(G110), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  OAI211_X1 g041(.A(KEYINPUT78), .B(new_n218), .C1(new_n222), .C2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G953), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(G221), .A3(G234), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n230), .B(KEYINPUT22), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n231), .B(G137), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n228), .A2(new_n233), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n226), .B(new_n219), .C1(new_n221), .C2(new_n220), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT78), .B1(new_n235), .B2(new_n218), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n218), .B1(new_n222), .B2(new_n227), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT78), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(new_n239), .A3(new_n232), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n187), .B1(new_n237), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT25), .ZN(new_n243));
  INV_X1    g057(.A(G217), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(G234), .B2(new_n187), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n238), .A2(new_n239), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(new_n228), .A3(new_n233), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n240), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT25), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n249), .A3(new_n187), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n243), .A2(new_n245), .A3(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n245), .A2(G902), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT79), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n251), .A2(KEYINPUT79), .A3(new_n253), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT31), .ZN(new_n259));
  INV_X1    g073(.A(G146), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G143), .ZN(new_n261));
  INV_X1    g075(.A(G143), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G146), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT1), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n265), .B1(G143), .B2(new_n260), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n264), .B1(new_n193), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT67), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n261), .A2(new_n263), .A3(new_n265), .A4(G128), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n264), .B(KEYINPUT67), .C1(new_n193), .C2(new_n266), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AND2_X1   g086(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n273));
  NOR2_X1   g087(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G134), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(G137), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT65), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n276), .A2(G137), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n279), .B1(KEYINPUT11), .B2(new_n277), .ZN(new_n280));
  INV_X1    g094(.A(G131), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT65), .ZN(new_n282));
  OAI221_X1 g096(.A(new_n282), .B1(new_n276), .B2(G137), .C1(new_n273), .C2(new_n274), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n278), .A2(new_n280), .A3(new_n281), .A4(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(G131), .B1(new_n279), .B2(new_n277), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n272), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  OR2_X1    g100(.A1(KEYINPUT0), .A2(G128), .ZN(new_n287));
  NAND2_X1  g101(.A1(KEYINPUT0), .A2(G128), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n264), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n261), .A2(new_n263), .A3(KEYINPUT0), .A4(G128), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n278), .A2(new_n280), .A3(new_n283), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G131), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n291), .B1(new_n293), .B2(new_n284), .ZN(new_n294));
  INV_X1    g108(.A(G119), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G116), .ZN(new_n296));
  INV_X1    g110(.A(G116), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G119), .ZN(new_n298));
  INV_X1    g112(.A(G113), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n299), .A2(KEYINPUT2), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n299), .A2(KEYINPUT2), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n296), .B(new_n298), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n296), .A2(new_n298), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT2), .B(G113), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n286), .A2(new_n294), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n293), .A2(new_n284), .ZN(new_n308));
  INV_X1    g122(.A(new_n291), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT30), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n272), .A2(new_n284), .A3(new_n285), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT30), .B1(new_n286), .B2(new_n294), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n307), .B1(new_n315), .B2(new_n306), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT26), .B(G101), .Z(new_n317));
  NOR2_X1   g131(.A1(G237), .A2(G953), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G210), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n317), .B(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n320), .B(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n259), .B1(new_n316), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n306), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(new_n313), .B2(new_n314), .ZN(new_n326));
  NOR4_X1   g140(.A1(new_n326), .A2(KEYINPUT31), .A3(new_n322), .A4(new_n307), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n310), .A2(new_n325), .A3(new_n312), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n306), .B1(new_n286), .B2(new_n294), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n323), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NOR3_X1   g149(.A1(new_n324), .A2(new_n327), .A3(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(G472), .A2(G902), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT32), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n315), .A2(new_n306), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n323), .A3(new_n328), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT31), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n332), .A2(new_n334), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n322), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n316), .A2(new_n259), .A3(new_n323), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT32), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n347), .A3(new_n337), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n339), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n332), .A2(new_n323), .A3(new_n334), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n322), .B1(new_n326), .B2(new_n307), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT29), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT70), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT71), .ZN(new_n356));
  INV_X1    g170(.A(new_n334), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n333), .B1(new_n328), .B2(new_n329), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n323), .A2(KEYINPUT29), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n356), .B(new_n187), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NOR3_X1   g175(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT71), .B1(new_n362), .B2(G902), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT70), .A4(new_n352), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n355), .A2(new_n361), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G472), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n349), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n258), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n258), .A2(KEYINPUT80), .A3(new_n367), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n193), .A2(G143), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n195), .A2(G143), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n373), .A2(new_n276), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G122), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G116), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n297), .A2(G122), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G107), .ZN(new_n381));
  INV_X1    g195(.A(G107), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n378), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT13), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n385), .B1(new_n193), .B2(G143), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT96), .ZN(new_n387));
  OR3_X1    g201(.A1(new_n386), .A2(new_n387), .A3(new_n374), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n375), .A2(new_n385), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n387), .B1(new_n386), .B2(new_n374), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n388), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n376), .B(new_n384), .C1(new_n392), .C2(new_n276), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n297), .A2(KEYINPUT14), .A3(G122), .ZN(new_n394));
  OAI211_X1 g208(.A(G107), .B(new_n394), .C1(new_n380), .C2(KEYINPUT14), .ZN(new_n395));
  XOR2_X1   g209(.A(new_n395), .B(KEYINPUT97), .Z(new_n396));
  INV_X1    g210(.A(new_n376), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n276), .B1(new_n373), .B2(new_n375), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n396), .B(new_n383), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  XOR2_X1   g213(.A(KEYINPUT9), .B(G234), .Z(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n401), .A2(new_n244), .A3(G953), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n393), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n402), .B1(new_n393), .B2(new_n399), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n187), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT98), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n393), .A2(new_n399), .ZN(new_n408));
  INV_X1    g222(.A(new_n402), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n403), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT98), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n412), .A3(new_n187), .ZN(new_n413));
  INV_X1    g227(.A(G478), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(KEYINPUT15), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n407), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  OR2_X1    g230(.A1(new_n406), .A2(new_n415), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G475), .ZN(new_n420));
  XNOR2_X1  g234(.A(G113), .B(G122), .ZN(new_n421));
  INV_X1    g235(.A(G104), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n421), .B(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT93), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G143), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n262), .A2(KEYINPUT93), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n425), .A2(new_n426), .A3(G214), .A4(new_n318), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n318), .A2(G214), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n427), .B1(new_n428), .B2(new_n425), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(G131), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n217), .A2(KEYINPUT19), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n208), .A2(new_n212), .A3(new_n213), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT94), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n434), .B(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT19), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n433), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n216), .B(new_n431), .C1(new_n438), .C2(G146), .ZN(new_n439));
  AND2_X1   g253(.A1(KEYINPUT18), .A2(G131), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n429), .B(new_n440), .ZN(new_n441));
  OR2_X1    g255(.A1(new_n434), .A2(KEYINPUT94), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n434), .A2(KEYINPUT94), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n260), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n217), .A2(G146), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n441), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n423), .B1(new_n439), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n220), .A2(new_n221), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT17), .ZN(new_n449));
  OR3_X1    g263(.A1(new_n429), .A2(new_n449), .A3(new_n281), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n430), .A2(new_n449), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n448), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n446), .A2(new_n452), .A3(new_n423), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n420), .B(new_n187), .C1(new_n447), .C2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT20), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n423), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n431), .A2(new_n216), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n442), .A2(new_n443), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n432), .B1(new_n460), .B2(KEYINPUT19), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n459), .B1(new_n461), .B2(new_n260), .ZN(new_n462));
  INV_X1    g276(.A(new_n446), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n458), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n453), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n465), .A2(KEYINPUT20), .A3(new_n420), .A4(new_n187), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n423), .B1(new_n446), .B2(new_n452), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n187), .B1(new_n454), .B2(new_n467), .ZN(new_n468));
  XOR2_X1   g282(.A(KEYINPUT95), .B(G475), .Z(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n457), .A2(new_n466), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n419), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G214), .B1(G237), .B2(G902), .ZN(new_n474));
  XNOR2_X1  g288(.A(G110), .B(G122), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G101), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n422), .A2(new_n382), .ZN(new_n478));
  OR2_X1    g292(.A1(KEYINPUT81), .A2(G104), .ZN(new_n479));
  NAND2_X1  g293(.A1(KEYINPUT81), .A2(G104), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI211_X1 g295(.A(new_n477), .B(new_n478), .C1(new_n481), .C2(new_n382), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n296), .A2(new_n298), .A3(KEYINPUT5), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(G113), .B1(new_n296), .B2(KEYINPUT5), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n302), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g300(.A1(KEYINPUT3), .A2(G107), .ZN(new_n487));
  NOR2_X1   g301(.A1(KEYINPUT3), .A2(G107), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n487), .B1(G104), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT3), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n382), .ZN(new_n491));
  AND2_X1   g305(.A1(KEYINPUT81), .A2(G104), .ZN(new_n492));
  NOR2_X1   g306(.A1(KEYINPUT81), .A2(G104), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT82), .B(G101), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n489), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT83), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n489), .A2(new_n494), .A3(KEYINPUT83), .A4(new_n495), .ZN(new_n499));
  AOI211_X1 g313(.A(new_n482), .B(new_n486), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT4), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n488), .B1(new_n479), .B2(new_n480), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n490), .A2(new_n382), .A3(G104), .ZN(new_n503));
  NAND2_X1  g317(.A1(KEYINPUT3), .A2(G107), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n501), .B(G101), .C1(new_n502), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n306), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n498), .A2(new_n499), .ZN(new_n508));
  OAI21_X1  g322(.A(G101), .B1(new_n502), .B2(new_n505), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n509), .A2(KEYINPUT4), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n507), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n476), .B1(new_n500), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n482), .ZN(new_n513));
  INV_X1    g327(.A(new_n486), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n508), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n509), .A2(KEYINPUT4), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n516), .B1(new_n498), .B2(new_n499), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n515), .B(new_n475), .C1(new_n517), .C2(new_n507), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n512), .A2(KEYINPUT6), .A3(new_n518), .ZN(new_n519));
  XOR2_X1   g333(.A(KEYINPUT76), .B(G125), .Z(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n291), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT89), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n269), .A2(new_n270), .A3(new_n271), .A4(new_n520), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT89), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n291), .A2(new_n525), .A3(new_n521), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G224), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(G953), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n527), .B(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT6), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n531), .B(new_n476), .C1(new_n500), .C2(new_n511), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n519), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT90), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n519), .A2(new_n530), .A3(new_n532), .A4(KEYINPUT90), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT91), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n483), .B1(new_n485), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n297), .A2(G119), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT5), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n299), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(KEYINPUT91), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n302), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n508), .A2(new_n544), .A3(new_n513), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n475), .B(KEYINPUT8), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n482), .B1(new_n498), .B2(new_n499), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n545), .B(new_n546), .C1(new_n547), .C2(new_n486), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n524), .A2(new_n522), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT7), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n549), .B1(new_n550), .B2(new_n529), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n525), .B1(new_n291), .B2(new_n521), .ZN(new_n552));
  AOI211_X1 g366(.A(KEYINPUT89), .B(new_n520), .C1(new_n289), .C2(new_n290), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n529), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n554), .A2(KEYINPUT7), .A3(new_n524), .A4(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n548), .A2(new_n518), .A3(new_n551), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n187), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT92), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n557), .A2(KEYINPUT92), .A3(new_n187), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(G210), .B1(G237), .B2(G902), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n537), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n563), .B1(new_n537), .B2(new_n562), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n474), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT99), .B(G952), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(G953), .ZN(new_n568));
  NAND2_X1  g382(.A1(G234), .A2(G237), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n569), .A2(G902), .A3(G953), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT21), .B(G898), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT100), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  OR3_X1    g390(.A1(new_n473), .A2(new_n566), .A3(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(G110), .B(G140), .Z(new_n578));
  AND2_X1   g392(.A1(new_n229), .A2(G227), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n308), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT84), .ZN(new_n583));
  INV_X1    g397(.A(new_n506), .ZN(new_n584));
  NOR4_X1   g398(.A1(new_n517), .A2(new_n583), .A3(new_n291), .A4(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n584), .B1(new_n508), .B2(new_n510), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT84), .B1(new_n586), .B2(new_n309), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n272), .A2(KEYINPUT10), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n264), .B1(new_n266), .B2(new_n195), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT85), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT85), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n264), .B(new_n592), .C1(new_n195), .C2(new_n266), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(new_n593), .A3(new_n270), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n508), .A2(new_n594), .A3(new_n513), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT10), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n547), .A2(new_n589), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n582), .B1(new_n588), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n508), .A2(new_n510), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n599), .A2(new_n309), .A3(new_n506), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n583), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n586), .A2(KEYINPUT84), .A3(new_n309), .ZN(new_n602));
  AND4_X1   g416(.A1(new_n582), .A2(new_n597), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n581), .B1(new_n598), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT87), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT87), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n606), .B(new_n581), .C1(new_n598), .C2(new_n603), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n603), .A2(new_n581), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n595), .B1(new_n547), .B2(new_n272), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT12), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n609), .A2(KEYINPUT86), .A3(new_n610), .A4(new_n308), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT86), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n609), .A2(new_n308), .B1(new_n612), .B2(KEYINPUT12), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n613), .B1(new_n612), .B2(KEYINPUT12), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n608), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n605), .A2(new_n607), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(G469), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n617), .A3(new_n187), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n597), .A2(new_n601), .A3(new_n582), .A4(new_n602), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n614), .A2(new_n619), .A3(new_n611), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n581), .ZN(new_n621));
  INV_X1    g435(.A(new_n598), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n608), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(new_n623), .A3(G469), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n617), .A2(new_n187), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n618), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(G221), .B1(new_n401), .B2(G902), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT88), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT88), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n627), .A2(new_n631), .A3(new_n628), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n577), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n372), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n634), .B(new_n495), .Z(G3));
  NAND2_X1  g449(.A1(new_n630), .A2(new_n632), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n251), .A2(KEYINPUT79), .A3(new_n253), .ZN(new_n637));
  AOI21_X1  g451(.A(KEYINPUT79), .B1(new_n251), .B2(new_n253), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(G472), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n346), .B2(new_n187), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n324), .A2(new_n327), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n338), .B1(new_n642), .B2(new_n344), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT101), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(G472), .B1(new_n336), .B2(G902), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n639), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n636), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n566), .A2(KEYINPUT102), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n652), .B(new_n474), .C1(new_n564), .C2(new_n565), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n407), .A2(new_n413), .A3(new_n414), .ZN(new_n656));
  NAND2_X1  g470(.A1(KEYINPUT103), .A2(KEYINPUT33), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n411), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT103), .B(KEYINPUT33), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n410), .A2(new_n403), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n658), .A2(new_n187), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n656), .B1(new_n414), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n471), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n576), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n655), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n650), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT104), .B(KEYINPUT34), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n422), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n666), .B(new_n668), .ZN(G6));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n418), .A2(new_n457), .A3(new_n466), .A4(new_n470), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n670), .B1(new_n671), .B2(new_n576), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n472), .A2(KEYINPUT105), .A3(new_n575), .A4(new_n418), .ZN(new_n673));
  AOI211_X1 g487(.A(new_n654), .B(new_n650), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT35), .B(G107), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  AOI21_X1  g490(.A(new_n249), .B1(new_n248), .B2(new_n187), .ZN(new_n677));
  AOI211_X1 g491(.A(KEYINPUT25), .B(G902), .C1(new_n247), .C2(new_n240), .ZN(new_n678));
  INV_X1    g492(.A(new_n245), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n233), .A2(KEYINPUT36), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n238), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n252), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(KEYINPUT106), .B1(new_n680), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n251), .A2(new_n686), .A3(new_n683), .ZN(new_n687));
  AND4_X1   g501(.A1(new_n644), .A2(new_n685), .A3(new_n647), .A4(new_n687), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n473), .A2(new_n566), .A3(new_n576), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n627), .A2(new_n631), .A3(new_n628), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n631), .B1(new_n627), .B2(new_n628), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n688), .B(new_n689), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n692), .B(KEYINPUT37), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G110), .ZN(G12));
  NAND3_X1  g508(.A1(new_n367), .A2(new_n685), .A3(new_n687), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n654), .ZN(new_n696));
  INV_X1    g510(.A(G900), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n571), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n570), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n671), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n636), .A2(new_n696), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G128), .ZN(G30));
  XNOR2_X1  g516(.A(new_n699), .B(KEYINPUT39), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n703), .B1(new_n630), .B2(new_n632), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT40), .ZN(new_n705));
  AOI211_X1 g519(.A(new_n472), .B(new_n419), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n251), .A2(new_n686), .A3(new_n683), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n686), .B1(new_n251), .B2(new_n683), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n474), .ZN(new_n711));
  INV_X1    g525(.A(new_n703), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n636), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n711), .B1(new_n713), .B2(KEYINPUT40), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n316), .A2(new_n322), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n187), .B1(new_n330), .B2(new_n323), .ZN(new_n716));
  OAI21_X1  g530(.A(G472), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n349), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n349), .A2(KEYINPUT107), .A3(new_n717), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n565), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n537), .A2(new_n562), .A3(new_n563), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n726), .B(KEYINPUT38), .Z(new_n727));
  NOR2_X1   g541(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n706), .A2(new_n710), .A3(new_n714), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G143), .ZN(G45));
  INV_X1    g544(.A(new_n699), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n662), .A2(new_n471), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n636), .A2(new_n696), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT108), .B(G146), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G48));
  NAND2_X1  g550(.A1(new_n616), .A2(new_n187), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(G469), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n628), .A3(new_n618), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n665), .A2(new_n368), .A3(new_n739), .ZN(new_n740));
  XOR2_X1   g554(.A(KEYINPUT41), .B(G113), .Z(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  AOI22_X1  g556(.A1(new_n339), .A2(new_n348), .B1(new_n365), .B2(G472), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n639), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n672), .A2(new_n673), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n738), .A2(new_n628), .A3(new_n618), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n744), .A2(new_n745), .A3(new_n655), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G116), .ZN(G18));
  NOR3_X1   g562(.A1(new_n743), .A2(new_n707), .A3(new_n708), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n473), .A2(new_n576), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n749), .A2(new_n655), .A3(new_n750), .A4(new_n746), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT109), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G119), .ZN(G21));
  AND2_X1   g567(.A1(new_n418), .A2(new_n471), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n651), .A2(new_n653), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT111), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n651), .A2(new_n754), .A3(new_n757), .A4(new_n653), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n254), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n346), .A2(new_n187), .ZN(new_n761));
  XOR2_X1   g575(.A(KEYINPUT110), .B(G472), .Z(new_n762));
  NAND2_X1  g576(.A1(new_n359), .A2(new_n322), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n642), .A2(new_n763), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n761), .A2(new_n762), .B1(new_n764), .B2(new_n337), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n739), .A2(new_n766), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n759), .A2(new_n575), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n377), .ZN(G24));
  NOR2_X1   g583(.A1(new_n654), .A2(new_n739), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n685), .A2(new_n687), .A3(new_n765), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n770), .A2(new_n733), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G125), .ZN(G27));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n624), .A2(KEYINPUT112), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n624), .A2(KEYINPUT112), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n618), .B(new_n626), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n628), .A2(new_n474), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n726), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n258), .A2(new_n367), .A3(new_n778), .A4(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n775), .B1(new_n781), .B2(new_n732), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n778), .A2(new_n780), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n744), .A2(new_n783), .A3(KEYINPUT113), .A4(new_n733), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT42), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n743), .A2(new_n254), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n783), .A2(KEYINPUT42), .A3(new_n733), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT114), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G131), .ZN(G33));
  NOR3_X1   g605(.A1(new_n781), .A2(new_n671), .A3(new_n699), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(new_n276), .ZN(G36));
  INV_X1    g607(.A(KEYINPUT46), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n621), .A2(new_n623), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT45), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n796), .A2(G469), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n794), .B1(new_n797), .B2(new_n625), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(G469), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(KEYINPUT46), .A3(new_n626), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n798), .A2(new_n618), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n628), .A3(new_n712), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n802), .A2(KEYINPUT115), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n472), .A2(new_n662), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT43), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n805), .B1(new_n471), .B2(KEYINPUT116), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n804), .A2(new_n806), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n648), .A3(new_n709), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT44), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n802), .A2(KEYINPUT115), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n803), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n810), .A2(new_n811), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n726), .A2(new_n711), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G137), .ZN(G39));
  NAND2_X1  g634(.A1(new_n801), .A2(new_n628), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT47), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n801), .A2(KEYINPUT47), .A3(new_n628), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n367), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n258), .A2(new_n817), .A3(new_n732), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G140), .ZN(G42));
  NAND2_X1  g642(.A1(new_n738), .A2(new_n618), .ZN(new_n829));
  OR3_X1    g643(.A1(new_n829), .A2(KEYINPUT117), .A3(KEYINPUT49), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n723), .A2(new_n830), .A3(new_n804), .ZN(new_n831));
  AOI211_X1 g645(.A(new_n779), .B(new_n254), .C1(KEYINPUT117), .C2(KEYINPUT49), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n829), .B1(KEYINPUT117), .B2(KEYINPUT49), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n831), .A2(new_n727), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n654), .A2(new_n771), .A3(new_n739), .A4(new_n732), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n709), .A2(new_n367), .A3(new_n651), .A4(new_n653), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(new_n632), .B2(new_n630), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n836), .B1(new_n838), .B2(new_n700), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n251), .A2(new_n778), .A3(new_n683), .A4(new_n731), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n759), .A2(new_n628), .A3(new_n722), .A4(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n839), .A2(KEYINPUT52), .A3(new_n734), .A4(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n841), .A2(new_n701), .A3(new_n734), .A4(new_n773), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n842), .A2(new_n845), .A3(KEYINPUT120), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT120), .B1(new_n842), .B2(new_n845), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n747), .A2(new_n751), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n768), .A2(new_n849), .A3(new_n740), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n792), .B1(new_n786), .B2(new_n788), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n783), .A2(new_n733), .A3(new_n765), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n473), .A2(new_n699), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n367), .B(new_n853), .C1(new_n690), .C2(new_n691), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n852), .B1(new_n854), .B2(new_n817), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n709), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n850), .A2(new_n851), .A3(new_n856), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n644), .B(new_n647), .C1(new_n637), .C2(new_n638), .ZN(new_n858));
  AOI211_X1 g672(.A(new_n566), .B(new_n858), .C1(new_n630), .C2(new_n632), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n859), .A2(new_n664), .B1(new_n372), .B2(new_n633), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n671), .A2(new_n566), .A3(new_n576), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n649), .B(new_n862), .C1(new_n690), .C2(new_n691), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT118), .B1(new_n863), .B2(new_n692), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n863), .A2(new_n692), .A3(KEYINPUT118), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n860), .B(new_n861), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n863), .A2(new_n692), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n863), .A2(new_n692), .A3(KEYINPUT118), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n861), .B1(new_n872), .B2(new_n860), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n857), .B1(new_n867), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n835), .B1(new_n848), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n850), .A2(new_n851), .A3(new_n856), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n860), .B1(new_n865), .B2(new_n864), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT119), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n877), .B1(new_n879), .B2(new_n866), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n842), .A2(new_n845), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(KEYINPUT53), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n875), .A2(new_n876), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n843), .A2(new_n844), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n843), .A2(new_n844), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n842), .A2(new_n845), .A3(KEYINPUT120), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n889), .A2(KEYINPUT53), .A3(new_n880), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n881), .B(new_n857), .C1(new_n867), .C2(new_n873), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n835), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  AOI22_X1  g707(.A1(new_n883), .A2(KEYINPUT121), .B1(KEYINPUT54), .B2(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n893), .A2(KEYINPUT121), .A3(KEYINPUT54), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n829), .A2(new_n726), .A3(new_n779), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n639), .A2(new_n570), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n723), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n898), .A2(new_n471), .A3(new_n662), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n570), .B1(new_n807), .B2(new_n808), .ZN(new_n900));
  INV_X1    g714(.A(new_n766), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n746), .A2(KEYINPUT122), .A3(new_n711), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n739), .A2(new_n474), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n727), .B1(new_n904), .B2(KEYINPUT122), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT50), .ZN(new_n906));
  OR3_X1    g720(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n906), .B1(new_n903), .B2(new_n905), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n899), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n900), .A2(new_n896), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n772), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n829), .A2(new_n628), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n823), .A2(new_n824), .A3(new_n912), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n900), .A2(new_n901), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n914), .A2(new_n816), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n909), .A2(new_n911), .A3(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT51), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n913), .A2(KEYINPUT123), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n823), .A2(new_n921), .A3(new_n824), .A4(new_n912), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n920), .A2(new_n915), .A3(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n923), .A2(KEYINPUT51), .A3(new_n911), .A4(new_n909), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n919), .A2(new_n924), .A3(new_n568), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n910), .A2(new_n787), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT48), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n898), .A2(new_n663), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n914), .A2(new_n770), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n925), .A2(new_n927), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n894), .A2(new_n895), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(G952), .A2(G953), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n834), .B1(new_n931), .B2(new_n932), .ZN(G75));
  AOI21_X1  g747(.A(new_n187), .B1(new_n875), .B2(new_n882), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(G210), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT56), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n519), .A2(new_n532), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(new_n530), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT55), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n935), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n939), .B1(new_n935), .B2(new_n936), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n229), .A2(G952), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(G51));
  OR2_X1    g757(.A1(new_n626), .A2(KEYINPUT57), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n626), .A2(KEYINPUT57), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT53), .B1(new_n889), .B2(new_n880), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n891), .A2(new_n835), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n946), .A2(new_n947), .A3(KEYINPUT54), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n876), .B1(new_n875), .B2(new_n882), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n944), .B(new_n945), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n616), .ZN(new_n951));
  OAI211_X1 g765(.A(G902), .B(new_n797), .C1(new_n946), .C2(new_n947), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT124), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n942), .B1(new_n951), .B2(new_n953), .ZN(G54));
  INV_X1    g768(.A(new_n942), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n934), .A2(KEYINPUT58), .A3(G475), .ZN(new_n956));
  INV_X1    g770(.A(new_n465), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI211_X1 g772(.A(KEYINPUT58), .B(G902), .C1(new_n946), .C2(new_n947), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n959), .B2(new_n420), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n956), .A2(KEYINPUT125), .A3(new_n957), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n958), .B1(new_n962), .B2(new_n963), .ZN(G60));
  NAND2_X1  g778(.A1(new_n658), .A2(new_n660), .ZN(new_n965));
  NAND2_X1  g779(.A1(G478), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT59), .Z(new_n967));
  NOR2_X1   g781(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n948), .B2(new_n949), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n955), .ZN(new_n970));
  INV_X1    g784(.A(new_n967), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(new_n894), .B2(new_n895), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n970), .B1(new_n965), .B2(new_n972), .ZN(G63));
  INV_X1    g787(.A(KEYINPUT61), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n875), .A2(new_n882), .ZN(new_n975));
  NAND2_X1  g789(.A1(G217), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT60), .Z(new_n977));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n682), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n955), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n248), .B1(new_n975), .B2(new_n977), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n974), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n980), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n982), .A2(KEYINPUT61), .A3(new_n955), .A4(new_n978), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n981), .A2(new_n983), .ZN(G66));
  OAI21_X1  g798(.A(G953), .B1(new_n572), .B2(new_n528), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n879), .A2(new_n866), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n986), .A2(new_n850), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n985), .B1(new_n987), .B2(G953), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n937), .B1(G898), .B2(new_n229), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n988), .B(new_n989), .ZN(G69));
  AOI22_X1  g804(.A1(new_n814), .A2(new_n818), .B1(new_n825), .B2(new_n826), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n839), .A2(new_n734), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n803), .A2(new_n759), .A3(new_n787), .A4(new_n813), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n991), .A2(new_n992), .A3(new_n851), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n229), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n229), .A2(G900), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT127), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n315), .B(KEYINPUT126), .Z(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(new_n461), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1000), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n729), .A2(new_n992), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT62), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n817), .B1(new_n663), .B2(new_n671), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n372), .A2(new_n704), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1005), .A2(new_n991), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1002), .B1(new_n1009), .B2(G953), .ZN(new_n1010));
  NAND2_X1  g824(.A1(G227), .A2(G900), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(G953), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1001), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  OAI211_X1 g827(.A(G953), .B(new_n1011), .C1(new_n998), .C2(new_n1002), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(G72));
  INV_X1    g829(.A(new_n715), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n316), .A2(new_n322), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(G472), .A2(G902), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n1020), .B(KEYINPUT63), .Z(new_n1021));
  NOR2_X1   g835(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  OAI22_X1  g836(.A1(new_n1008), .A2(new_n1016), .B1(new_n994), .B2(new_n1017), .ZN(new_n1023));
  AOI211_X1 g837(.A(new_n942), .B(new_n1022), .C1(new_n1023), .C2(new_n987), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n893), .A2(new_n1021), .A3(new_n1019), .ZN(new_n1025));
  AND2_X1   g839(.A1(new_n1024), .A2(new_n1025), .ZN(G57));
endmodule


