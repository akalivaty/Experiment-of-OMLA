//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n823, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n202));
  AND2_X1   g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G141gat), .ZN(new_n206));
  INV_X1    g005(.A(G148gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(KEYINPUT73), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n205), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AND2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n208), .B(new_n209), .C1(new_n213), .C2(new_n214), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT74), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(new_n213), .B2(new_n211), .ZN(new_n220));
  NAND2_X1  g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(KEYINPUT74), .A3(KEYINPUT2), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n216), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G113gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT68), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT68), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G113gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n229), .A3(G120gat), .ZN(new_n230));
  INV_X1    g029(.A(G120gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G113gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G127gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G134gat), .ZN(new_n235));
  INV_X1    g034(.A(G134gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G127gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT1), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n233), .A2(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n226), .A2(G120gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n231), .A2(G113gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n238), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n247));
  NOR3_X1   g046(.A1(new_n246), .A2(new_n247), .A3(new_n234), .ZN(new_n248));
  INV_X1    g047(.A(new_n235), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n244), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n241), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT4), .B1(new_n225), .B2(new_n251), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n215), .A2(new_n212), .B1(new_n218), .B2(new_n223), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n239), .B1(new_n232), .B2(new_n230), .ZN(new_n254));
  OR2_X1    g053(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(G127gat), .A3(new_n245), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n226), .A2(G120gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n232), .A2(new_n257), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n256), .A2(new_n235), .B1(new_n258), .B2(new_n238), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n253), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT78), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n252), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n215), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n208), .A2(new_n209), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT2), .B1(new_n266), .B2(new_n202), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n265), .B1(new_n267), .B2(new_n210), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n217), .B1(new_n220), .B2(new_n222), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT3), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT3), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n216), .A2(new_n271), .A3(new_n224), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT75), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(new_n254), .B2(new_n259), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n241), .A2(new_n250), .A3(KEYINPUT75), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n270), .A2(new_n272), .A3(new_n274), .A4(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n253), .A2(new_n260), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(KEYINPUT78), .A3(KEYINPUT4), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n264), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G225gat), .A2(G233gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n274), .A2(new_n225), .A3(new_n275), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(new_n277), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n282), .B(KEYINPUT39), .C1(new_n281), .C2(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(G1gat), .B(G29gat), .Z(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G57gat), .B(G85gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n285), .B(new_n290), .C1(KEYINPUT39), .C2(new_n282), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT40), .ZN(new_n292));
  OR2_X1    g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n290), .ZN(new_n294));
  XOR2_X1   g093(.A(KEYINPUT76), .B(KEYINPUT5), .Z(new_n295));
  AOI21_X1  g094(.A(new_n295), .B1(new_n284), .B2(new_n281), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n252), .A2(new_n262), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n297), .A2(new_n276), .A3(new_n280), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n264), .A2(new_n278), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n276), .A2(new_n280), .A3(new_n295), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n294), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n291), .A2(new_n292), .ZN(new_n304));
  XOR2_X1   g103(.A(G211gat), .B(G218gat), .Z(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(G197gat), .A2(G204gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(G197gat), .A2(G204gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n310));
  NOR3_X1   g109(.A1(new_n309), .A2(KEYINPUT70), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT70), .ZN(new_n312));
  XNOR2_X1  g111(.A(G197gat), .B(G204gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n310), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n306), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n313), .A2(new_n312), .A3(new_n314), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(new_n305), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321));
  INV_X1    g120(.A(G169gat), .ZN(new_n322));
  INV_X1    g121(.A(G176gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT26), .ZN(new_n325));
  NAND2_X1  g124(.A1(G169gat), .A2(G176gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT26), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n325), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT27), .B(G183gat), .ZN(new_n331));
  INV_X1    g130(.A(G190gat), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT28), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G183gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT27), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT27), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G183gat), .ZN(new_n337));
  AND4_X1   g136(.A1(KEYINPUT28), .A2(new_n335), .A3(new_n337), .A4(new_n332), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n321), .B(new_n330), .C1(new_n333), .C2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n327), .A2(KEYINPUT23), .ZN(new_n340));
  OR2_X1    g139(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT23), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n342), .B1(G169gat), .B2(G176gat), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n340), .B(new_n341), .C1(new_n343), .C2(new_n327), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT24), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n321), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n346), .B(new_n347), .C1(G183gat), .C2(G190gat), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n342), .A2(G169gat), .A3(G176gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n326), .A2(KEYINPUT23), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n349), .B1(new_n324), .B2(new_n350), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n344), .B(new_n348), .C1(new_n351), .C2(KEYINPUT64), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n340), .B1(new_n343), .B2(new_n327), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT66), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(G183gat), .B2(G190gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n334), .A2(new_n332), .A3(KEYINPUT66), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n345), .A2(new_n334), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n355), .A2(new_n356), .B1(new_n357), .B2(G190gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n321), .A2(KEYINPUT65), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT65), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(G183gat), .A3(G190gat), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(new_n361), .A3(new_n345), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n353), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT25), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n339), .B(new_n352), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  AND2_X1   g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT29), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n366), .B1(new_n365), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n320), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  OR2_X1    g170(.A1(new_n333), .A2(new_n338), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n330), .A2(new_n321), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n355), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n362), .A2(new_n374), .A3(new_n347), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n351), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n372), .A2(new_n373), .B1(new_n376), .B2(KEYINPUT25), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT29), .B1(new_n377), .B2(new_n352), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n319), .B(new_n367), .C1(new_n378), .C2(new_n366), .ZN(new_n379));
  XNOR2_X1  g178(.A(G8gat), .B(G36gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(KEYINPUT71), .ZN(new_n381));
  XNOR2_X1  g180(.A(G64gat), .B(G92gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n371), .A2(new_n379), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT30), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n379), .ZN(new_n387));
  INV_X1    g186(.A(new_n383), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n371), .A2(new_n379), .A3(KEYINPUT30), .A4(new_n383), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n293), .A2(new_n303), .A3(new_n304), .A4(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(KEYINPUT79), .B(G22gat), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G78gat), .B(G106gat), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT70), .B1(new_n309), .B2(new_n310), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n305), .B1(new_n396), .B2(new_n317), .ZN(new_n397));
  INV_X1    g196(.A(new_n318), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n369), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n253), .B1(new_n399), .B2(new_n271), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n319), .B1(new_n369), .B2(new_n272), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n395), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT31), .B(G50gat), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT29), .B1(new_n316), .B2(new_n318), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n225), .B1(new_n404), .B2(KEYINPUT3), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n272), .A2(new_n369), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n320), .ZN(new_n407));
  INV_X1    g206(.A(new_n395), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n405), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n402), .A2(new_n403), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n403), .B1(new_n402), .B2(new_n409), .ZN(new_n411));
  NAND2_X1  g210(.A1(G228gat), .A2(G233gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NOR3_X1   g212(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n403), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n400), .A2(new_n401), .A3(new_n395), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n408), .B1(new_n405), .B2(new_n407), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n409), .A3(new_n403), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n412), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n394), .B1(new_n414), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n413), .B1(new_n410), .B2(new_n411), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n418), .A2(new_n412), .A3(new_n419), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n393), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n296), .A2(new_n298), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n427), .B(new_n290), .C1(new_n300), .C2(new_n301), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n303), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  OAI211_X1 g228(.A(KEYINPUT6), .B(new_n294), .C1(new_n299), .C2(new_n302), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n384), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n383), .B1(new_n387), .B2(KEYINPUT37), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n434), .B1(KEYINPUT37), .B2(new_n387), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n435), .B(KEYINPUT38), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n392), .B(new_n425), .C1(new_n433), .C2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n365), .A2(new_n260), .ZN(new_n438));
  INV_X1    g237(.A(G227gat), .ZN(new_n439));
  INV_X1    g238(.A(G233gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n376), .A2(KEYINPUT25), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n442), .A2(new_n251), .A3(new_n352), .A4(new_n339), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n438), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT33), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT69), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n444), .A2(KEYINPUT69), .A3(new_n445), .ZN(new_n449));
  XNOR2_X1  g248(.A(G15gat), .B(G43gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(G71gat), .B(G99gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n452), .B1(new_n444), .B2(KEYINPUT32), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n448), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n441), .B1(new_n438), .B2(new_n443), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(KEYINPUT34), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n444), .B(KEYINPUT32), .C1(new_n445), .C2(new_n452), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n454), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n456), .B1(new_n454), .B2(new_n457), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(KEYINPUT36), .ZN(new_n461));
  INV_X1    g260(.A(new_n386), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n462), .B1(new_n429), .B2(new_n430), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT72), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n389), .A2(new_n464), .A3(new_n390), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n464), .B1(new_n389), .B2(new_n390), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n437), .B(new_n461), .C1(new_n425), .C2(new_n468), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n421), .A2(new_n424), .ZN(new_n470));
  INV_X1    g269(.A(new_n460), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n391), .ZN(new_n473));
  XOR2_X1   g272(.A(KEYINPUT80), .B(KEYINPUT35), .Z(new_n474));
  NAND4_X1  g273(.A1(new_n472), .A2(new_n431), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n425), .A2(new_n460), .A3(new_n463), .A4(new_n467), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT81), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT35), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n477), .B1(new_n476), .B2(KEYINPUT35), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n469), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G22gat), .ZN(new_n482));
  INV_X1    g281(.A(G1gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT16), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n485), .B1(G1gat), .B2(new_n482), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(G8gat), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n486), .A2(G8gat), .ZN(new_n488));
  OR2_X1    g287(.A1(G71gat), .A2(G78gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(G71gat), .A2(G78gat), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT9), .ZN(new_n492));
  XNOR2_X1  g291(.A(G57gat), .B(G64gat), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT89), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n491), .B(KEYINPUT89), .C1(new_n492), .C2(new_n493), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT90), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n493), .B(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n490), .B1(new_n489), .B2(new_n492), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT21), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n487), .B(new_n488), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n505), .A2(KEYINPUT91), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(KEYINPUT91), .ZN(new_n507));
  XOR2_X1   g306(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(G155gat), .ZN(new_n509));
  OR3_X1    g308(.A1(new_n506), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n509), .B1(new_n506), .B2(new_n507), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n503), .A2(new_n504), .ZN(new_n514));
  NAND2_X1  g313(.A1(G231gat), .A2(G233gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(new_n234), .ZN(new_n517));
  XNOR2_X1  g316(.A(G183gat), .B(G211gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n516), .B(G127gat), .ZN(new_n520));
  INV_X1    g319(.A(new_n518), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n513), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n513), .B1(new_n519), .B2(new_n522), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G29gat), .A2(G36gat), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NOR3_X1   g327(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G43gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G50gat), .ZN(new_n532));
  INV_X1    g331(.A(G50gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(G43gat), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n530), .A2(KEYINPUT15), .A3(new_n532), .A4(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(new_n534), .A3(KEYINPUT82), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT15), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n536), .B(new_n537), .C1(KEYINPUT82), .C2(new_n532), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n532), .A2(new_n534), .A3(KEYINPUT15), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(new_n526), .A3(new_n539), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n529), .A2(KEYINPUT83), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n529), .A2(KEYINPUT83), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n528), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n535), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT84), .B(KEYINPUT17), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g345(.A(KEYINPUT17), .B(new_n535), .C1(new_n540), .C2(new_n543), .ZN(new_n547));
  NAND2_X1  g346(.A1(G85gat), .A2(G92gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT7), .ZN(new_n549));
  NAND2_X1  g348(.A1(G99gat), .A2(G106gat), .ZN(new_n550));
  INV_X1    g349(.A(G85gat), .ZN(new_n551));
  INV_X1    g350(.A(G92gat), .ZN(new_n552));
  AOI22_X1  g351(.A1(KEYINPUT8), .A2(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G99gat), .B(G106gat), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n554), .B(new_n555), .Z(new_n556));
  NAND3_X1  g355(.A1(new_n546), .A2(new_n547), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n554), .B(new_n555), .ZN(new_n558));
  AND2_X1   g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n544), .A2(new_n558), .B1(KEYINPUT41), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n557), .A2(KEYINPUT93), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT93), .B1(new_n557), .B2(new_n560), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n557), .A2(new_n560), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT93), .ZN(new_n567));
  INV_X1    g366(.A(new_n562), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT92), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n559), .A2(KEYINPUT41), .ZN(new_n572));
  OR3_X1    g371(.A1(new_n565), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n572), .B1(new_n565), .B2(new_n571), .ZN(new_n574));
  XOR2_X1   g373(.A(G134gat), .B(G162gat), .Z(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n573), .A2(new_n574), .ZN(new_n577));
  INV_X1    g376(.A(new_n575), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n496), .A2(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n580), .A2(new_n558), .A3(KEYINPUT10), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n549), .A2(new_n555), .A3(new_n553), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT94), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n558), .B1(new_n503), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n556), .A2(new_n580), .A3(new_n583), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g386(.A(KEYINPUT95), .B(new_n581), .C1(new_n587), .C2(KEYINPUT10), .ZN(new_n588));
  NAND2_X1  g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT95), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT10), .B1(new_n585), .B2(new_n586), .ZN(new_n591));
  INV_X1    g390(.A(new_n581), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n588), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G120gat), .B(G148gat), .Z(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT96), .ZN(new_n596));
  XNOR2_X1  g395(.A(G176gat), .B(G204gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n596), .B(new_n597), .Z(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n589), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n599), .B1(new_n587), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n594), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n600), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT97), .B1(new_n605), .B2(new_n599), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT97), .ZN(new_n607));
  AOI211_X1 g406(.A(new_n607), .B(new_n598), .C1(new_n603), .C2(new_n604), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n602), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n525), .A2(new_n576), .A3(new_n579), .A4(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G229gat), .A2(G233gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n612), .B(KEYINPUT13), .Z(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n488), .A2(new_n487), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n615), .A2(new_n544), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n544), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(KEYINPUT85), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT85), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n488), .A2(new_n620), .A3(new_n487), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n619), .A2(new_n546), .A3(new_n547), .A4(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT18), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n623), .B1(G229gat), .B2(G233gat), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n617), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT86), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n618), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G113gat), .B(G141gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G197gat), .ZN(new_n629));
  XOR2_X1   g428(.A(KEYINPUT11), .B(G169gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n631), .B(KEYINPUT12), .Z(new_n632));
  NAND3_X1  g431(.A1(new_n622), .A2(new_n617), .A3(new_n612), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n632), .B1(new_n633), .B2(new_n623), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n622), .A2(KEYINPUT86), .A3(new_n617), .A4(new_n624), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n627), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT88), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n627), .A2(new_n634), .A3(KEYINPUT88), .A4(new_n635), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n627), .A2(KEYINPUT87), .A3(new_n635), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT87), .B1(new_n627), .B2(new_n635), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n633), .A2(new_n623), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n632), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n611), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n481), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(new_n431), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(new_n483), .ZN(G1324gat));
  NAND3_X1  g450(.A1(new_n481), .A2(new_n391), .A3(new_n648), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT16), .B(G8gat), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n654), .A2(KEYINPUT42), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(KEYINPUT42), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n652), .A2(G8gat), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(G1325gat));
  OAI21_X1  g457(.A(G15gat), .B1(new_n649), .B2(new_n461), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n471), .A2(G15gat), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n659), .B1(new_n649), .B2(new_n660), .ZN(G1326gat));
  NOR2_X1   g460(.A1(new_n649), .A2(new_n425), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT43), .B(G22gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1327gat));
  NOR3_X1   g463(.A1(new_n647), .A2(new_n525), .A3(new_n609), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT98), .Z(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT99), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n480), .A2(new_n668), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n475), .B(KEYINPUT99), .C1(new_n478), .C2(new_n479), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n469), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n579), .A2(new_n576), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n673), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n678), .B1(new_n469), .B2(new_n480), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(new_n674), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n667), .B1(new_n677), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(G29gat), .B1(new_n683), .B2(new_n431), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n679), .A2(new_n665), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n685), .A2(G29gat), .A3(new_n431), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT45), .Z(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(new_n687), .ZN(G1328gat));
  OAI21_X1  g487(.A(G36gat), .B1(new_n683), .B2(new_n473), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n473), .A2(G36gat), .ZN(new_n690));
  OAI21_X1  g489(.A(KEYINPUT46), .B1(new_n685), .B2(new_n690), .ZN(new_n691));
  OR3_X1    g490(.A1(new_n685), .A2(KEYINPUT46), .A3(new_n690), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(KEYINPUT100), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT100), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n689), .A2(new_n695), .A3(new_n691), .A4(new_n692), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(G1329gat));
  OAI21_X1  g496(.A(new_n531), .B1(new_n685), .B2(new_n471), .ZN(new_n698));
  INV_X1    g497(.A(new_n461), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(G43gat), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n683), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g501(.A(new_n675), .B1(new_n671), .B2(new_n469), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n470), .B(new_n666), .C1(new_n703), .C2(new_n680), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(G50gat), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n685), .A2(G50gat), .A3(new_n425), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT102), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n705), .A2(KEYINPUT101), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT48), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n713), .B1(new_n704), .B2(G50gat), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(KEYINPUT102), .A3(KEYINPUT48), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n708), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n710), .A2(new_n709), .A3(new_n711), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n706), .A2(new_n707), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT102), .B1(new_n714), .B2(KEYINPUT48), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n716), .A2(new_n720), .ZN(G1331gat));
  INV_X1    g520(.A(new_n525), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(new_n673), .ZN(new_n723));
  AND4_X1   g522(.A1(new_n647), .A2(new_n672), .A3(new_n723), .A4(new_n609), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n432), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n391), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT49), .B(G64gat), .Z(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n727), .B2(new_n729), .ZN(G1333gat));
  NAND2_X1  g529(.A1(new_n724), .A2(new_n699), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n471), .A2(G71gat), .ZN(new_n732));
  AOI22_X1  g531(.A1(new_n731), .A2(G71gat), .B1(new_n724), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g533(.A1(new_n724), .A2(new_n470), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g535(.A1(new_n722), .A2(new_n647), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n610), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n703), .B2(new_n680), .ZN(new_n739));
  OAI21_X1  g538(.A(G85gat), .B1(new_n739), .B2(new_n431), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n737), .A2(new_n678), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n672), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT51), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n672), .A2(KEYINPUT51), .A3(new_n741), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n432), .A2(new_n609), .A3(new_n551), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n740), .B1(new_n747), .B2(new_n748), .ZN(G1336gat));
  NAND3_X1  g548(.A1(new_n609), .A2(new_n552), .A3(new_n391), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT104), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n751), .B1(new_n744), .B2(new_n745), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(KEYINPUT52), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n391), .B(new_n738), .C1(new_n703), .C2(new_n680), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G92gat), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n753), .A2(KEYINPUT105), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT105), .B1(new_n753), .B2(new_n755), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n754), .A2(KEYINPUT103), .A3(G92gat), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT103), .B1(new_n754), .B2(G92gat), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n758), .A2(new_n759), .A3(new_n752), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761));
  OAI22_X1  g560(.A1(new_n756), .A2(new_n757), .B1(new_n760), .B2(new_n761), .ZN(G1337gat));
  OAI21_X1  g561(.A(KEYINPUT106), .B1(new_n739), .B2(new_n461), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G99gat), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n739), .A2(KEYINPUT106), .A3(new_n461), .ZN(new_n765));
  OR3_X1    g564(.A1(new_n610), .A2(new_n471), .A3(G99gat), .ZN(new_n766));
  OAI22_X1  g565(.A1(new_n764), .A2(new_n765), .B1(new_n747), .B2(new_n766), .ZN(G1338gat));
  NOR3_X1   g566(.A1(new_n610), .A2(G106gat), .A3(new_n425), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n746), .A2(new_n768), .ZN(new_n769));
  XOR2_X1   g568(.A(KEYINPUT107), .B(G106gat), .Z(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n739), .B2(new_n425), .ZN(new_n771));
  XNOR2_X1  g570(.A(KEYINPUT108), .B(KEYINPUT53), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n769), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n769), .A2(KEYINPUT109), .A3(new_n771), .A4(new_n772), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n769), .A2(new_n771), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT53), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(G1339gat));
  NAND3_X1  g578(.A1(new_n646), .A2(new_n227), .A3(new_n229), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT114), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n431), .A2(new_n391), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n611), .A2(new_n646), .ZN(new_n783));
  INV_X1    g582(.A(new_n602), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n591), .A2(new_n592), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n786), .B2(new_n600), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n594), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n785), .B(new_n589), .C1(new_n591), .C2(new_n592), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n789), .A2(KEYINPUT110), .A3(new_n599), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT110), .B1(new_n789), .B2(new_n599), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT55), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n788), .B(new_n794), .C1(new_n790), .C2(new_n791), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n784), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n612), .B1(new_n622), .B2(new_n617), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n797), .A2(KEYINPUT111), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n616), .A2(new_n617), .A3(new_n614), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n799), .B1(new_n797), .B2(KEYINPUT111), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n631), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n796), .A2(new_n673), .A3(new_n640), .A4(new_n801), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n640), .A2(new_n609), .A3(new_n801), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n796), .B2(new_n646), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n804), .B2(new_n673), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n783), .B1(new_n805), .B2(new_n722), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(KEYINPUT112), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n808));
  AOI211_X1 g607(.A(new_n808), .B(new_n783), .C1(new_n805), .C2(new_n722), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n472), .B(new_n782), .C1(new_n807), .C2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n810), .A2(KEYINPUT113), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n810), .A2(KEYINPUT113), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n781), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(G113gat), .B1(new_n810), .B2(new_n647), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(G1340gat));
  OAI211_X1 g614(.A(new_n231), .B(new_n609), .C1(new_n811), .C2(new_n812), .ZN(new_n816));
  OAI21_X1  g615(.A(G120gat), .B1(new_n810), .B2(new_n610), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n816), .A2(KEYINPUT115), .A3(new_n817), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(G1341gat));
  NOR2_X1   g621(.A1(new_n810), .A2(new_n722), .ZN(new_n823));
  XNOR2_X1  g622(.A(KEYINPUT116), .B(G127gat), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n823), .B(new_n824), .ZN(G1342gat));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n678), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n255), .A2(new_n245), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n826), .A2(KEYINPUT56), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT56), .B1(new_n826), .B2(new_n828), .ZN(new_n830));
  OAI21_X1  g629(.A(G134gat), .B1(new_n810), .B2(new_n678), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(G1343gat));
  INV_X1    g631(.A(KEYINPUT58), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n805), .A2(new_n722), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n808), .B1(new_n834), .B2(new_n783), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n806), .A2(KEYINPUT112), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n837), .A2(KEYINPUT118), .A3(new_n432), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n432), .B1(new_n807), .B2(new_n809), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n699), .A2(new_n425), .A3(new_n391), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n647), .A2(G141gat), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n838), .A2(new_n841), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n833), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT57), .B1(new_n806), .B2(new_n425), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n847), .A2(new_n461), .A3(new_n782), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n849), .B(new_n470), .C1(new_n807), .C2(new_n809), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G141gat), .B1(new_n851), .B2(new_n647), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n844), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n846), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n852), .B(new_n844), .C1(new_n845), .C2(new_n833), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(G1344gat));
  NOR2_X1   g655(.A1(new_n610), .A2(G148gat), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n838), .A2(new_n841), .A3(new_n842), .A4(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n851), .A2(new_n610), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n859), .A2(KEYINPUT59), .A3(new_n207), .ZN(new_n860));
  XOR2_X1   g659(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n861));
  OAI211_X1 g660(.A(KEYINPUT57), .B(new_n470), .C1(new_n807), .C2(new_n809), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n849), .B1(new_n806), .B2(new_n425), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n864), .A2(new_n461), .A3(new_n609), .A4(new_n782), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n861), .B1(new_n865), .B2(G148gat), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n858), .B1(new_n860), .B2(new_n866), .ZN(G1345gat));
  OAI21_X1  g666(.A(G155gat), .B1(new_n851), .B2(new_n722), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n722), .A2(G155gat), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n838), .A2(new_n841), .A3(new_n842), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(G1346gat));
  OAI21_X1  g670(.A(G162gat), .B1(new_n851), .B2(new_n678), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n678), .A2(G162gat), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n838), .A2(new_n841), .A3(new_n842), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(G1347gat));
  INV_X1    g674(.A(new_n472), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n876), .B1(new_n835), .B2(new_n836), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n432), .A2(new_n473), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n647), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(new_n322), .ZN(G1348gat));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n610), .B1(new_n882), .B2(new_n323), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n877), .A2(new_n878), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n882), .A2(new_n323), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n884), .B(new_n885), .ZN(G1349gat));
  OAI21_X1  g685(.A(new_n334), .B1(new_n879), .B2(new_n722), .ZN(new_n887));
  INV_X1    g686(.A(new_n331), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n877), .A2(new_n888), .A3(new_n525), .A4(new_n878), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT60), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n890), .B(new_n891), .ZN(G1350gat));
  OAI21_X1  g691(.A(G190gat), .B1(new_n879), .B2(new_n678), .ZN(new_n893));
  NOR2_X1   g692(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n877), .A2(new_n332), .A3(new_n673), .A4(new_n878), .ZN(new_n896));
  XNOR2_X1  g695(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n895), .B(new_n896), .C1(new_n893), .C2(new_n897), .ZN(G1351gat));
  NAND3_X1  g697(.A1(new_n461), .A2(new_n470), .A3(new_n391), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n899), .A2(new_n900), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n901), .A2(new_n902), .A3(new_n432), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n837), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT123), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n837), .A2(new_n906), .A3(new_n903), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n908), .A2(new_n647), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(G197gat), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n864), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n862), .A2(KEYINPUT124), .A3(new_n863), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n461), .A2(new_n878), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT125), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n912), .A2(new_n913), .A3(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(G197gat), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n917), .A2(new_n918), .A3(new_n647), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n910), .A2(new_n919), .ZN(G1352gat));
  NOR3_X1   g719(.A1(new_n904), .A2(G204gat), .A3(new_n610), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT62), .ZN(new_n922));
  OAI21_X1  g721(.A(G204gat), .B1(new_n917), .B2(new_n610), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1353gat));
  AND2_X1   g723(.A1(new_n862), .A2(new_n863), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n916), .A2(new_n525), .ZN(new_n926));
  OAI21_X1  g725(.A(G211gat), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  XOR2_X1   g726(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n722), .A2(G211gat), .ZN(new_n930));
  OR2_X1    g729(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n931));
  OAI221_X1 g730(.A(new_n929), .B1(new_n908), .B2(new_n930), .C1(new_n927), .C2(new_n931), .ZN(G1354gat));
  NAND2_X1  g731(.A1(new_n673), .A2(G218gat), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n933), .B1(new_n917), .B2(KEYINPUT127), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n912), .A2(new_n935), .A3(new_n913), .A4(new_n916), .ZN(new_n936));
  INV_X1    g735(.A(G218gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n905), .A2(new_n673), .A3(new_n907), .ZN(new_n938));
  AOI22_X1  g737(.A1(new_n934), .A2(new_n936), .B1(new_n937), .B2(new_n938), .ZN(G1355gat));
endmodule


