//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n604, new_n605, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT66), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  NAND2_X1  g033(.A1(new_n453), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(new_n456), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n464), .A2(G137), .A3(new_n463), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  OR2_X1    g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n475));
  OR2_X1    g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n463), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n475), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(G136), .B2(new_n482), .ZN(G162));
  AND2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  OAI211_X1 g060(.A(G126), .B(G2105), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n487), .A2(new_n489), .A3(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n463), .C1(new_n484), .C2(new_n485), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n464), .A2(new_n494), .A3(G138), .A4(new_n463), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(G164));
  NAND2_X1  g071(.A1(KEYINPUT69), .A2(G651), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT68), .A2(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT6), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT68), .B1(KEYINPUT69), .B2(G651), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n500), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G50), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT70), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n497), .A2(new_n498), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT6), .A3(new_n501), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n508), .B1(new_n510), .B2(new_n500), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(new_n512), .A3(G50), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n517), .B1(new_n510), .B2(new_n500), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G62), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n518), .A2(G88), .B1(new_n521), .B2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n514), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND2_X1  g099(.A1(new_n511), .A2(G51), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n518), .A2(G89), .ZN(new_n526));
  INV_X1    g101(.A(new_n517), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n527), .A2(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n525), .A2(new_n526), .A3(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  AOI22_X1  g109(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G651), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n511), .A2(G52), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n518), .A2(G90), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  AOI22_X1  g116(.A1(G43), .A2(new_n511), .B1(new_n518), .B2(G81), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n517), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT71), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n547));
  OAI211_X1 g122(.A(new_n547), .B(new_n543), .C1(new_n517), .C2(new_n544), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n546), .A2(G651), .A3(new_n548), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n542), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT9), .B1(new_n505), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n511), .A2(new_n558), .A3(G53), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OR2_X1    g136(.A1(KEYINPUT5), .A2(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(KEYINPUT5), .A2(G543), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AND2_X1   g139(.A1(G78), .A2(G543), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n518), .A2(G91), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n560), .A2(new_n566), .A3(new_n567), .ZN(G299));
  NAND2_X1  g143(.A1(new_n511), .A2(G49), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n518), .A2(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  NAND3_X1  g147(.A1(new_n504), .A2(G48), .A3(G543), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n562), .B2(new_n563), .ZN(new_n575));
  AND2_X1   g150(.A1(G73), .A2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n504), .A2(new_n527), .A3(G86), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G305));
  NAND2_X1  g155(.A1(new_n511), .A2(G47), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n504), .A2(new_n527), .ZN(new_n582));
  XNOR2_X1  g157(.A(KEYINPUT72), .B(G85), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n527), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  OAI221_X1 g159(.A(new_n581), .B1(new_n582), .B2(new_n583), .C1(new_n536), .C2(new_n584), .ZN(G290));
  INV_X1    g160(.A(KEYINPUT73), .ZN(new_n586));
  INV_X1    g161(.A(G79), .ZN(new_n587));
  INV_X1    g162(.A(G66), .ZN(new_n588));
  OAI221_X1 g163(.A(new_n586), .B1(new_n587), .B2(new_n508), .C1(new_n517), .C2(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n588), .B1(new_n562), .B2(new_n563), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n587), .A2(new_n508), .ZN(new_n591));
  OAI21_X1  g166(.A(KEYINPUT73), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n589), .A2(G651), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n511), .A2(G54), .ZN(new_n594));
  AOI21_X1  g169(.A(KEYINPUT10), .B1(new_n518), .B2(G92), .ZN(new_n595));
  AND4_X1   g170(.A1(KEYINPUT10), .A2(new_n504), .A3(new_n527), .A4(G92), .ZN(new_n596));
  OAI211_X1 g171(.A(new_n593), .B(new_n594), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(G171), .B2(new_n598), .ZN(G321));
  XOR2_X1   g175(.A(G321), .B(KEYINPUT74), .Z(G284));
  NAND2_X1  g176(.A1(G286), .A2(G868), .ZN(new_n602));
  INV_X1    g177(.A(G91), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n566), .B1(new_n582), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n604), .B1(new_n557), .B2(new_n559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n602), .B1(new_n605), .B2(G868), .ZN(G297));
  OAI21_X1  g181(.A(new_n602), .B1(new_n605), .B2(G868), .ZN(G280));
  INV_X1    g182(.A(new_n597), .ZN(new_n608));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n542), .A2(new_n549), .ZN(new_n611));
  OR3_X1    g186(.A1(new_n597), .A2(KEYINPUT75), .A3(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(KEYINPUT75), .B1(new_n597), .B2(G559), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  MUX2_X1   g189(.A(new_n611), .B(new_n614), .S(G868), .Z(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g191(.A1(new_n464), .A2(new_n470), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT12), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  XOR2_X1   g194(.A(KEYINPUT76), .B(G2100), .Z(new_n620));
  OR2_X1    g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n482), .A2(G135), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n478), .A2(G123), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n463), .A2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NAND3_X1  g203(.A1(new_n621), .A2(new_n622), .A3(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT77), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2430), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2443), .B(G2446), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G1341), .B(G1348), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT78), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(G14), .A3(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(G401));
  INV_X1    g222(.A(KEYINPUT18), .ZN(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n648), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2100), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n651), .B2(KEYINPUT18), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2096), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(G227));
  XNOR2_X1  g234(.A(G1961), .B(G1966), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT79), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1956), .B(G2474), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT20), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n661), .A2(new_n662), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n669), .A2(new_n665), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT80), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n663), .A2(new_n669), .A3(new_n665), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n668), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n679), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(G229));
  NAND2_X1  g257(.A1(G290), .A2(G16), .ZN(new_n683));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G24), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT83), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(G1986), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n478), .A2(G119), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT81), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n482), .A2(G131), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n463), .A2(G107), .ZN(new_n692));
  OAI21_X1  g267(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n690), .B(new_n691), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G25), .B(new_n694), .S(G29), .Z(new_n695));
  XOR2_X1   g270(.A(KEYINPUT35), .B(G1991), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT82), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n688), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n698), .B2(new_n697), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n684), .A2(G22), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G166), .B2(new_n684), .ZN(new_n702));
  INV_X1    g277(.A(G1971), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  MUX2_X1   g279(.A(G6), .B(G305), .S(G16), .Z(new_n705));
  XOR2_X1   g280(.A(KEYINPUT32), .B(G1981), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT84), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n705), .B(new_n707), .ZN(new_n708));
  MUX2_X1   g283(.A(G23), .B(G288), .S(G16), .Z(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT33), .B(G1976), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n704), .A2(new_n708), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(KEYINPUT34), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(KEYINPUT34), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n700), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT85), .ZN(new_n716));
  OR3_X1    g291(.A1(new_n715), .A2(new_n716), .A3(KEYINPUT36), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT85), .B(KEYINPUT36), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT30), .B(G28), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  OR2_X1    g296(.A1(KEYINPUT31), .A2(G11), .ZN(new_n722));
  NAND2_X1  g297(.A1(KEYINPUT31), .A2(G11), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n720), .A2(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n627), .B2(new_n721), .ZN(new_n725));
  NOR2_X1   g300(.A1(G171), .A2(new_n684), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G5), .B2(new_n684), .ZN(new_n727));
  INV_X1    g302(.A(G1961), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n684), .A2(G21), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G168), .B2(new_n684), .ZN(new_n730));
  OAI22_X1  g305(.A1(new_n727), .A2(new_n728), .B1(G1966), .B2(new_n730), .ZN(new_n731));
  AOI211_X1 g306(.A(new_n725), .B(new_n731), .C1(G1966), .C2(new_n730), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n732), .A2(KEYINPUT92), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(KEYINPUT92), .ZN(new_n734));
  NOR2_X1   g309(.A1(G29), .A2(G35), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G162), .B2(G29), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G2090), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT94), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n721), .A2(G32), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n470), .A2(G105), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT91), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n482), .A2(G141), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n478), .A2(G129), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(KEYINPUT26), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(KEYINPUT26), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n747), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n746), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n742), .B1(new_n752), .B2(new_n721), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT27), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1996), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n721), .A2(G27), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G164), .B2(new_n721), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G2078), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n727), .B2(new_n728), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n741), .A2(new_n755), .A3(new_n759), .ZN(new_n760));
  NOR3_X1   g335(.A1(new_n733), .A2(new_n734), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n721), .A2(G33), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT88), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT25), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n464), .A2(G127), .ZN(new_n766));
  INV_X1    g341(.A(G115), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(new_n469), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n768), .A2(G2105), .B1(G139), .B2(new_n482), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT89), .Z(new_n771));
  OAI21_X1  g346(.A(new_n762), .B1(new_n771), .B2(new_n721), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(G2072), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n684), .A2(G20), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT23), .Z(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G299), .B2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1956), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT24), .ZN(new_n778));
  INV_X1    g353(.A(G34), .ZN(new_n779));
  AOI21_X1  g354(.A(G29), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n778), .B2(new_n779), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G160), .B2(new_n721), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT90), .Z(new_n783));
  OAI22_X1  g358(.A1(new_n738), .A2(new_n739), .B1(new_n783), .B2(G2084), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G2084), .B2(new_n783), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n773), .A2(new_n777), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n684), .A2(G4), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n608), .B2(new_n684), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1348), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n721), .A2(G26), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT28), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n482), .A2(G140), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n478), .A2(G128), .ZN(new_n793));
  OR2_X1    g368(.A1(G104), .A2(G2105), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n794), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n792), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(G29), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n797), .A2(KEYINPUT86), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(KEYINPUT86), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n791), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G2067), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n684), .A2(G19), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n550), .B2(new_n684), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1341), .ZN(new_n804));
  OR3_X1    g379(.A1(new_n789), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n805), .A2(KEYINPUT87), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n805), .A2(KEYINPUT87), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n786), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n717), .A2(new_n719), .A3(new_n761), .A4(new_n808), .ZN(G150));
  INV_X1    g384(.A(G150), .ZN(G311));
  NAND2_X1  g385(.A1(G80), .A2(G543), .ZN(new_n811));
  INV_X1    g386(.A(G67), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n517), .B2(new_n812), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n518), .A2(G93), .B1(new_n813), .B2(G651), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n511), .A2(G55), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G860), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT96), .B(KEYINPUT37), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n608), .A2(G559), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT95), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT38), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n611), .A2(new_n816), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n542), .A2(new_n549), .A3(new_n815), .A4(new_n814), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n822), .B(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n826), .A2(KEYINPUT39), .ZN(new_n827));
  INV_X1    g402(.A(G860), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n826), .B2(KEYINPUT39), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n819), .B1(new_n827), .B2(new_n829), .ZN(G145));
  NAND2_X1  g405(.A1(new_n493), .A2(new_n495), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT97), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n491), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n486), .A2(KEYINPUT97), .A3(new_n490), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n831), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n796), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n482), .A2(G142), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n478), .A2(G130), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n463), .A2(G118), .ZN(new_n839));
  OAI21_X1  g414(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n837), .B(new_n838), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n836), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n771), .A2(new_n752), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n770), .B(KEYINPUT89), .ZN(new_n845));
  INV_X1    g420(.A(new_n752), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n694), .B(new_n618), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n844), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n849), .B1(new_n844), .B2(new_n847), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n843), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(G160), .B(new_n627), .Z(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(G162), .Z(new_n855));
  NAND2_X1  g430(.A1(new_n844), .A2(new_n847), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n848), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n857), .A2(new_n842), .A3(new_n850), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n853), .A2(new_n855), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G37), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n855), .B1(new_n853), .B2(new_n858), .ZN(new_n862));
  OAI21_X1  g437(.A(KEYINPUT98), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n853), .A2(new_n858), .ZN(new_n864));
  INV_X1    g439(.A(new_n855), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT98), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n866), .A2(new_n859), .A3(new_n867), .A4(new_n860), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT40), .ZN(G395));
  AND2_X1   g445(.A1(new_n614), .A2(new_n825), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n614), .A2(new_n825), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n597), .A2(new_n605), .A3(KEYINPUT99), .ZN(new_n874));
  AOI21_X1  g449(.A(KEYINPUT99), .B1(new_n597), .B2(new_n605), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n597), .A2(new_n605), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n881));
  NOR4_X1   g456(.A1(new_n874), .A2(new_n875), .A3(new_n877), .A4(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n875), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT100), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n597), .A2(new_n605), .A3(KEYINPUT99), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(KEYINPUT100), .B1(new_n874), .B2(new_n875), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n886), .A2(new_n887), .A3(new_n878), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n882), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n880), .B1(new_n873), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT102), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(new_n892), .A3(KEYINPUT42), .ZN(new_n893));
  XNOR2_X1  g468(.A(G303), .B(G290), .ZN(new_n894));
  XOR2_X1   g469(.A(G305), .B(G288), .Z(new_n895));
  XNOR2_X1  g470(.A(new_n894), .B(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n896), .B1(KEYINPUT102), .B2(new_n897), .ZN(new_n898));
  OAI221_X1 g473(.A(new_n880), .B1(KEYINPUT102), .B2(new_n897), .C1(new_n873), .C2(new_n890), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n893), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n898), .B1(new_n893), .B2(new_n899), .ZN(new_n901));
  OAI21_X1  g476(.A(G868), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n816), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n902), .B1(G868), .B2(new_n903), .ZN(G295));
  OAI21_X1  g479(.A(new_n902), .B1(G868), .B2(new_n903), .ZN(G331));
  NAND3_X1  g480(.A1(new_n823), .A2(G301), .A3(new_n824), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(G301), .B1(new_n823), .B2(new_n824), .ZN(new_n908));
  OAI21_X1  g483(.A(G286), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n908), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(G168), .A3(new_n906), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n879), .ZN(new_n913));
  INV_X1    g488(.A(new_n896), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n913), .B(new_n914), .C1(new_n890), .C2(new_n912), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n913), .B1(new_n890), .B2(new_n912), .ZN(new_n917));
  AOI21_X1  g492(.A(G37), .B1(new_n917), .B2(new_n896), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n912), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n877), .B1(new_n876), .B2(new_n884), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT41), .B1(new_n922), .B2(new_n887), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n921), .B1(new_n923), .B2(new_n882), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n914), .B1(new_n924), .B2(new_n913), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT103), .B1(new_n925), .B2(G37), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT43), .B1(new_n920), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n913), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n879), .A2(new_n881), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT104), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n879), .A2(new_n931), .A3(new_n881), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n930), .B(new_n932), .C1(new_n889), .C2(new_n888), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n928), .B1(new_n933), .B2(new_n921), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n860), .B(new_n915), .C1(new_n934), .C2(new_n914), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT44), .B1(new_n927), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n936), .B1(new_n920), .B2(new_n926), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n935), .A2(KEYINPUT43), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n938), .A2(new_n942), .ZN(G397));
  INV_X1    g518(.A(G1384), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT45), .B1(new_n835), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(KEYINPUT105), .B(G40), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(G160), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n796), .B(G2067), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n951), .B(KEYINPUT108), .Z(new_n952));
  INV_X1    g527(.A(G1996), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n752), .B(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n950), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT109), .ZN(new_n956));
  INV_X1    g531(.A(new_n950), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n694), .B(new_n696), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(G290), .A2(G1986), .ZN(new_n960));
  XOR2_X1   g535(.A(new_n960), .B(KEYINPUT106), .Z(new_n961));
  NAND2_X1  g536(.A1(G290), .A2(G1986), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT107), .ZN(new_n963));
  OR2_X1    g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n959), .B1(new_n950), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT54), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n835), .A2(KEYINPUT45), .A3(new_n944), .ZN(new_n967));
  INV_X1    g542(.A(G2078), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n467), .A2(new_n472), .A3(new_n947), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(G164), .B2(G1384), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n967), .A2(new_n968), .A3(new_n969), .A4(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT124), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT124), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n972), .A2(new_n976), .A3(new_n973), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT50), .B1(new_n835), .B2(new_n944), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n980));
  NOR3_X1   g555(.A1(G164), .A2(new_n980), .A3(G1384), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n969), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n728), .ZN(new_n983));
  INV_X1    g558(.A(new_n491), .ZN(new_n984));
  AOI21_X1  g559(.A(G1384), .B1(new_n831), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT45), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n968), .A2(KEYINPUT53), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n946), .A2(new_n969), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(G301), .B1(new_n978), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT125), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n472), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n465), .A2(new_n466), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(G2105), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n468), .A2(KEYINPUT125), .A3(new_n471), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n987), .A2(G40), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n992), .A2(new_n994), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n835), .A2(new_n944), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n997), .B1(new_n998), .B2(new_n970), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n982), .A2(new_n728), .B1(new_n999), .B2(new_n967), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n972), .A2(new_n976), .A3(new_n973), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n976), .B1(new_n972), .B2(new_n973), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1000), .B(G301), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n966), .B1(new_n990), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1966), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n986), .A2(new_n969), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1006), .B1(new_n1007), .B2(new_n945), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n949), .A2(G2084), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n979), .B2(new_n981), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1008), .A2(G168), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G8), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1012), .A2(KEYINPUT122), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT51), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1016), .A2(G8), .A3(G286), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1011), .A2(new_n1018), .A3(new_n1013), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1015), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n983), .A2(G301), .A3(new_n988), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n966), .B1(new_n1021), .B2(new_n978), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1000), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(G171), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1005), .A2(new_n1020), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n998), .A2(KEYINPUT50), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n1028), .A3(new_n969), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n980), .B1(new_n835), .B2(new_n944), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT115), .B1(new_n1030), .B2(new_n949), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n985), .A2(new_n980), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1029), .A2(new_n1031), .A3(new_n739), .A4(new_n1032), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n835), .A2(KEYINPUT45), .A3(new_n944), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n969), .B1(new_n985), .B2(KEYINPUT45), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n703), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1012), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(G166), .B2(new_n1012), .ZN(new_n1039));
  NAND3_X1  g614(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n1037), .A2(new_n1041), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n739), .B(new_n969), .C1(new_n979), .C2(new_n981), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1036), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT110), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT110), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1036), .A2(new_n1043), .A3(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1045), .A2(G8), .A3(new_n1041), .A4(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n969), .A2(new_n944), .A3(new_n835), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G8), .ZN(new_n1050));
  INV_X1    g625(.A(G1981), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n578), .A2(KEYINPUT111), .A3(new_n1051), .A4(new_n579), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n579), .A2(new_n573), .A3(new_n577), .A4(new_n1051), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT111), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT112), .B(G86), .Z(new_n1057));
  OAI211_X1 g632(.A(new_n573), .B(new_n577), .C1(new_n582), .C2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(G1981), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n1061));
  AOI21_X1  g636(.A(new_n1050), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1052), .A2(new_n1055), .B1(new_n1058), .B2(G1981), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1063), .A2(KEYINPUT114), .A3(KEYINPUT49), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT114), .B1(new_n1063), .B2(KEYINPUT49), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1062), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n1067));
  INV_X1    g642(.A(G1976), .ZN(new_n1068));
  NOR2_X1   g643(.A1(G288), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT52), .B1(new_n1050), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1069), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT52), .B1(G288), .B2(new_n1068), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1071), .A2(new_n1072), .A3(G8), .A4(new_n1049), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1066), .A2(new_n1067), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1067), .B1(new_n1066), .B2(new_n1074), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1042), .B(new_n1048), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT126), .B1(new_n1026), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1048), .B1(new_n1041), .B2(new_n1037), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1066), .A2(new_n1074), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT116), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1066), .A2(new_n1067), .A3(new_n1074), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT126), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1019), .A2(new_n1017), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1086), .A2(new_n1015), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1083), .A2(new_n1084), .A3(new_n1005), .A4(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1029), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1089));
  INV_X1    g664(.A(G1956), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT56), .B(G2072), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1095), .B1(G299), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n605), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n1100));
  NAND3_X1  g675(.A1(G299), .A2(new_n1100), .A3(new_n1096), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT119), .B1(new_n605), .B2(KEYINPUT57), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1091), .A2(new_n1094), .A3(new_n1104), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n949), .B1(new_n998), .B2(KEYINPUT50), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1107), .A2(new_n1028), .B1(new_n980), .B2(new_n985), .ZN(new_n1108));
  AOI21_X1  g683(.A(G1956), .B1(new_n1108), .B2(new_n1031), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1094), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1106), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n998), .A2(new_n980), .ZN(new_n1113));
  INV_X1    g688(.A(new_n981), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n949), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI22_X1  g690(.A1(new_n1115), .A2(G1348), .B1(G2067), .B2(new_n1049), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1116), .A2(new_n608), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1105), .B1(new_n1112), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1111), .A2(KEYINPUT61), .A3(new_n1105), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT60), .ZN(new_n1120));
  OR3_X1    g695(.A1(new_n1116), .A2(new_n1120), .A3(new_n608), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n597), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n1120), .B2(new_n1116), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n1124));
  NAND2_X1  g699(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n967), .A2(new_n953), .A3(new_n969), .A4(new_n971), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT58), .B(G1341), .Z(new_n1127));
  NAND2_X1  g702(.A1(new_n1049), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n611), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  MUX2_X1   g704(.A(new_n1124), .B(new_n1125), .S(new_n1129), .Z(new_n1130));
  NAND4_X1  g705(.A1(new_n1119), .A2(new_n1121), .A3(new_n1123), .A4(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT61), .B1(new_n1111), .B2(new_n1105), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1118), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1078), .A2(new_n1088), .A3(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(G288), .A2(G1976), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1066), .A2(new_n1135), .B1(new_n1055), .B2(new_n1052), .ZN(new_n1136));
  OAI22_X1  g711(.A1(new_n1136), .A2(new_n1050), .B1(new_n1080), .B2(new_n1048), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1018), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1138));
  OAI211_X1 g713(.A(KEYINPUT127), .B(KEYINPUT62), .C1(new_n1085), .C2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n990), .B1(new_n1020), .B2(KEYINPUT62), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT127), .B1(new_n1020), .B2(KEYINPUT62), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1077), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1137), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1134), .A2(new_n1145), .ZN(new_n1146));
  AOI211_X1 g721(.A(new_n1012), .B(G286), .C1(new_n1008), .C2(new_n1010), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1048), .A2(KEYINPUT63), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1080), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1045), .A2(G8), .A3(new_n1047), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1150), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1149), .A2(new_n1151), .A3(KEYINPUT118), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1148), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1157), .A2(new_n1048), .A3(new_n1042), .A4(new_n1147), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT117), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT63), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1083), .A2(KEYINPUT117), .A3(new_n1147), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1156), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n965), .B1(new_n1146), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n961), .A2(new_n950), .ZN(new_n1164));
  XOR2_X1   g739(.A(new_n1164), .B(KEYINPUT48), .Z(new_n1165));
  NOR2_X1   g740(.A1(new_n959), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n696), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n694), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n956), .A2(new_n1168), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n796), .A2(G2067), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n957), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OR2_X1    g746(.A1(new_n952), .A2(new_n846), .ZN(new_n1172));
  OR3_X1    g747(.A1(new_n957), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT46), .B1(new_n957), .B2(G1996), .ZN(new_n1174));
  AOI22_X1  g749(.A1(new_n1172), .A2(new_n950), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT47), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1166), .A2(new_n1171), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1163), .A2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g753(.A1(new_n461), .A2(G227), .ZN(new_n1180));
  NAND2_X1  g754(.A1(new_n646), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g755(.A(new_n1181), .B1(new_n680), .B2(new_n681), .ZN(new_n1182));
  OAI211_X1 g756(.A(new_n869), .B(new_n1182), .C1(new_n940), .C2(new_n941), .ZN(G225));
  INV_X1    g757(.A(G225), .ZN(G308));
endmodule


