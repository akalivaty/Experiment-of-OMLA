

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593;

  XOR2_X1 U326 ( .A(KEYINPUT41), .B(n582), .Z(n558) );
  XNOR2_X1 U327 ( .A(n330), .B(n329), .ZN(n396) );
  NOR2_X2 U328 ( .A1(n479), .A2(n458), .ZN(n549) );
  NOR2_X2 U329 ( .A1(n479), .A2(n467), .ZN(n570) );
  NOR2_X1 U330 ( .A1(n398), .A2(n582), .ZN(n399) );
  XNOR2_X1 U331 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n403) );
  XNOR2_X1 U332 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U333 ( .A(G36GAT), .B(G190GAT), .Z(n434) );
  XNOR2_X1 U334 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U335 ( .A(n368), .B(n367), .ZN(n370) );
  XOR2_X1 U336 ( .A(n424), .B(n423), .Z(n573) );
  XOR2_X1 U337 ( .A(n457), .B(KEYINPUT28), .Z(n540) );
  XNOR2_X1 U338 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U339 ( .A(n459), .B(G127GAT), .ZN(n460) );
  XNOR2_X1 U340 ( .A(n471), .B(n470), .ZN(G1349GAT) );
  XOR2_X1 U341 ( .A(G120GAT), .B(G71GAT), .Z(n365) );
  XOR2_X1 U342 ( .A(G15GAT), .B(G127GAT), .Z(n378) );
  XNOR2_X1 U343 ( .A(n365), .B(n378), .ZN(n296) );
  XOR2_X1 U344 ( .A(KEYINPUT84), .B(KEYINPUT0), .Z(n295) );
  XNOR2_X1 U345 ( .A(G113GAT), .B(G134GAT), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n420) );
  XNOR2_X1 U347 ( .A(n296), .B(n420), .ZN(n302) );
  XOR2_X1 U348 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n298) );
  XNOR2_X1 U349 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n426) );
  XOR2_X1 U351 ( .A(G176GAT), .B(n426), .Z(n300) );
  NAND2_X1 U352 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U354 ( .A(n302), .B(n301), .Z(n310) );
  XOR2_X1 U355 ( .A(KEYINPUT20), .B(G190GAT), .Z(n304) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(G99GAT), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U358 ( .A(G183GAT), .B(KEYINPUT65), .Z(n306) );
  XNOR2_X1 U359 ( .A(KEYINPUT86), .B(KEYINPUT85), .ZN(n305) );
  XNOR2_X1 U360 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U362 ( .A(n310), .B(n309), .Z(n537) );
  INV_X1 U363 ( .A(n537), .ZN(n479) );
  XOR2_X1 U364 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n312) );
  XNOR2_X1 U365 ( .A(G43GAT), .B(G29GAT), .ZN(n311) );
  XNOR2_X1 U366 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U367 ( .A(KEYINPUT69), .B(n313), .Z(n343) );
  XOR2_X1 U368 ( .A(G92GAT), .B(n434), .Z(n315) );
  XNOR2_X1 U369 ( .A(G99GAT), .B(G85GAT), .ZN(n369) );
  XOR2_X1 U370 ( .A(G218GAT), .B(n369), .Z(n314) );
  XNOR2_X1 U371 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U372 ( .A(n343), .B(n316), .Z(n318) );
  NAND2_X1 U373 ( .A1(G232GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U375 ( .A(n319), .B(KEYINPUT9), .Z(n330) );
  XOR2_X1 U376 ( .A(KEYINPUT11), .B(KEYINPUT66), .Z(n321) );
  XNOR2_X1 U377 ( .A(G106GAT), .B(KEYINPUT77), .ZN(n320) );
  XNOR2_X1 U378 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U379 ( .A(KEYINPUT78), .B(KEYINPUT76), .Z(n323) );
  XNOR2_X1 U380 ( .A(KEYINPUT10), .B(KEYINPUT79), .ZN(n322) );
  XNOR2_X1 U381 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U382 ( .A(n325), .B(n324), .Z(n328) );
  XNOR2_X1 U383 ( .A(G50GAT), .B(KEYINPUT75), .ZN(n326) );
  XNOR2_X1 U384 ( .A(n326), .B(G162GAT), .ZN(n446) );
  XNOR2_X1 U385 ( .A(G134GAT), .B(n446), .ZN(n327) );
  XOR2_X1 U386 ( .A(KEYINPUT70), .B(G1GAT), .Z(n386) );
  XOR2_X1 U387 ( .A(G15GAT), .B(G50GAT), .Z(n332) );
  XNOR2_X1 U388 ( .A(G169GAT), .B(G36GAT), .ZN(n331) );
  XNOR2_X1 U389 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U390 ( .A(n386), .B(n333), .Z(n335) );
  NAND2_X1 U391 ( .A1(G229GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U393 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n337) );
  XNOR2_X1 U394 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U396 ( .A(n339), .B(n338), .Z(n345) );
  XOR2_X1 U397 ( .A(G22GAT), .B(G197GAT), .Z(n341) );
  XNOR2_X1 U398 ( .A(G113GAT), .B(G141GAT), .ZN(n340) );
  XNOR2_X1 U399 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U401 ( .A(n345), .B(n344), .Z(n519) );
  INV_X1 U402 ( .A(n519), .ZN(n577) );
  INV_X1 U403 ( .A(G148GAT), .ZN(n346) );
  NAND2_X1 U404 ( .A1(n346), .A2(G78GAT), .ZN(n349) );
  INV_X1 U405 ( .A(G78GAT), .ZN(n347) );
  NAND2_X1 U406 ( .A1(n347), .A2(G148GAT), .ZN(n348) );
  NAND2_X1 U407 ( .A1(n349), .A2(n348), .ZN(n351) );
  XNOR2_X1 U408 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n351), .B(n350), .ZN(n353) );
  INV_X1 U410 ( .A(n353), .ZN(n449) );
  INV_X1 U411 ( .A(KEYINPUT33), .ZN(n352) );
  NAND2_X1 U412 ( .A1(n449), .A2(n352), .ZN(n355) );
  NAND2_X1 U413 ( .A1(n353), .A2(KEYINPUT33), .ZN(n354) );
  NAND2_X1 U414 ( .A1(n355), .A2(n354), .ZN(n357) );
  AND2_X1 U415 ( .A1(G230GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U416 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U417 ( .A(KEYINPUT73), .B(KEYINPUT32), .Z(n359) );
  XNOR2_X1 U418 ( .A(KEYINPUT31), .B(KEYINPUT74), .ZN(n358) );
  XOR2_X1 U419 ( .A(n359), .B(n358), .Z(n360) );
  XNOR2_X1 U420 ( .A(n361), .B(n360), .ZN(n368) );
  XNOR2_X1 U421 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n362), .B(KEYINPUT13), .ZN(n377) );
  XOR2_X1 U423 ( .A(G64GAT), .B(G92GAT), .Z(n364) );
  XNOR2_X1 U424 ( .A(G176GAT), .B(G204GAT), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n425) );
  XNOR2_X1 U426 ( .A(n377), .B(n425), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n370), .B(n369), .ZN(n582) );
  NAND2_X1 U428 ( .A1(n577), .A2(n558), .ZN(n372) );
  INV_X1 U429 ( .A(KEYINPUT46), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n391) );
  XOR2_X1 U431 ( .A(KEYINPUT80), .B(KEYINPUT12), .Z(n374) );
  XNOR2_X1 U432 ( .A(G78GAT), .B(KEYINPUT14), .ZN(n373) );
  XNOR2_X1 U433 ( .A(n374), .B(n373), .ZN(n390) );
  XOR2_X1 U434 ( .A(G8GAT), .B(G183GAT), .Z(n430) );
  XOR2_X1 U435 ( .A(G22GAT), .B(G155GAT), .Z(n443) );
  XOR2_X1 U436 ( .A(n430), .B(n443), .Z(n376) );
  XNOR2_X1 U437 ( .A(G71GAT), .B(G211GAT), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n376), .B(n375), .ZN(n382) );
  XOR2_X1 U439 ( .A(n378), .B(n377), .Z(n380) );
  NAND2_X1 U440 ( .A1(G231GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U441 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U442 ( .A(n382), .B(n381), .Z(n388) );
  XOR2_X1 U443 ( .A(G64GAT), .B(KEYINPUT82), .Z(n384) );
  XNOR2_X1 U444 ( .A(KEYINPUT15), .B(KEYINPUT81), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U446 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U447 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n585) );
  NOR2_X1 U449 ( .A1(n391), .A2(n585), .ZN(n392) );
  XOR2_X1 U450 ( .A(n392), .B(KEYINPUT112), .Z(n393) );
  NOR2_X1 U451 ( .A1(n396), .A2(n393), .ZN(n394) );
  XNOR2_X1 U452 ( .A(KEYINPUT113), .B(n394), .ZN(n395) );
  XNOR2_X1 U453 ( .A(KEYINPUT47), .B(n395), .ZN(n402) );
  INV_X1 U454 ( .A(n585), .ZN(n503) );
  XOR2_X1 U455 ( .A(n396), .B(KEYINPUT36), .Z(n590) );
  NOR2_X1 U456 ( .A1(n503), .A2(n590), .ZN(n397) );
  XOR2_X1 U457 ( .A(n397), .B(KEYINPUT45), .Z(n398) );
  XOR2_X1 U458 ( .A(KEYINPUT114), .B(n399), .Z(n400) );
  NOR2_X1 U459 ( .A1(n577), .A2(n400), .ZN(n401) );
  NOR2_X1 U460 ( .A1(n402), .A2(n401), .ZN(n404) );
  XNOR2_X1 U461 ( .A(n404), .B(n403), .ZN(n463) );
  XOR2_X1 U462 ( .A(KEYINPUT4), .B(KEYINPUT92), .Z(n406) );
  XNOR2_X1 U463 ( .A(KEYINPUT91), .B(KEYINPUT1), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n424) );
  XOR2_X1 U465 ( .A(G155GAT), .B(G162GAT), .Z(n408) );
  XNOR2_X1 U466 ( .A(G120GAT), .B(G127GAT), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U468 ( .A(KEYINPUT93), .B(G57GAT), .Z(n410) );
  XNOR2_X1 U469 ( .A(G1GAT), .B(G148GAT), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U471 ( .A(n412), .B(n411), .Z(n418) );
  XNOR2_X1 U472 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n413) );
  XNOR2_X1 U473 ( .A(n413), .B(KEYINPUT2), .ZN(n451) );
  XOR2_X1 U474 ( .A(G85GAT), .B(n451), .Z(n415) );
  NAND2_X1 U475 ( .A1(G225GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U477 ( .A(G29GAT), .B(n416), .ZN(n417) );
  XNOR2_X1 U478 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U479 ( .A(n419), .B(KEYINPUT6), .Z(n422) );
  XNOR2_X1 U480 ( .A(n420), .B(KEYINPUT5), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n426), .B(n425), .ZN(n438) );
  XOR2_X1 U483 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n432) );
  XOR2_X1 U484 ( .A(KEYINPUT88), .B(G218GAT), .Z(n428) );
  XNOR2_X1 U485 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U487 ( .A(G197GAT), .B(n429), .Z(n452) );
  XNOR2_X1 U488 ( .A(n452), .B(n430), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U490 ( .A(n434), .B(n433), .Z(n436) );
  NAND2_X1 U491 ( .A1(G226GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U493 ( .A(n438), .B(n437), .Z(n534) );
  XNOR2_X1 U494 ( .A(n534), .B(KEYINPUT27), .ZN(n483) );
  NAND2_X1 U495 ( .A1(n573), .A2(n483), .ZN(n474) );
  NOR2_X1 U496 ( .A1(n463), .A2(n474), .ZN(n439) );
  XNOR2_X1 U497 ( .A(KEYINPUT115), .B(n439), .ZN(n555) );
  XOR2_X1 U498 ( .A(KEYINPUT23), .B(KEYINPUT87), .Z(n441) );
  XNOR2_X1 U499 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n440) );
  XNOR2_X1 U500 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U501 ( .A(n442), .B(KEYINPUT90), .Z(n445) );
  XNOR2_X1 U502 ( .A(n443), .B(KEYINPUT89), .ZN(n444) );
  XNOR2_X1 U503 ( .A(n445), .B(n444), .ZN(n456) );
  XOR2_X1 U504 ( .A(n446), .B(G204GAT), .Z(n448) );
  NAND2_X1 U505 ( .A1(G228GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n448), .B(n447), .ZN(n450) );
  XOR2_X1 U507 ( .A(n450), .B(n353), .Z(n454) );
  XNOR2_X1 U508 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U509 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U510 ( .A(n456), .B(n455), .Z(n480) );
  XNOR2_X1 U511 ( .A(n480), .B(KEYINPUT67), .ZN(n457) );
  OR2_X1 U512 ( .A1(n555), .A2(n540), .ZN(n458) );
  NAND2_X1 U513 ( .A1(n549), .A2(n585), .ZN(n461) );
  XOR2_X1 U514 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n459) );
  XNOR2_X1 U515 ( .A(n461), .B(n460), .ZN(G1342GAT) );
  XNOR2_X1 U516 ( .A(KEYINPUT106), .B(n558), .ZN(n546) );
  XOR2_X1 U517 ( .A(n534), .B(KEYINPUT124), .Z(n462) );
  NOR2_X1 U518 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U519 ( .A(n464), .B(KEYINPUT54), .ZN(n576) );
  NOR2_X1 U520 ( .A1(n573), .A2(n480), .ZN(n465) );
  AND2_X1 U521 ( .A1(n576), .A2(n465), .ZN(n466) );
  XNOR2_X1 U522 ( .A(n466), .B(KEYINPUT55), .ZN(n467) );
  NAND2_X1 U523 ( .A1(n546), .A2(n570), .ZN(n471) );
  XOR2_X1 U524 ( .A(G176GAT), .B(KEYINPUT57), .Z(n469) );
  XOR2_X1 U525 ( .A(KEYINPUT56), .B(KEYINPUT125), .Z(n468) );
  XOR2_X1 U526 ( .A(KEYINPUT34), .B(KEYINPUT99), .Z(n493) );
  OR2_X1 U527 ( .A1(n503), .A2(n396), .ZN(n472) );
  XNOR2_X1 U528 ( .A(n472), .B(KEYINPUT16), .ZN(n473) );
  XNOR2_X1 U529 ( .A(n473), .B(KEYINPUT83), .ZN(n490) );
  NOR2_X1 U530 ( .A1(n474), .A2(n540), .ZN(n475) );
  XNOR2_X1 U531 ( .A(KEYINPUT96), .B(n475), .ZN(n476) );
  NAND2_X1 U532 ( .A1(n479), .A2(n476), .ZN(n489) );
  AND2_X1 U533 ( .A1(n537), .A2(n534), .ZN(n477) );
  NOR2_X1 U534 ( .A1(n480), .A2(n477), .ZN(n478) );
  XNOR2_X1 U535 ( .A(n478), .B(KEYINPUT25), .ZN(n485) );
  XOR2_X1 U536 ( .A(KEYINPUT26), .B(KEYINPUT97), .Z(n482) );
  NAND2_X1 U537 ( .A1(n480), .A2(n479), .ZN(n481) );
  XOR2_X1 U538 ( .A(n482), .B(n481), .Z(n554) );
  NAND2_X1 U539 ( .A1(n483), .A2(n554), .ZN(n484) );
  NAND2_X1 U540 ( .A1(n485), .A2(n484), .ZN(n487) );
  INV_X1 U541 ( .A(n573), .ZN(n486) );
  NAND2_X1 U542 ( .A1(n487), .A2(n486), .ZN(n488) );
  NAND2_X1 U543 ( .A1(n489), .A2(n488), .ZN(n502) );
  NAND2_X1 U544 ( .A1(n490), .A2(n502), .ZN(n520) );
  OR2_X1 U545 ( .A1(n519), .A2(n582), .ZN(n507) );
  NOR2_X1 U546 ( .A1(n520), .A2(n507), .ZN(n491) );
  XNOR2_X1 U547 ( .A(n491), .B(KEYINPUT98), .ZN(n499) );
  NAND2_X1 U548 ( .A1(n573), .A2(n499), .ZN(n492) );
  XNOR2_X1 U549 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U550 ( .A(G1GAT), .B(n494), .ZN(G1324GAT) );
  NAND2_X1 U551 ( .A1(n499), .A2(n534), .ZN(n495) );
  XNOR2_X1 U552 ( .A(n495), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n497) );
  NAND2_X1 U554 ( .A1(n499), .A2(n537), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U556 ( .A(G15GAT), .B(n498), .ZN(G1326GAT) );
  XOR2_X1 U557 ( .A(G22GAT), .B(KEYINPUT101), .Z(n501) );
  NAND2_X1 U558 ( .A1(n499), .A2(n540), .ZN(n500) );
  XNOR2_X1 U559 ( .A(n501), .B(n500), .ZN(G1327GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n511) );
  NAND2_X1 U561 ( .A1(n503), .A2(n502), .ZN(n504) );
  NOR2_X1 U562 ( .A1(n590), .A2(n504), .ZN(n506) );
  XOR2_X1 U563 ( .A(KEYINPUT103), .B(KEYINPUT37), .Z(n505) );
  XNOR2_X1 U564 ( .A(n506), .B(n505), .ZN(n529) );
  NOR2_X1 U565 ( .A1(n529), .A2(n507), .ZN(n509) );
  XNOR2_X1 U566 ( .A(KEYINPUT104), .B(KEYINPUT38), .ZN(n508) );
  XNOR2_X1 U567 ( .A(n509), .B(n508), .ZN(n517) );
  NAND2_X1 U568 ( .A1(n517), .A2(n573), .ZN(n510) );
  XNOR2_X1 U569 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U570 ( .A(G29GAT), .B(n512), .ZN(G1328GAT) );
  NAND2_X1 U571 ( .A1(n534), .A2(n517), .ZN(n513) );
  XNOR2_X1 U572 ( .A(n513), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n515) );
  NAND2_X1 U574 ( .A1(n517), .A2(n537), .ZN(n514) );
  XNOR2_X1 U575 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U576 ( .A(G43GAT), .B(n516), .ZN(G1330GAT) );
  NAND2_X1 U577 ( .A1(n540), .A2(n517), .ZN(n518) );
  XNOR2_X1 U578 ( .A(n518), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n522) );
  NAND2_X1 U580 ( .A1(n546), .A2(n519), .ZN(n530) );
  NOR2_X1 U581 ( .A1(n530), .A2(n520), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n526), .A2(n573), .ZN(n521) );
  XNOR2_X1 U583 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U584 ( .A(G57GAT), .B(n523), .ZN(G1332GAT) );
  NAND2_X1 U585 ( .A1(n534), .A2(n526), .ZN(n524) );
  XNOR2_X1 U586 ( .A(n524), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U587 ( .A1(n537), .A2(n526), .ZN(n525) );
  XNOR2_X1 U588 ( .A(n525), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U589 ( .A(G78GAT), .B(KEYINPUT43), .Z(n528) );
  NAND2_X1 U590 ( .A1(n526), .A2(n540), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n528), .B(n527), .ZN(G1335GAT) );
  XOR2_X1 U592 ( .A(G85GAT), .B(KEYINPUT109), .Z(n533) );
  NOR2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U594 ( .A(n531), .B(KEYINPUT108), .ZN(n541) );
  NAND2_X1 U595 ( .A1(n573), .A2(n541), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(G1336GAT) );
  NAND2_X1 U597 ( .A1(n541), .A2(n534), .ZN(n535) );
  XNOR2_X1 U598 ( .A(n535), .B(KEYINPUT110), .ZN(n536) );
  XNOR2_X1 U599 ( .A(G92GAT), .B(n536), .ZN(G1337GAT) );
  XOR2_X1 U600 ( .A(G99GAT), .B(KEYINPUT111), .Z(n539) );
  NAND2_X1 U601 ( .A1(n541), .A2(n537), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n539), .B(n538), .ZN(G1338GAT) );
  NAND2_X1 U603 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U604 ( .A(n542), .B(KEYINPUT44), .ZN(n543) );
  XNOR2_X1 U605 ( .A(G106GAT), .B(n543), .ZN(G1339GAT) );
  NAND2_X1 U606 ( .A1(n549), .A2(n577), .ZN(n544) );
  XNOR2_X1 U607 ( .A(n544), .B(KEYINPUT116), .ZN(n545) );
  XNOR2_X1 U608 ( .A(G113GAT), .B(n545), .ZN(G1340GAT) );
  XOR2_X1 U609 ( .A(G120GAT), .B(KEYINPUT49), .Z(n548) );
  NAND2_X1 U610 ( .A1(n549), .A2(n546), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n548), .B(n547), .ZN(G1341GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U613 ( .A1(n549), .A2(n396), .ZN(n550) );
  XNOR2_X1 U614 ( .A(n551), .B(n550), .ZN(n553) );
  XOR2_X1 U615 ( .A(G134GAT), .B(KEYINPUT119), .Z(n552) );
  XNOR2_X1 U616 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  INV_X1 U617 ( .A(n554), .ZN(n574) );
  NOR2_X1 U618 ( .A1(n574), .A2(n555), .ZN(n564) );
  NAND2_X1 U619 ( .A1(n577), .A2(n564), .ZN(n556) );
  XNOR2_X1 U620 ( .A(KEYINPUT120), .B(n556), .ZN(n557) );
  XNOR2_X1 U621 ( .A(G141GAT), .B(n557), .ZN(G1344GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n560) );
  NAND2_X1 U623 ( .A1(n564), .A2(n558), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(n561), .ZN(G1345GAT) );
  XOR2_X1 U626 ( .A(G155GAT), .B(KEYINPUT121), .Z(n563) );
  NAND2_X1 U627 ( .A1(n564), .A2(n585), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(G1346GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n566) );
  NAND2_X1 U630 ( .A1(n564), .A2(n396), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(G162GAT), .B(n567), .ZN(G1347GAT) );
  NAND2_X1 U633 ( .A1(n570), .A2(n577), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U635 ( .A1(n585), .A2(n570), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U637 ( .A1(n570), .A2(n396), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(KEYINPUT58), .ZN(n572) );
  XNOR2_X1 U639 ( .A(G190GAT), .B(n572), .ZN(G1351GAT) );
  XNOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT126), .ZN(n581) );
  XOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT59), .Z(n579) );
  NOR2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n575) );
  AND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n588) );
  NAND2_X1 U644 ( .A1(n588), .A2(n577), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  NAND2_X1 U648 ( .A1(n588), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  XOR2_X1 U650 ( .A(G211GAT), .B(KEYINPUT127), .Z(n587) );
  NAND2_X1 U651 ( .A1(n588), .A2(n585), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1354GAT) );
  INV_X1 U653 ( .A(n588), .ZN(n589) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n592) );
  INV_X1 U655 ( .A(KEYINPUT62), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U657 ( .A(n593), .B(G218GAT), .ZN(G1355GAT) );
endmodule

