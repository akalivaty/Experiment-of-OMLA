//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1203;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  AND3_X1   g040(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT65), .ZN(new_n466));
  AOI21_X1  g041(.A(KEYINPUT65), .B1(new_n463), .B2(new_n465), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n461), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n462), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n473), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n464), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n474), .A2(new_n475), .A3(new_n461), .A4(new_n463), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n470), .A2(new_n478), .ZN(G160));
  NAND4_X1  g054(.A1(new_n474), .A2(new_n475), .A3(G2105), .A4(new_n463), .ZN(new_n480));
  INV_X1    g055(.A(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n461), .A2(G112), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  OAI22_X1  g058(.A1(new_n480), .A2(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n476), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(G136), .B2(new_n485), .ZN(G162));
  INV_X1    g061(.A(KEYINPUT65), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n464), .A2(G2104), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT65), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n493), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n493), .A2(G2105), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n474), .A2(new_n475), .A3(new_n495), .A4(new_n463), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n492), .A2(new_n494), .B1(KEYINPUT4), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n461), .A2(G114), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  OAI22_X1  g076(.A1(new_n480), .A2(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR3_X1   g077(.A1(new_n497), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n494), .B1(new_n466), .B2(new_n467), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n500), .A2(new_n501), .ZN(new_n507));
  INV_X1    g082(.A(new_n480), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(G126), .ZN(new_n509));
  AOI21_X1  g084(.A(KEYINPUT67), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n503), .A2(new_n510), .ZN(G164));
  XNOR2_X1  g086(.A(KEYINPUT68), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT6), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(G651), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n517), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G88), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(new_n512), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n513), .A2(G543), .A3(new_n516), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G50), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n526), .A2(new_n528), .A3(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n513), .A2(new_n516), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n536), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n535), .B1(new_n537), .B2(new_n524), .ZN(new_n538));
  INV_X1    g113(.A(G51), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT71), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n536), .A2(new_n540), .A3(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n529), .A2(KEYINPUT71), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n538), .A2(new_n543), .ZN(G168));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G64), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n524), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n512), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n525), .A2(G90), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G52), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n551), .B1(new_n541), .B2(new_n542), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n550), .A2(new_n552), .ZN(G171));
  NAND2_X1  g128(.A1(new_n541), .A2(new_n542), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G43), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT72), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n525), .A2(G81), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(G43), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(new_n541), .B2(new_n542), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT72), .B1(new_n561), .B2(new_n557), .ZN(new_n562));
  NAND2_X1  g137(.A1(G68), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G56), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n524), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n559), .A2(new_n562), .B1(new_n548), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n530), .A2(new_n572), .A3(G53), .ZN(new_n573));
  INV_X1    g148(.A(G53), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT9), .B1(new_n529), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n536), .A2(new_n523), .ZN(new_n577));
  INV_X1    g152(.A(G91), .ZN(new_n578));
  INV_X1    g153(.A(G651), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n523), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n577), .A2(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G299));
  INV_X1    g158(.A(G171), .ZN(G301));
  INV_X1    g159(.A(G168), .ZN(G286));
  NAND2_X1  g160(.A1(new_n525), .A2(G87), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n530), .A2(G49), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(new_n525), .A2(G86), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n523), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n591), .A2(new_n512), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n530), .A2(G48), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n590), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT73), .Z(G305));
  INV_X1    g170(.A(G85), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n577), .A2(new_n596), .B1(new_n512), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(G47), .B2(new_n554), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n554), .A2(G54), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT74), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(G66), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(G66), .ZN(new_n605));
  AND3_X1   g180(.A1(new_n523), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AND2_X1   g181(.A1(G79), .A2(G543), .ZN(new_n607));
  OAI21_X1  g182(.A(G651), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n513), .A2(new_n523), .A3(new_n516), .A4(G92), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n602), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n601), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n601), .B1(new_n613), .B2(G868), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n582), .ZN(G297));
  OAI21_X1  g192(.A(new_n616), .B1(G868), .B2(new_n582), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n613), .B1(new_n619), .B2(G860), .ZN(G148));
  INV_X1    g195(.A(new_n566), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n612), .A2(G559), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT75), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n622), .B1(new_n624), .B2(G868), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n492), .A2(new_n471), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT76), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT77), .B(KEYINPUT13), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT78), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n485), .A2(G135), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n508), .A2(G123), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n461), .A2(G111), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2096), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n640), .B1(new_n631), .B2(new_n632), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n634), .A2(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(KEYINPUT14), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n648), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2443), .B(G2446), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT79), .Z(new_n657));
  INV_X1    g232(.A(G14), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n654), .B2(new_n655), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT17), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n665), .B2(new_n662), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n666), .B1(KEYINPUT80), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(KEYINPUT80), .B2(new_n668), .ZN(new_n670));
  INV_X1    g245(.A(new_n662), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n671), .A2(new_n667), .A3(new_n664), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT18), .Z(new_n673));
  NAND3_X1  g248(.A1(new_n663), .A2(new_n667), .A3(new_n665), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2096), .B(G2100), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1971), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n678), .B(new_n679), .Z(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT20), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n681), .A2(KEYINPUT82), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n682), .A2(new_n683), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(new_n680), .B2(new_n684), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n687), .B(new_n689), .Z(new_n690));
  NAND2_X1  g265(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1981), .B(G1986), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT83), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n693), .B(new_n697), .ZN(G229));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G32), .ZN(new_n700));
  NAND3_X1  g275(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT95), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT26), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n485), .A2(G141), .B1(G105), .B2(new_n471), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n508), .A2(G129), .ZN(new_n705));
  AND3_X1   g280(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n700), .B1(new_n706), .B2(new_n699), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT96), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT27), .B(G1996), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT97), .Z(new_n711));
  NAND2_X1  g286(.A1(G164), .A2(G29), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G27), .B2(G29), .ZN(new_n713));
  INV_X1    g288(.A(G2078), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n699), .A2(G33), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT93), .B(KEYINPUT25), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n492), .A2(G127), .ZN(new_n720));
  NAND2_X1  g295(.A1(G115), .A2(G2104), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n461), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AOI211_X1 g297(.A(new_n719), .B(new_n722), .C1(G139), .C2(new_n485), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n716), .B1(new_n723), .B2(new_n699), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n724), .A2(G2072), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT94), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n713), .A2(new_n714), .ZN(new_n727));
  NOR4_X1   g302(.A1(new_n711), .A2(new_n715), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G16), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G20), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT23), .Z(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G299), .B2(G16), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G1956), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n699), .A2(G35), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G162), .B2(new_n699), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT29), .Z(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(G2090), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n699), .A2(G26), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT28), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n508), .A2(G128), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT92), .ZN(new_n742));
  OAI21_X1  g317(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n743));
  INV_X1    g318(.A(G116), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(G2105), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n485), .B2(G140), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n740), .B1(new_n747), .B2(new_n699), .ZN(new_n748));
  INV_X1    g323(.A(G2067), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n737), .A2(G2090), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n733), .A2(new_n738), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G171), .A2(new_n729), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G5), .B2(new_n729), .ZN(new_n754));
  INV_X1    g329(.A(G1961), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(G168), .A2(new_n729), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n729), .B2(G21), .ZN(new_n758));
  INV_X1    g333(.A(G1966), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n754), .A2(new_n755), .ZN(new_n761));
  INV_X1    g336(.A(G34), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n762), .A2(KEYINPUT24), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(KEYINPUT24), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n699), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G160), .B2(new_n699), .ZN(new_n766));
  INV_X1    g341(.A(G2084), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n756), .A2(new_n760), .A3(new_n761), .A4(new_n768), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT31), .B(G11), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT98), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT30), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n772), .A2(G28), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n699), .B1(new_n772), .B2(G28), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n771), .B1(new_n773), .B2(new_n774), .C1(new_n639), .C2(new_n699), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n724), .B2(G2072), .ZN(new_n776));
  OAI221_X1 g351(.A(new_n776), .B1(new_n708), .B2(new_n709), .C1(new_n759), .C2(new_n758), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n752), .A2(new_n769), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n729), .A2(G19), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n566), .B2(new_n729), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(G1341), .Z(new_n781));
  NOR2_X1   g356(.A1(G4), .A2(G16), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n613), .B2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT91), .ZN(new_n784));
  INV_X1    g359(.A(G1348), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n728), .A2(new_n778), .A3(new_n781), .A4(new_n786), .ZN(new_n787));
  MUX2_X1   g362(.A(G6), .B(G305), .S(G16), .Z(new_n788));
  XOR2_X1   g363(.A(KEYINPUT32), .B(G1981), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT87), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n788), .B(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(KEYINPUT88), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(KEYINPUT88), .ZN(new_n793));
  NOR2_X1   g368(.A1(G16), .A2(G22), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G166), .B2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT90), .B(G1971), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n729), .A2(G23), .ZN(new_n798));
  INV_X1    g373(.A(G288), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n729), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT33), .B(G1976), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT89), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n800), .B(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n792), .A2(new_n793), .A3(new_n797), .A4(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT86), .B(KEYINPUT34), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n729), .A2(G24), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n599), .B2(new_n729), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1986), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n699), .A2(G25), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(KEYINPUT84), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n811), .A2(KEYINPUT84), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n485), .A2(G131), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n508), .A2(G119), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n461), .A2(G107), .ZN(new_n816));
  OAI21_X1  g391(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n814), .B(new_n815), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT85), .ZN(new_n819));
  AOI211_X1 g394(.A(new_n812), .B(new_n813), .C1(new_n819), .C2(G29), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT35), .B(G1991), .Z(new_n821));
  AND2_X1   g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n810), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n806), .A2(new_n807), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(KEYINPUT36), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT36), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n806), .A2(new_n827), .A3(new_n807), .A4(new_n824), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n787), .B1(new_n826), .B2(new_n828), .ZN(G311));
  NAND2_X1  g404(.A1(new_n826), .A2(new_n828), .ZN(new_n830));
  INV_X1    g405(.A(new_n787), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(G150));
  NAND2_X1  g407(.A1(G80), .A2(G543), .ZN(new_n833));
  INV_X1    g408(.A(G67), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n524), .B2(new_n834), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n525), .A2(G93), .B1(new_n835), .B2(new_n548), .ZN(new_n836));
  INV_X1    g411(.A(new_n554), .ZN(new_n837));
  INV_X1    g412(.A(G55), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G860), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT101), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT100), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n843), .B(new_n836), .C1(new_n837), .C2(new_n838), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n565), .A2(new_n548), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n556), .B1(new_n555), .B2(new_n558), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n561), .A2(KEYINPUT72), .A3(new_n557), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n844), .B(new_n845), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n839), .A2(KEYINPUT100), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n849), .B1(new_n566), .B2(new_n844), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n613), .A2(G559), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n858), .A2(KEYINPUT39), .ZN(new_n859));
  INV_X1    g434(.A(G860), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n858), .B2(KEYINPUT39), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n842), .B1(new_n859), .B2(new_n861), .ZN(G145));
  INV_X1    g437(.A(G37), .ZN(new_n863));
  XNOR2_X1  g438(.A(G160), .B(new_n639), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(G162), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n485), .A2(G142), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT102), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n508), .A2(G130), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n461), .A2(G118), .ZN(new_n869));
  OAI21_X1  g444(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n867), .B(new_n868), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n818), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n723), .B(new_n706), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n506), .A2(new_n509), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n747), .B(new_n875), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(new_n629), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n874), .B(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(new_n865), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n879), .A2(KEYINPUT103), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(KEYINPUT103), .ZN(new_n881));
  OAI221_X1 g456(.A(new_n863), .B1(new_n865), .B2(new_n878), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g458(.A(new_n853), .B(new_n624), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n612), .A2(new_n582), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n612), .A2(new_n582), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(KEYINPUT104), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n612), .A2(new_n582), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n886), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n885), .A2(new_n895), .ZN(new_n897));
  AOI22_X1  g472(.A1(new_n896), .A2(KEYINPUT105), .B1(new_n887), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n899), .A3(new_n895), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n890), .B1(new_n884), .B2(new_n901), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n902), .A2(KEYINPUT42), .ZN(new_n903));
  XNOR2_X1  g478(.A(G305), .B(G303), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n599), .B(new_n799), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n904), .B1(KEYINPUT106), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(KEYINPUT106), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n906), .B(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n902), .A2(KEYINPUT42), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n903), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n909), .B1(new_n903), .B2(new_n910), .ZN(new_n912));
  OAI21_X1  g487(.A(G868), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n839), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n913), .B1(G868), .B2(new_n914), .ZN(G295));
  OAI21_X1  g490(.A(new_n913), .B1(G868), .B2(new_n914), .ZN(G331));
  INV_X1    g491(.A(KEYINPUT110), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n909), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(G171), .A2(KEYINPUT107), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(new_n550), .B2(new_n552), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(G168), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(G301), .A2(G286), .A3(new_n920), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n851), .B2(new_n852), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n848), .A2(new_n850), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n566), .A2(new_n849), .A3(new_n844), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n926), .A2(new_n927), .A3(new_n923), .A4(new_n922), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(KEYINPUT108), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n930), .B(new_n924), .C1(new_n851), .C2(new_n852), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(KEYINPUT109), .A3(new_n888), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n925), .A2(new_n928), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n901), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n889), .B1(new_n929), .B2(new_n931), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n937), .A2(KEYINPUT109), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n918), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n940));
  AOI22_X1  g515(.A1(new_n937), .A2(KEYINPUT109), .B1(new_n901), .B2(new_n934), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n932), .A2(new_n888), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n909), .A2(new_n917), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n941), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n939), .A2(new_n940), .A3(new_n946), .A4(new_n863), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT111), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n891), .A2(new_n893), .ZN(new_n951));
  AOI22_X1  g526(.A1(new_n951), .A2(new_n897), .B1(new_n888), .B2(new_n895), .ZN(new_n952));
  OAI22_X1  g527(.A1(new_n932), .A2(new_n952), .B1(new_n889), .B2(new_n934), .ZN(new_n953));
  AOI21_X1  g528(.A(G37), .B1(new_n953), .B2(new_n909), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n941), .A2(new_n944), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n954), .B1(new_n955), .B2(new_n909), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n950), .B1(new_n956), .B2(KEYINPUT43), .ZN(new_n957));
  AOI21_X1  g532(.A(G37), .B1(new_n955), .B2(new_n918), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n958), .A2(KEYINPUT111), .A3(new_n940), .A4(new_n946), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n949), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n940), .B1(new_n958), .B2(new_n946), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n950), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n960), .A2(new_n963), .ZN(G397));
  INV_X1    g539(.A(KEYINPUT127), .ZN(new_n965));
  INV_X1    g540(.A(new_n478), .ZN(new_n966));
  INV_X1    g541(.A(new_n469), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(new_n492), .B2(G125), .ZN(new_n968));
  OAI211_X1 g543(.A(G40), .B(new_n966), .C1(new_n968), .C2(new_n461), .ZN(new_n969));
  AOI21_X1  g544(.A(G1384), .B1(new_n506), .B2(new_n509), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n969), .A2(new_n970), .A3(KEYINPUT45), .ZN(new_n971));
  OR2_X1    g546(.A1(new_n971), .A2(KEYINPUT112), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(KEYINPUT112), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n747), .B(G2067), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n706), .B(G1996), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n818), .B(new_n821), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n599), .B(G1986), .Z(new_n979));
  OAI21_X1  g554(.A(new_n974), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G8), .ZN(new_n982));
  INV_X1    g557(.A(G40), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n470), .A2(new_n983), .A3(new_n478), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n982), .B1(new_n984), .B2(new_n970), .ZN(new_n985));
  INV_X1    g560(.A(G1976), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n985), .B1(new_n986), .B2(G288), .ZN(new_n987));
  NAND2_X1  g562(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OR3_X1    g564(.A1(new_n799), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n987), .A2(new_n988), .ZN(new_n992));
  INV_X1    g567(.A(G1981), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n993), .B1(new_n592), .B2(new_n994), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n995), .A2(new_n594), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n594), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(KEYINPUT49), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT49), .B1(new_n996), .B2(new_n997), .ZN(new_n999));
  INV_X1    g574(.A(new_n985), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n991), .A2(new_n992), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(G303), .A2(G8), .ZN(new_n1003));
  XOR2_X1   g578(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1005), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n969), .B1(new_n1008), .B2(new_n970), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n498), .B1(new_n497), .B2(new_n502), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n506), .A2(new_n509), .A3(KEYINPUT67), .ZN(new_n1011));
  AOI21_X1  g586(.A(G1384), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1009), .B1(new_n1012), .B2(new_n1008), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1013), .A2(G2090), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n970), .A2(KEYINPUT45), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT113), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n1012), .B2(KEYINPUT45), .ZN(new_n1017));
  INV_X1    g592(.A(G1384), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(new_n503), .B2(new_n510), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(KEYINPUT113), .A3(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1017), .A2(new_n1021), .A3(new_n984), .ZN(new_n1022));
  INV_X1    g597(.A(G1971), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1014), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1022), .A2(KEYINPUT114), .A3(new_n1023), .ZN(new_n1027));
  AOI211_X1 g602(.A(new_n982), .B(new_n1007), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(KEYINPUT45), .B(new_n1018), .C1(new_n503), .C2(new_n510), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1018), .B1(new_n497), .B2(new_n502), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n969), .B1(new_n1020), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n759), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1009), .B(new_n767), .C1(new_n1008), .C2(new_n1012), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n982), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT63), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1036), .A3(G168), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1024), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1030), .A2(KEYINPUT50), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1039), .A2(KEYINPUT118), .A3(new_n984), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1008), .B(new_n1018), .C1(new_n503), .C2(new_n510), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT118), .B1(new_n1039), .B2(new_n984), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1042), .A2(G2090), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(G8), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1037), .B1(new_n1045), .B2(new_n1007), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1002), .B1(new_n1028), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1007), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1014), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(new_n1027), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1048), .B1(new_n1051), .B2(G8), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1002), .A2(G168), .A3(new_n1035), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT63), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI211_X1 g629(.A(G1976), .B(G288), .C1(new_n1001), .C2(new_n998), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n594), .A2(G1981), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n985), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1047), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n582), .B(KEYINPUT57), .ZN(new_n1059));
  INV_X1    g634(.A(G1956), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT56), .B(G2072), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1017), .A2(new_n1021), .A3(new_n984), .A4(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1059), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1061), .A2(new_n1063), .A3(new_n1059), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n984), .A2(new_n1066), .A3(new_n970), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT119), .B1(new_n969), .B2(new_n1030), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1013), .A2(new_n785), .B1(new_n1069), .B2(new_n749), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(new_n612), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1064), .B1(new_n1065), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1061), .A2(new_n1063), .A3(new_n1059), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1074), .A2(new_n1064), .ZN(new_n1075));
  INV_X1    g650(.A(G1996), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1017), .A2(new_n1021), .A3(new_n1076), .A4(new_n984), .ZN(new_n1077));
  XOR2_X1   g652(.A(KEYINPUT58), .B(G1341), .Z(new_n1078));
  NAND3_X1  g653(.A1(new_n1067), .A2(new_n1068), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n566), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT59), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(new_n1083), .A3(new_n566), .ZN(new_n1084));
  AOI22_X1  g659(.A1(KEYINPUT61), .A2(new_n1075), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1059), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n1065), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT61), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1013), .A2(new_n785), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1069), .A2(new_n749), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(KEYINPUT60), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n613), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1070), .A2(KEYINPUT60), .A3(new_n612), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1070), .A2(KEYINPUT60), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1089), .A2(new_n1090), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1073), .B1(new_n1085), .B2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(G171), .B(KEYINPUT54), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1008), .B(new_n1018), .C1(new_n497), .C2(new_n502), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n984), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n1019), .B2(KEYINPUT50), .ZN(new_n1103));
  OR3_X1    g678(.A1(new_n1103), .A2(KEYINPUT122), .A3(G1961), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT122), .B1(new_n1103), .B2(G1961), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1031), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n970), .A2(KEYINPUT45), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT123), .B1(new_n1108), .B2(new_n969), .ZN(new_n1109));
  OR2_X1    g684(.A1(KEYINPUT124), .A2(G2078), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(KEYINPUT124), .B2(G2078), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1015), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1107), .A2(new_n1109), .A3(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1104), .A2(new_n1105), .A3(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1111), .B1(new_n1022), .B2(G2078), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1100), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1032), .A2(new_n1111), .A3(G2078), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n755), .B2(new_n1013), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1100), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(new_n1116), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1103), .A2(new_n767), .B1(new_n1032), .B2(new_n759), .ZN(new_n1124));
  NOR2_X1   g699(.A1(G168), .A2(new_n982), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1125), .B1(KEYINPUT120), .B2(KEYINPUT51), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1124), .B2(new_n982), .ZN(new_n1129));
  NOR2_X1   g704(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1127), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1130), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1128), .B(new_n1132), .C1(new_n1124), .C2(new_n982), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT121), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1126), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1130), .B1(new_n1035), .B2(new_n1136), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1138));
  AND4_X1   g713(.A1(KEYINPUT121), .A2(new_n1137), .A3(new_n1133), .A4(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1123), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1099), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n992), .A2(new_n990), .A3(new_n989), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1001), .A2(new_n998), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1144), .B1(new_n1045), .B2(new_n1007), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1051), .A2(G8), .A3(new_n1048), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT125), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1145), .A2(new_n1146), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1058), .B1(new_n1141), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1131), .A2(KEYINPUT121), .A3(new_n1133), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1137), .A2(new_n1133), .A3(new_n1138), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1153), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(KEYINPUT62), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1159));
  AOI21_X1  g734(.A(G301), .B1(new_n1120), .B2(new_n1116), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1151), .A2(new_n1158), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n981), .B1(new_n1152), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n974), .A2(new_n1076), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT46), .ZN(new_n1164));
  INV_X1    g739(.A(new_n974), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n975), .A2(new_n706), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT47), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1167), .B(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(new_n819), .ZN(new_n1170));
  AND4_X1   g745(.A1(new_n821), .A2(new_n975), .A3(new_n1170), .A4(new_n976), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n747), .A2(new_n749), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n974), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT126), .ZN(new_n1174));
  NOR2_X1   g749(.A1(G290), .A2(G1986), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n974), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1177), .A2(KEYINPUT48), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n1177), .A2(KEYINPUT48), .ZN(new_n1179));
  AOI211_X1 g754(.A(new_n1178), .B(new_n1179), .C1(new_n974), .C2(new_n978), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1169), .A2(new_n1174), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n965), .B1(new_n1162), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1088), .A2(KEYINPUT61), .A3(new_n1065), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1090), .B1(new_n1074), .B2(new_n1064), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1072), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1190));
  AOI22_X1  g765(.A1(new_n1153), .A2(new_n1156), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1191));
  AND3_X1   g766(.A1(new_n1145), .A2(new_n1146), .A3(new_n1149), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1149), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1190), .B(new_n1191), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1194));
  AND3_X1   g769(.A1(new_n1047), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1159), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1197));
  OAI211_X1 g772(.A(new_n1194), .B(new_n1195), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1198), .A2(new_n980), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1199), .A2(KEYINPUT127), .A3(new_n1181), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1183), .A2(new_n1200), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g776(.A1(G401), .A2(new_n459), .A3(G227), .A4(G229), .ZN(new_n1203));
  OAI211_X1 g777(.A(new_n882), .B(new_n1203), .C1(new_n961), .C2(new_n962), .ZN(G225));
  INV_X1    g778(.A(G225), .ZN(G308));
endmodule


