//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT15), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(KEYINPUT87), .A3(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G36gat), .ZN(new_n206));
  AND2_X1   g005(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G29gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n210), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT87), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT15), .B1(new_n202), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n205), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(KEYINPUT88), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n209), .A2(KEYINPUT15), .A3(new_n202), .A4(new_n211), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G15gat), .B(G22gat), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n219), .A2(G1gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT89), .ZN(new_n221));
  AOI21_X1  g020(.A(G8gat), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT16), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n219), .B1(new_n223), .B2(G1gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(new_n222), .B(new_n225), .Z(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n218), .A2(new_n227), .ZN(new_n228));
  AND3_X1   g027(.A1(new_n216), .A2(KEYINPUT17), .A3(new_n217), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n229), .A2(KEYINPUT90), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n229), .A2(KEYINPUT90), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n218), .A2(KEYINPUT17), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(new_n226), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n228), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G229gat), .A2(G233gat), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT18), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n234), .B1(new_n230), .B2(new_n231), .ZN(new_n238));
  INV_X1    g037(.A(new_n228), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n238), .A2(KEYINPUT18), .A3(new_n239), .A4(new_n236), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n218), .A2(new_n227), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(new_n236), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n237), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT91), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n240), .A2(new_n248), .A3(new_n245), .ZN(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G141gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(G197gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT11), .B(G169gat), .ZN(new_n252));
  XOR2_X1   g051(.A(new_n251), .B(new_n252), .Z(new_n253));
  XOR2_X1   g052(.A(KEYINPUT86), .B(KEYINPUT12), .Z(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n249), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n247), .A2(new_n256), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n249), .B(new_n255), .C1(new_n237), .C2(new_n246), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G15gat), .B(G43gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(G71gat), .B(G99gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G227gat), .ZN(new_n264));
  INV_X1    g063(.A(G233gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G113gat), .B(G120gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n270));
  XNOR2_X1  g069(.A(G127gat), .B(G134gat), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n268), .B(new_n269), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(G127gat), .B(G134gat), .Z(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n269), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n273), .B(new_n274), .C1(new_n267), .C2(KEYINPUT1), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT23), .ZN(new_n277));
  NOR3_X1   g076(.A1(new_n277), .A2(G169gat), .A3(G176gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT66), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT66), .ZN(new_n282));
  INV_X1    g081(.A(G169gat), .ZN(new_n283));
  INV_X1    g082(.A(G176gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n282), .B(new_n279), .C1(new_n285), .C2(new_n277), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT25), .ZN(new_n288));
  NOR2_X1   g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT65), .B1(new_n289), .B2(KEYINPUT23), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT65), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n291), .B(new_n277), .C1(G169gat), .C2(G176gat), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n288), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n294));
  INV_X1    g093(.A(G183gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G190gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT69), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n296), .A2(new_n301), .A3(new_n297), .A4(new_n298), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT67), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n305), .A2(new_n306), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n304), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n287), .B(new_n293), .C1(new_n303), .C2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n297), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n297), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n304), .B(new_n311), .C1(new_n312), .C2(KEYINPUT24), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n290), .A2(new_n292), .ZN(new_n314));
  OR2_X1    g113(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n315), .A2(KEYINPUT23), .A3(new_n283), .A4(new_n316), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n313), .A2(new_n314), .A3(new_n279), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n288), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n310), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT70), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT70), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n310), .A2(new_n322), .A3(new_n319), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT27), .B(G183gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n297), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n312), .B1(new_n326), .B2(KEYINPUT28), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n296), .A2(KEYINPUT27), .A3(new_n298), .ZN(new_n328));
  OR3_X1    g127(.A1(new_n295), .A2(KEYINPUT71), .A3(KEYINPUT27), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT71), .B1(new_n295), .B2(KEYINPUT27), .ZN(new_n330));
  NOR2_X1   g129(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n328), .A2(new_n329), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n280), .B1(KEYINPUT26), .B2(new_n285), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n333), .B1(KEYINPUT26), .B2(new_n285), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n327), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n276), .B1(new_n324), .B2(new_n335), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n310), .A2(new_n322), .A3(new_n319), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n322), .B1(new_n310), .B2(new_n319), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n276), .B(new_n335), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n266), .B1(new_n336), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n263), .B1(new_n341), .B2(KEYINPUT32), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT73), .ZN(new_n343));
  INV_X1    g142(.A(new_n266), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n335), .B1(new_n337), .B2(new_n338), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n272), .A2(new_n275), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n344), .B1(new_n347), .B2(new_n339), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n343), .B1(new_n348), .B2(KEYINPUT33), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT33), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n341), .A2(KEYINPUT73), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n342), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n341), .B(KEYINPUT32), .C1(new_n350), .C2(new_n263), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n347), .A2(new_n344), .A3(new_n339), .ZN(new_n354));
  XNOR2_X1  g153(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n354), .B(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n352), .A2(new_n353), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT75), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n352), .A2(new_n360), .A3(new_n353), .A4(new_n357), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT36), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n364));
  INV_X1    g163(.A(new_n353), .ZN(new_n365));
  NOR3_X1   g164(.A1(new_n348), .A2(new_n343), .A3(KEYINPUT33), .ZN(new_n366));
  INV_X1    g165(.A(new_n263), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT32), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n367), .B1(new_n348), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n365), .B1(new_n370), .B2(new_n349), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n364), .B1(new_n371), .B2(new_n357), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n352), .A2(new_n353), .ZN(new_n373));
  INV_X1    g172(.A(new_n357), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(KEYINPUT76), .A3(new_n374), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n362), .A2(new_n363), .A3(new_n372), .A4(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n374), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n358), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT36), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G228gat), .A2(G233gat), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n383));
  XOR2_X1   g182(.A(G211gat), .B(G218gat), .Z(new_n384));
  XOR2_X1   g183(.A(G197gat), .B(G204gat), .Z(new_n385));
  AOI21_X1  g184(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G211gat), .B(G218gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(G197gat), .B(G204gat), .ZN(new_n389));
  INV_X1    g188(.A(G211gat), .ZN(new_n390));
  INV_X1    g189(.A(G218gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n388), .B(new_n389), .C1(KEYINPUT22), .C2(new_n392), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n387), .A2(KEYINPUT80), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT29), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n395), .B1(new_n393), .B2(KEYINPUT80), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n383), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(G141gat), .A2(G148gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G155gat), .A2(G162gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT2), .ZN(new_n401));
  NAND2_X1  g200(.A1(G141gat), .A2(G148gat), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n400), .ZN(new_n404));
  NOR2_X1   g203(.A1(G155gat), .A2(G162gat), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT78), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(G155gat), .ZN(new_n407));
  INV_X1    g206(.A(G162gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT78), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(new_n400), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n403), .A2(new_n406), .A3(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n404), .A2(new_n405), .ZN(new_n413));
  AND2_X1   g212(.A1(G141gat), .A2(G148gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(new_n398), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n413), .A2(new_n415), .A3(new_n410), .A4(new_n401), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n387), .A2(new_n393), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT3), .B1(new_n412), .B2(new_n416), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n419), .B1(new_n420), .B2(KEYINPUT29), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT81), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n397), .A2(new_n417), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n419), .B(KEYINPUT81), .C1(new_n420), .C2(KEYINPUT29), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n382), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT29), .B1(new_n387), .B2(new_n393), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n417), .B1(new_n426), .B2(KEYINPUT3), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n421), .A2(new_n427), .A3(new_n382), .ZN(new_n428));
  OAI21_X1  g227(.A(G22gat), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n397), .A2(new_n417), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n421), .A2(new_n422), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n424), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n428), .B1(new_n432), .B2(new_n381), .ZN(new_n433));
  INV_X1    g232(.A(G22gat), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT82), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n434), .ZN(new_n436));
  XOR2_X1   g235(.A(G78gat), .B(G106gat), .Z(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT31), .B(G50gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  AND4_X1   g238(.A1(new_n429), .A2(new_n435), .A3(new_n436), .A4(new_n439), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n435), .A2(new_n439), .B1(new_n429), .B2(new_n436), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G1gat), .B(G29gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(KEYINPUT0), .ZN(new_n444));
  XNOR2_X1  g243(.A(G57gat), .B(G85gat), .ZN(new_n445));
  XOR2_X1   g244(.A(new_n444), .B(new_n445), .Z(new_n446));
  NAND2_X1  g245(.A1(new_n412), .A2(new_n416), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n346), .B(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(G225gat), .A2(G233gat), .ZN(new_n449));
  OR2_X1    g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n276), .A2(KEYINPUT4), .A3(new_n447), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT4), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n452), .B1(new_n417), .B2(new_n346), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n447), .A2(new_n383), .B1(new_n272), .B2(new_n275), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n417), .A2(KEYINPUT3), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT79), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT79), .B1(new_n455), .B2(new_n456), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n454), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n449), .ZN(new_n460));
  OAI211_X1 g259(.A(KEYINPUT5), .B(new_n450), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n451), .A2(new_n453), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n455), .A2(new_n456), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT79), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT79), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT5), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n468), .A3(new_n449), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n446), .B1(new_n461), .B2(new_n469), .ZN(new_n470));
  XOR2_X1   g269(.A(KEYINPUT84), .B(KEYINPUT39), .Z(new_n471));
  NOR3_X1   g270(.A1(new_n467), .A2(KEYINPUT83), .A3(new_n449), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT83), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n473), .B1(new_n459), .B2(new_n460), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n471), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT83), .B1(new_n467), .B2(new_n449), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n459), .A2(new_n473), .A3(new_n460), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n448), .A2(new_n449), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT39), .A4(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n475), .A2(new_n446), .A3(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(KEYINPUT85), .B(KEYINPUT40), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n470), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT77), .ZN(new_n483));
  NAND2_X1  g282(.A1(G226gat), .A2(G233gat), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n345), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n484), .B1(new_n324), .B2(new_n335), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT29), .B1(new_n320), .B2(new_n335), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT77), .B1(new_n488), .B2(new_n485), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n486), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n418), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n320), .A2(new_n335), .A3(new_n485), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n485), .A2(KEYINPUT29), .ZN(new_n493));
  AOI211_X1 g292(.A(new_n418), .B(new_n492), .C1(new_n345), .C2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G8gat), .B(G36gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(G64gat), .B(G92gat), .ZN(new_n497));
  XOR2_X1   g296(.A(new_n496), .B(new_n497), .Z(new_n498));
  NAND3_X1  g297(.A1(new_n491), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n498), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n327), .A2(new_n332), .A3(new_n334), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n501), .B1(new_n319), .B2(new_n310), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n484), .B1(new_n502), .B2(KEYINPUT29), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n501), .B1(new_n321), .B2(new_n323), .ZN(new_n504));
  OAI211_X1 g303(.A(KEYINPUT77), .B(new_n503), .C1(new_n504), .C2(new_n484), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n419), .B1(new_n505), .B2(new_n486), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n500), .B1(new_n506), .B2(new_n494), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n499), .A2(new_n507), .A3(KEYINPUT30), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n494), .B1(new_n490), .B2(new_n418), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT30), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n510), .A3(new_n498), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n475), .A2(new_n479), .A3(KEYINPUT40), .A4(new_n446), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n482), .A2(new_n508), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT37), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n498), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n490), .A2(new_n419), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n492), .B1(new_n345), .B2(new_n493), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n514), .B1(new_n517), .B2(new_n418), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT38), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n461), .A2(new_n469), .A3(new_n446), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT6), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n470), .ZN(new_n524));
  INV_X1    g323(.A(new_n470), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(new_n522), .A3(new_n521), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n520), .A2(new_n524), .A3(new_n526), .A4(new_n499), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT38), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT37), .B1(new_n506), .B2(new_n494), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n528), .B1(new_n515), .B2(new_n529), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n442), .B(new_n513), .C1(new_n527), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n508), .A2(new_n511), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n526), .A2(new_n524), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n442), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n376), .A2(new_n380), .A3(new_n531), .A4(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT76), .B1(new_n373), .B2(new_n374), .ZN(new_n538));
  AOI211_X1 g337(.A(new_n364), .B(new_n357), .C1(new_n352), .C2(new_n353), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT35), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n532), .A2(new_n533), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n540), .A2(new_n542), .A3(new_n362), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n377), .A2(new_n358), .A3(new_n442), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT35), .B1(new_n544), .B2(new_n534), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n260), .B1(new_n537), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(G57gat), .B(G64gat), .ZN(new_n549));
  XOR2_X1   g348(.A(G71gat), .B(G78gat), .Z(new_n550));
  INV_X1    g349(.A(KEYINPUT93), .ZN(new_n551));
  AOI211_X1 g350(.A(new_n548), .B(new_n549), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n550), .A2(new_n551), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT94), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT21), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G127gat), .B(G155gat), .Z(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n227), .B1(new_n556), .B2(new_n557), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n561), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G231gat), .A2(G233gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT95), .ZN(new_n566));
  XOR2_X1   g365(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G183gat), .B(G211gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n564), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n562), .A2(new_n563), .A3(new_n570), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n218), .ZN(new_n576));
  NOR2_X1   g375(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n577));
  INV_X1    g376(.A(G85gat), .ZN(new_n578));
  INV_X1    g377(.A(G92gat), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(G99gat), .ZN(new_n581));
  INV_X1    g380(.A(G106gat), .ZN(new_n582));
  OAI21_X1  g381(.A(KEYINPUT8), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n580), .B(new_n583), .C1(G85gat), .C2(G92gat), .ZN(new_n584));
  AND2_X1   g383(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n585));
  NOR4_X1   g384(.A1(new_n585), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT97), .ZN(new_n588));
  XOR2_X1   g387(.A(G99gat), .B(G106gat), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n587), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(KEYINPUT97), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594));
  AOI22_X1  g393(.A1(new_n576), .A2(new_n593), .B1(KEYINPUT41), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n233), .A2(new_n593), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n596), .B1(new_n232), .B2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(G190gat), .B(G218gat), .Z(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n597), .B1(new_n230), .B2(new_n231), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n601), .A2(new_n599), .A3(new_n595), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT98), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n601), .A2(KEYINPUT98), .A3(new_n599), .A4(new_n595), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n600), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT99), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n607), .B1(new_n604), .B2(new_n605), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n594), .A2(KEYINPUT41), .ZN(new_n609));
  XNOR2_X1  g408(.A(G134gat), .B(G162gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NOR3_X1   g411(.A1(new_n606), .A2(new_n608), .A3(new_n612), .ZN(new_n613));
  AOI221_X4 g412(.A(new_n600), .B1(new_n607), .B2(new_n611), .C1(new_n604), .C2(new_n605), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n575), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT100), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT98), .B1(new_n598), .B2(new_n599), .ZN(new_n618));
  INV_X1    g417(.A(new_n605), .ZN(new_n619));
  OAI22_X1  g418(.A1(new_n618), .A2(new_n619), .B1(new_n599), .B2(new_n598), .ZN(new_n620));
  OAI21_X1  g419(.A(KEYINPUT99), .B1(new_n618), .B2(new_n619), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n620), .A2(new_n621), .A3(new_n611), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n606), .B1(new_n608), .B2(new_n612), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(KEYINPUT100), .A3(new_n575), .ZN(new_n625));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n587), .B1(KEYINPUT101), .B2(new_n590), .ZN(new_n628));
  OR3_X1    g427(.A1(new_n587), .A2(KEYINPUT101), .A3(new_n590), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n554), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(KEYINPUT102), .B(KEYINPUT10), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n554), .B(KEYINPUT94), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n630), .B(new_n631), .C1(new_n632), .C2(new_n593), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n632), .A2(KEYINPUT10), .A3(new_n593), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n627), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n630), .B1(new_n632), .B2(new_n593), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n635), .B1(new_n627), .B2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G120gat), .B(G148gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(G176gat), .B(G204gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n638), .B(new_n639), .Z(new_n640));
  OR2_X1    g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n635), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n636), .A2(new_n627), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(new_n643), .A3(new_n640), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  AND4_X1   g445(.A1(new_n547), .A2(new_n617), .A3(new_n625), .A4(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n533), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G1gat), .ZN(G1324gat));
  INV_X1    g449(.A(new_n532), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT16), .B(G8gat), .Z(new_n652));
  AND3_X1   g451(.A1(new_n647), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(G8gat), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n654), .B1(new_n647), .B2(new_n651), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT42), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(KEYINPUT42), .B2(new_n653), .ZN(G1325gat));
  INV_X1    g456(.A(G15gat), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n540), .A2(new_n362), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n647), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n376), .A2(new_n380), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n647), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n661), .B1(new_n663), .B2(new_n658), .ZN(G1326gat));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n535), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT43), .B(G22gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1327gat));
  NOR2_X1   g466(.A1(new_n613), .A2(new_n614), .ZN(new_n668));
  AND4_X1   g467(.A1(new_n547), .A2(new_n668), .A3(new_n574), .A4(new_n646), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n669), .A2(new_n210), .A3(new_n648), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT45), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n537), .A2(new_n546), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT104), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n537), .A2(new_n546), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n668), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n624), .B1(new_n537), .B2(new_n546), .ZN(new_n679));
  OAI22_X1  g478(.A1(new_n676), .A2(new_n678), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n645), .B(KEYINPUT103), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n681), .A2(new_n260), .A3(new_n575), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n533), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n671), .B1(new_n210), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT105), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n671), .B(new_n687), .C1(new_n210), .C2(new_n684), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(G1328gat));
  NAND3_X1  g488(.A1(new_n669), .A2(new_n206), .A3(new_n651), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT46), .Z(new_n691));
  OAI21_X1  g490(.A(G36gat), .B1(new_n683), .B2(new_n532), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(G1329gat));
  INV_X1    g492(.A(new_n662), .ZN(new_n694));
  OAI21_X1  g493(.A(G43gat), .B1(new_n683), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(G43gat), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n669), .A2(new_n696), .A3(new_n660), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1330gat));
  AND3_X1   g499(.A1(new_n537), .A2(new_n546), .A3(new_n674), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n674), .B1(new_n537), .B2(new_n546), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n701), .A2(new_n702), .A3(new_n678), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n679), .A2(new_n677), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n535), .B(new_n682), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT107), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n680), .A2(new_n707), .A3(new_n535), .A4(new_n682), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n706), .A2(new_n708), .A3(G50gat), .ZN(new_n709));
  INV_X1    g508(.A(G50gat), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n669), .A2(new_n710), .A3(new_n535), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT48), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n705), .A2(G50gat), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n711), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT48), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n714), .A2(KEYINPUT108), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n710), .B1(new_n705), .B2(KEYINPUT107), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n712), .B1(new_n721), .B2(new_n708), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT48), .B1(new_n715), .B2(new_n711), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n720), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n719), .A2(new_n724), .ZN(G1331gat));
  NOR2_X1   g524(.A1(new_n701), .A2(new_n702), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT100), .B1(new_n624), .B2(new_n575), .ZN(new_n727));
  AOI211_X1 g526(.A(new_n616), .B(new_n574), .C1(new_n622), .C2(new_n623), .ZN(new_n728));
  INV_X1    g527(.A(new_n681), .ZN(new_n729));
  NOR4_X1   g528(.A1(new_n727), .A2(new_n728), .A3(new_n729), .A4(new_n259), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n533), .B(KEYINPUT109), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g534(.A1(new_n731), .A2(new_n532), .ZN(new_n736));
  NOR2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  AND2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n736), .B2(new_n737), .ZN(G1333gat));
  OAI21_X1  g539(.A(G71gat), .B1(new_n731), .B2(new_n694), .ZN(new_n741));
  OR2_X1    g540(.A1(new_n659), .A2(G71gat), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n731), .B2(new_n742), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g543(.A1(new_n731), .A2(new_n442), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT110), .B(G78gat), .Z(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1335gat));
  NAND3_X1  g546(.A1(new_n679), .A2(new_n260), .A3(new_n574), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT51), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(new_n646), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n750), .A2(new_n578), .A3(new_n648), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n259), .A2(new_n575), .A3(new_n646), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n680), .A2(new_n752), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n753), .A2(new_n648), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n751), .B1(new_n754), .B2(new_n578), .ZN(G1336gat));
  AOI21_X1  g554(.A(new_n579), .B1(new_n753), .B2(new_n651), .ZN(new_n756));
  NOR2_X1   g555(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n748), .B(new_n757), .Z(new_n758));
  NAND3_X1  g557(.A1(new_n681), .A2(new_n579), .A3(new_n651), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT52), .B1(new_n756), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n749), .B2(new_n759), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n756), .B2(new_n763), .ZN(G1337gat));
  NAND3_X1  g563(.A1(new_n750), .A2(new_n581), .A3(new_n660), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n753), .A2(new_n662), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n765), .B1(new_n766), .B2(new_n581), .ZN(G1338gat));
  NAND3_X1  g566(.A1(new_n680), .A2(new_n535), .A3(new_n752), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n582), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n769), .B2(new_n768), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n729), .A2(G106gat), .A3(new_n442), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n749), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(KEYINPUT53), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n768), .A2(G106gat), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n758), .A2(new_n773), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT53), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n779), .ZN(G1339gat));
  INV_X1    g579(.A(new_n733), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n633), .A2(new_n627), .A3(new_n634), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n642), .A2(KEYINPUT54), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n640), .B1(new_n635), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n783), .A2(KEYINPUT55), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n644), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT55), .B1(new_n783), .B2(new_n785), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT113), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n783), .A2(new_n785), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n792), .A2(new_n793), .A3(new_n644), .A4(new_n786), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n259), .A2(new_n789), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n255), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n238), .A2(new_n239), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n797), .A2(G229gat), .A3(G233gat), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n242), .A2(new_n244), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI22_X1  g599(.A1(new_n247), .A2(new_n796), .B1(new_n253), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n645), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n668), .B1(new_n795), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n622), .A2(new_n801), .A3(new_n623), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n794), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n574), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n617), .A2(new_n260), .A3(new_n625), .A4(new_n646), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n781), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n544), .A2(new_n651), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(G113gat), .B1(new_n811), .B2(new_n259), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n535), .B1(new_n807), .B2(new_n808), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n651), .A2(new_n533), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(new_n660), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(G113gat), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n815), .A2(new_n816), .A3(new_n260), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n812), .A2(new_n817), .ZN(G1340gat));
  AOI21_X1  g617(.A(G120gat), .B1(new_n811), .B2(new_n645), .ZN(new_n819));
  INV_X1    g618(.A(G120gat), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n815), .A2(new_n820), .A3(new_n729), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n819), .A2(new_n821), .ZN(G1341gat));
  OAI21_X1  g621(.A(G127gat), .B1(new_n815), .B2(new_n574), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n809), .A2(new_n810), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n574), .A2(G127gat), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(G1342gat));
  INV_X1    g625(.A(KEYINPUT56), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n824), .A2(G134gat), .A3(new_n624), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n624), .A2(G134gat), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n811), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(KEYINPUT114), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n827), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(G134gat), .B1(new_n815), .B2(new_n624), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n828), .A2(new_n829), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n832), .A2(KEYINPUT114), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n836), .A2(new_n837), .A3(KEYINPUT56), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n834), .A2(new_n835), .A3(new_n838), .ZN(G1343gat));
  INV_X1    g638(.A(new_n814), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n662), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g640(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n842), .B1(new_n783), .B2(new_n785), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n787), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n259), .A2(new_n844), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n845), .A2(new_n802), .B1(new_n623), .B2(new_n622), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n574), .B1(new_n846), .B2(new_n806), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n442), .B1(new_n847), .B2(new_n808), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n841), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI211_X1 g649(.A(KEYINPUT57), .B(new_n442), .C1(new_n807), .C2(new_n808), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n850), .A2(new_n851), .A3(new_n260), .ZN(new_n852));
  INV_X1    g651(.A(G141gat), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT118), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT116), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n809), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n694), .A2(new_n535), .A3(new_n532), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n857), .B1(new_n809), .B2(new_n855), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n259), .A2(new_n853), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT117), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n856), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n861), .B1(new_n852), .B2(new_n853), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n854), .A2(new_n862), .A3(KEYINPUT58), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT58), .ZN(new_n864));
  OAI221_X1 g663(.A(new_n861), .B1(KEYINPUT118), .B2(new_n864), .C1(new_n852), .C2(new_n853), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(G1344gat));
  AND2_X1   g665(.A1(new_n856), .A2(new_n858), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n646), .A2(G148gat), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n867), .A2(KEYINPUT119), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT119), .B1(new_n867), .B2(new_n868), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(G148gat), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n850), .A2(new_n851), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(new_n645), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n442), .A2(KEYINPUT57), .ZN(new_n875));
  INV_X1    g674(.A(new_n808), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n845), .A2(new_n802), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n624), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n787), .A2(new_n788), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n668), .A2(new_n801), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n575), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n875), .B1(new_n876), .B2(new_n881), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n662), .A2(new_n646), .A3(new_n840), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n442), .B1(new_n807), .B2(new_n808), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n882), .B(new_n883), .C1(new_n884), .C2(new_n849), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n871), .B1(new_n885), .B2(G148gat), .ZN(new_n886));
  OAI22_X1  g685(.A1(new_n869), .A2(new_n870), .B1(new_n874), .B2(new_n886), .ZN(G1345gat));
  NAND3_X1  g686(.A1(new_n867), .A2(new_n407), .A3(new_n575), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n850), .A2(new_n851), .A3(new_n574), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(new_n407), .ZN(G1346gat));
  AOI21_X1  g689(.A(G162gat), .B1(new_n867), .B2(new_n668), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n624), .A2(new_n408), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n873), .B2(new_n892), .ZN(G1347gat));
  AOI21_X1  g692(.A(new_n648), .B1(new_n807), .B2(new_n808), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n544), .A2(new_n532), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(G169gat), .B1(new_n896), .B2(new_n259), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n733), .A2(new_n532), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n659), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n813), .A2(new_n900), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n901), .A2(new_n283), .A3(new_n260), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n897), .A2(new_n902), .ZN(G1348gat));
  AOI21_X1  g702(.A(G176gat), .B1(new_n896), .B2(new_n645), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n904), .A2(KEYINPUT120), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(KEYINPUT120), .ZN(new_n906));
  INV_X1    g705(.A(new_n901), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n729), .B1(new_n315), .B2(new_n316), .ZN(new_n908));
  AOI22_X1  g707(.A1(new_n905), .A2(new_n906), .B1(new_n907), .B2(new_n908), .ZN(G1349gat));
  NAND3_X1  g708(.A1(new_n896), .A2(new_n325), .A3(new_n575), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n296), .A2(new_n298), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n911), .B1(new_n901), .B2(new_n574), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g712(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n913), .B(new_n915), .ZN(G1350gat));
  NAND3_X1  g715(.A1(new_n896), .A2(new_n297), .A3(new_n668), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n813), .A2(new_n668), .A3(new_n900), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G190gat), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT122), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n918), .A2(new_n922), .A3(G190gat), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n921), .B1(new_n920), .B2(new_n923), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n917), .B1(new_n924), .B2(new_n925), .ZN(G1351gat));
  XNOR2_X1  g725(.A(KEYINPUT123), .B(G197gat), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n899), .A2(new_n662), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n882), .B(new_n928), .C1(new_n884), .C2(new_n849), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n927), .B1(new_n929), .B2(new_n260), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n662), .A2(new_n442), .A3(new_n532), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n894), .A2(new_n931), .ZN(new_n932));
  OR3_X1    g731(.A1(new_n932), .A2(new_n260), .A3(new_n927), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n930), .A2(new_n933), .A3(KEYINPUT124), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1352gat));
  INV_X1    g737(.A(new_n932), .ZN(new_n939));
  INV_X1    g738(.A(G204gat), .ZN(new_n940));
  NAND2_X1  g739(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n939), .A2(new_n940), .A3(new_n645), .A4(new_n941), .ZN(new_n942));
  XNOR2_X1  g741(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n645), .A2(new_n940), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n932), .B2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n946), .B1(new_n929), .B2(new_n729), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(G204gat), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n929), .A2(new_n946), .A3(new_n729), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n942), .B(new_n945), .C1(new_n948), .C2(new_n949), .ZN(G1353gat));
  NAND3_X1  g749(.A1(new_n939), .A2(new_n390), .A3(new_n575), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n929), .A2(new_n574), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT63), .B1(new_n952), .B2(G211gat), .ZN(new_n953));
  OAI211_X1 g752(.A(KEYINPUT63), .B(G211gat), .C1(new_n929), .C2(new_n574), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n951), .B1(new_n953), .B2(new_n955), .ZN(G1354gat));
  OAI21_X1  g755(.A(G218gat), .B1(new_n929), .B2(new_n624), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n939), .A2(new_n391), .A3(new_n668), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1355gat));
endmodule


