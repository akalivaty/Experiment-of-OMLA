

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593;

  NOR2_X2 U326 ( .A1(n412), .A2(n411), .ZN(n413) );
  XNOR2_X1 U327 ( .A(n495), .B(KEYINPUT37), .ZN(n496) );
  XNOR2_X1 U328 ( .A(n325), .B(n324), .ZN(n528) );
  XNOR2_X1 U329 ( .A(KEYINPUT47), .B(KEYINPUT114), .ZN(n405) );
  INV_X1 U330 ( .A(KEYINPUT80), .ZN(n315) );
  XNOR2_X1 U331 ( .A(n327), .B(KEYINPUT73), .ZN(n328) );
  XNOR2_X1 U332 ( .A(n406), .B(n405), .ZN(n412) );
  XNOR2_X1 U333 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U334 ( .A(n452), .B(n328), .ZN(n332) );
  NOR2_X1 U335 ( .A1(n551), .A2(n488), .ZN(n537) );
  XNOR2_X1 U336 ( .A(n318), .B(n317), .ZN(n320) );
  XNOR2_X1 U337 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U338 ( .A(n497), .B(n496), .ZN(n525) );
  XNOR2_X1 U339 ( .A(n339), .B(n338), .ZN(n582) );
  XNOR2_X1 U340 ( .A(n402), .B(n401), .ZN(n560) );
  XNOR2_X1 U341 ( .A(n501), .B(n500), .ZN(n509) );
  XNOR2_X1 U342 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U343 ( .A(n462), .B(n461), .ZN(G1351GAT) );
  XOR2_X1 U344 ( .A(G15GAT), .B(G127GAT), .Z(n365) );
  XOR2_X1 U345 ( .A(G134GAT), .B(G190GAT), .Z(n295) );
  XNOR2_X1 U346 ( .A(G43GAT), .B(G99GAT), .ZN(n294) );
  XNOR2_X1 U347 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U348 ( .A(n365), .B(n296), .Z(n298) );
  NAND2_X1 U349 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n312) );
  XOR2_X1 U351 ( .A(G71GAT), .B(KEYINPUT85), .Z(n300) );
  XNOR2_X1 U352 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U354 ( .A(G176GAT), .B(KEYINPUT20), .Z(n302) );
  XNOR2_X1 U355 ( .A(G169GAT), .B(KEYINPUT86), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U357 ( .A(n304), .B(n303), .Z(n310) );
  XOR2_X1 U358 ( .A(G120GAT), .B(KEYINPUT0), .Z(n306) );
  XNOR2_X1 U359 ( .A(G113GAT), .B(KEYINPUT82), .ZN(n305) );
  XNOR2_X1 U360 ( .A(n306), .B(n305), .ZN(n416) );
  XOR2_X1 U361 ( .A(G183GAT), .B(KEYINPUT19), .Z(n308) );
  XNOR2_X1 U362 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n307) );
  XNOR2_X1 U363 ( .A(n308), .B(n307), .ZN(n323) );
  XNOR2_X1 U364 ( .A(n416), .B(n323), .ZN(n309) );
  XNOR2_X1 U365 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U366 ( .A(n312), .B(n311), .ZN(n530) );
  XOR2_X1 U367 ( .A(G36GAT), .B(G190GAT), .Z(n392) );
  XOR2_X1 U368 ( .A(G64GAT), .B(G92GAT), .Z(n314) );
  XNOR2_X1 U369 ( .A(G176GAT), .B(G204GAT), .ZN(n313) );
  XNOR2_X1 U370 ( .A(n314), .B(n313), .ZN(n335) );
  XOR2_X1 U371 ( .A(n392), .B(n335), .Z(n318) );
  NAND2_X1 U372 ( .A1(G226GAT), .A2(G233GAT), .ZN(n316) );
  XOR2_X1 U373 ( .A(G169GAT), .B(G8GAT), .Z(n352) );
  XNOR2_X1 U374 ( .A(n352), .B(KEYINPUT93), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n325) );
  XOR2_X1 U376 ( .A(G211GAT), .B(KEYINPUT21), .Z(n322) );
  XNOR2_X1 U377 ( .A(G197GAT), .B(G218GAT), .ZN(n321) );
  XNOR2_X1 U378 ( .A(n322), .B(n321), .ZN(n453) );
  XOR2_X1 U379 ( .A(n323), .B(n453), .Z(n324) );
  XNOR2_X1 U380 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n340) );
  XNOR2_X1 U381 ( .A(G106GAT), .B(G78GAT), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n326), .B(G148GAT), .ZN(n452) );
  AND2_X1 U383 ( .A1(G230GAT), .A2(G233GAT), .ZN(n327) );
  XOR2_X1 U384 ( .A(KEYINPUT33), .B(KEYINPUT74), .Z(n330) );
  XNOR2_X1 U385 ( .A(KEYINPUT75), .B(KEYINPUT32), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U387 ( .A(n332), .B(n331), .Z(n339) );
  XOR2_X1 U388 ( .A(G99GAT), .B(G85GAT), .Z(n386) );
  XNOR2_X1 U389 ( .A(G120GAT), .B(n386), .ZN(n333) );
  XNOR2_X1 U390 ( .A(n333), .B(KEYINPUT31), .ZN(n337) );
  XNOR2_X1 U391 ( .A(G71GAT), .B(G57GAT), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n334), .B(KEYINPUT13), .ZN(n368) );
  XNOR2_X1 U393 ( .A(n335), .B(n368), .ZN(n336) );
  XNOR2_X1 U394 ( .A(n340), .B(n582), .ZN(n555) );
  XOR2_X1 U395 ( .A(KEYINPUT72), .B(KEYINPUT29), .Z(n342) );
  XNOR2_X1 U396 ( .A(KEYINPUT67), .B(KEYINPUT69), .ZN(n341) );
  XNOR2_X1 U397 ( .A(n342), .B(n341), .ZN(n356) );
  XOR2_X1 U398 ( .A(G15GAT), .B(G113GAT), .Z(n344) );
  XNOR2_X1 U399 ( .A(G36GAT), .B(G50GAT), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U401 ( .A(KEYINPUT68), .B(G22GAT), .Z(n346) );
  XNOR2_X1 U402 ( .A(G197GAT), .B(G141GAT), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U404 ( .A(n348), .B(n347), .Z(n354) );
  XOR2_X1 U405 ( .A(KEYINPUT71), .B(G1GAT), .Z(n375) );
  XOR2_X1 U406 ( .A(n375), .B(KEYINPUT30), .Z(n350) );
  NAND2_X1 U407 ( .A1(G229GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U410 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U412 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n358) );
  XNOR2_X1 U413 ( .A(G43GAT), .B(G29GAT), .ZN(n357) );
  XNOR2_X1 U414 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U415 ( .A(KEYINPUT7), .B(n359), .ZN(n399) );
  XOR2_X1 U416 ( .A(n360), .B(n399), .Z(n512) );
  INV_X1 U417 ( .A(n512), .ZN(n579) );
  NAND2_X1 U418 ( .A1(n555), .A2(n579), .ZN(n362) );
  XOR2_X1 U419 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n404) );
  XOR2_X1 U421 ( .A(KEYINPUT80), .B(G78GAT), .Z(n364) );
  XNOR2_X1 U422 ( .A(G183GAT), .B(G211GAT), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n364), .B(n363), .ZN(n379) );
  XOR2_X1 U424 ( .A(G22GAT), .B(G155GAT), .Z(n440) );
  XOR2_X1 U425 ( .A(n440), .B(n365), .Z(n367) );
  NAND2_X1 U426 ( .A1(G231GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n367), .B(n366), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n368), .B(KEYINPUT81), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n369), .B(KEYINPUT12), .ZN(n370) );
  XOR2_X1 U430 ( .A(n371), .B(n370), .Z(n377) );
  XOR2_X1 U431 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n373) );
  XNOR2_X1 U432 ( .A(G8GAT), .B(G64GAT), .ZN(n372) );
  XNOR2_X1 U433 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U435 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n585) );
  XNOR2_X1 U437 ( .A(G106GAT), .B(G92GAT), .ZN(n381) );
  INV_X1 U438 ( .A(KEYINPUT9), .ZN(n380) );
  XNOR2_X1 U439 ( .A(n381), .B(n380), .ZN(n383) );
  XOR2_X1 U440 ( .A(KEYINPUT79), .B(KEYINPUT66), .Z(n382) );
  XNOR2_X1 U441 ( .A(n383), .B(n382), .ZN(n385) );
  XOR2_X1 U442 ( .A(G134GAT), .B(KEYINPUT77), .Z(n428) );
  XNOR2_X1 U443 ( .A(G218GAT), .B(n428), .ZN(n384) );
  XNOR2_X1 U444 ( .A(n385), .B(n384), .ZN(n388) );
  NAND2_X1 U445 ( .A1(n388), .A2(n387), .ZN(n390) );
  INV_X1 U446 ( .A(n386), .ZN(n387) );
  OR2_X1 U447 ( .A1(n388), .A2(n387), .ZN(n389) );
  NAND2_X1 U448 ( .A1(n390), .A2(n389), .ZN(n394) );
  XNOR2_X1 U449 ( .A(G50GAT), .B(KEYINPUT76), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n391), .B(G162GAT), .ZN(n445) );
  XNOR2_X1 U451 ( .A(n445), .B(n392), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U453 ( .A(KEYINPUT10), .B(KEYINPUT78), .Z(n396) );
  NAND2_X1 U454 ( .A1(G232GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U455 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U456 ( .A(n398), .B(n397), .ZN(n402) );
  INV_X1 U457 ( .A(n399), .ZN(n400) );
  XOR2_X1 U458 ( .A(n400), .B(KEYINPUT11), .Z(n401) );
  NOR2_X1 U459 ( .A1(n585), .A2(n560), .ZN(n403) );
  NAND2_X1 U460 ( .A1(n404), .A2(n403), .ZN(n406) );
  XOR2_X1 U461 ( .A(KEYINPUT36), .B(n560), .Z(n590) );
  INV_X1 U462 ( .A(n585), .ZN(n493) );
  NOR2_X1 U463 ( .A1(n590), .A2(n493), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n407), .B(KEYINPUT45), .ZN(n410) );
  INV_X1 U465 ( .A(n582), .ZN(n408) );
  NOR2_X1 U466 ( .A1(n579), .A2(n408), .ZN(n409) );
  AND2_X1 U467 ( .A1(n410), .A2(n409), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n413), .B(KEYINPUT48), .ZN(n553) );
  NOR2_X1 U469 ( .A1(n528), .A2(n553), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n414), .B(KEYINPUT54), .ZN(n437) );
  XNOR2_X1 U471 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n415), .B(KEYINPUT2), .ZN(n439) );
  XNOR2_X1 U473 ( .A(n416), .B(n439), .ZN(n436) );
  XOR2_X1 U474 ( .A(G57GAT), .B(G155GAT), .Z(n418) );
  XNOR2_X1 U475 ( .A(G1GAT), .B(G148GAT), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U477 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n420) );
  XNOR2_X1 U478 ( .A(KEYINPUT4), .B(KEYINPUT90), .ZN(n419) );
  XNOR2_X1 U479 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U480 ( .A(n422), .B(n421), .Z(n434) );
  XOR2_X1 U481 ( .A(KEYINPUT5), .B(KEYINPUT89), .Z(n424) );
  XNOR2_X1 U482 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n423) );
  XNOR2_X1 U483 ( .A(n424), .B(n423), .ZN(n432) );
  XOR2_X1 U484 ( .A(G85GAT), .B(G162GAT), .Z(n426) );
  XNOR2_X1 U485 ( .A(G29GAT), .B(G127GAT), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U487 ( .A(n428), .B(n427), .Z(n430) );
  NAND2_X1 U488 ( .A1(G225GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U490 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n526) );
  NAND2_X1 U493 ( .A1(n437), .A2(n526), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n438), .B(KEYINPUT65), .ZN(n576) );
  XOR2_X1 U495 ( .A(n440), .B(n439), .Z(n442) );
  NAND2_X1 U496 ( .A1(G228GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n444) );
  INV_X1 U498 ( .A(KEYINPUT88), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n447) );
  XNOR2_X1 U500 ( .A(n445), .B(KEYINPUT87), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n447), .B(n446), .ZN(n451) );
  XOR2_X1 U502 ( .A(G204GAT), .B(KEYINPUT24), .Z(n449) );
  XNOR2_X1 U503 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n448) );
  XOR2_X1 U504 ( .A(n449), .B(n448), .Z(n450) );
  XNOR2_X1 U505 ( .A(n451), .B(n450), .ZN(n455) );
  XNOR2_X1 U506 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n455), .B(n454), .ZN(n474) );
  NAND2_X1 U508 ( .A1(n576), .A2(n474), .ZN(n456) );
  XOR2_X1 U509 ( .A(n456), .B(KEYINPUT55), .Z(n457) );
  NOR2_X1 U510 ( .A1(n530), .A2(n457), .ZN(n458) );
  XNOR2_X1 U511 ( .A(n458), .B(KEYINPUT118), .ZN(n567) );
  BUF_X1 U512 ( .A(n567), .Z(n572) );
  NAND2_X1 U513 ( .A1(n572), .A2(n560), .ZN(n462) );
  XOR2_X1 U514 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n460) );
  XNOR2_X1 U515 ( .A(G190GAT), .B(KEYINPUT122), .ZN(n459) );
  NAND2_X1 U516 ( .A1(n579), .A2(n582), .ZN(n498) );
  NOR2_X1 U517 ( .A1(n560), .A2(n493), .ZN(n463) );
  XNOR2_X1 U518 ( .A(KEYINPUT16), .B(n463), .ZN(n478) );
  OR2_X1 U519 ( .A1(n530), .A2(n528), .ZN(n464) );
  NAND2_X1 U520 ( .A1(n474), .A2(n464), .ZN(n465) );
  XNOR2_X1 U521 ( .A(n465), .B(KEYINPUT25), .ZN(n469) );
  XNOR2_X1 U522 ( .A(KEYINPUT26), .B(KEYINPUT95), .ZN(n467) );
  INV_X1 U523 ( .A(n530), .ZN(n538) );
  NOR2_X1 U524 ( .A1(n538), .A2(n474), .ZN(n466) );
  XNOR2_X1 U525 ( .A(n467), .B(n466), .ZN(n578) );
  XNOR2_X1 U526 ( .A(KEYINPUT27), .B(n528), .ZN(n472) );
  NOR2_X1 U527 ( .A1(n578), .A2(n472), .ZN(n468) );
  NOR2_X1 U528 ( .A1(n469), .A2(n468), .ZN(n470) );
  XOR2_X1 U529 ( .A(KEYINPUT96), .B(n470), .Z(n471) );
  NAND2_X1 U530 ( .A1(n471), .A2(n526), .ZN(n476) );
  NOR2_X1 U531 ( .A1(n526), .A2(n472), .ZN(n473) );
  XOR2_X1 U532 ( .A(KEYINPUT94), .B(n473), .Z(n551) );
  XOR2_X1 U533 ( .A(n474), .B(KEYINPUT28), .Z(n488) );
  NAND2_X1 U534 ( .A1(n537), .A2(n530), .ZN(n475) );
  NAND2_X1 U535 ( .A1(n476), .A2(n475), .ZN(n477) );
  XOR2_X1 U536 ( .A(KEYINPUT97), .B(n477), .Z(n492) );
  NAND2_X1 U537 ( .A1(n478), .A2(n492), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n479), .B(KEYINPUT98), .ZN(n513) );
  NOR2_X1 U539 ( .A1(n498), .A2(n513), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n480), .B(KEYINPUT99), .ZN(n489) );
  NOR2_X1 U541 ( .A1(n526), .A2(n489), .ZN(n482) );
  XNOR2_X1 U542 ( .A(KEYINPUT34), .B(KEYINPUT100), .ZN(n481) );
  XNOR2_X1 U543 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U544 ( .A(G1GAT), .B(n483), .Z(G1324GAT) );
  NOR2_X1 U545 ( .A1(n528), .A2(n489), .ZN(n484) );
  XOR2_X1 U546 ( .A(G8GAT), .B(n484), .Z(G1325GAT) );
  NOR2_X1 U547 ( .A1(n530), .A2(n489), .ZN(n486) );
  XNOR2_X1 U548 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n485) );
  XNOR2_X1 U549 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U550 ( .A(G15GAT), .B(n487), .Z(G1326GAT) );
  INV_X1 U551 ( .A(n488), .ZN(n533) );
  NOR2_X1 U552 ( .A1(n533), .A2(n489), .ZN(n490) );
  XOR2_X1 U553 ( .A(KEYINPUT102), .B(n490), .Z(n491) );
  XNOR2_X1 U554 ( .A(G22GAT), .B(n491), .ZN(G1327GAT) );
  INV_X1 U555 ( .A(KEYINPUT38), .ZN(n501) );
  NAND2_X1 U556 ( .A1(n493), .A2(n492), .ZN(n494) );
  NOR2_X1 U557 ( .A1(n590), .A2(n494), .ZN(n497) );
  INV_X1 U558 ( .A(KEYINPUT103), .ZN(n495) );
  NOR2_X1 U559 ( .A1(n498), .A2(n525), .ZN(n499) );
  XNOR2_X1 U560 ( .A(KEYINPUT104), .B(n499), .ZN(n500) );
  NOR2_X1 U561 ( .A1(n526), .A2(n509), .ZN(n503) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  NOR2_X1 U564 ( .A1(n528), .A2(n509), .ZN(n504) );
  XOR2_X1 U565 ( .A(G36GAT), .B(n504), .Z(G1329GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n506) );
  XNOR2_X1 U567 ( .A(G43GAT), .B(KEYINPUT105), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n506), .B(n505), .ZN(n508) );
  NOR2_X1 U569 ( .A1(n530), .A2(n509), .ZN(n507) );
  XOR2_X1 U570 ( .A(n508), .B(n507), .Z(G1330GAT) );
  NOR2_X1 U571 ( .A1(n533), .A2(n509), .ZN(n511) );
  XNOR2_X1 U572 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n511), .B(n510), .ZN(G1331GAT) );
  XNOR2_X1 U574 ( .A(KEYINPUT108), .B(n555), .ZN(n566) );
  NAND2_X1 U575 ( .A1(n512), .A2(n566), .ZN(n524) );
  OR2_X1 U576 ( .A1(n513), .A2(n524), .ZN(n521) );
  NOR2_X1 U577 ( .A1(n526), .A2(n521), .ZN(n515) );
  XNOR2_X1 U578 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U580 ( .A(G57GAT), .B(n516), .ZN(G1332GAT) );
  NOR2_X1 U581 ( .A1(n528), .A2(n521), .ZN(n517) );
  XOR2_X1 U582 ( .A(KEYINPUT110), .B(n517), .Z(n518) );
  XNOR2_X1 U583 ( .A(G64GAT), .B(n518), .ZN(G1333GAT) );
  NOR2_X1 U584 ( .A1(n530), .A2(n521), .ZN(n520) );
  XNOR2_X1 U585 ( .A(G71GAT), .B(KEYINPUT111), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(G1334GAT) );
  NOR2_X1 U587 ( .A1(n533), .A2(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(G1335GAT) );
  OR2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n532) );
  NOR2_X1 U591 ( .A1(n526), .A2(n532), .ZN(n527) );
  XOR2_X1 U592 ( .A(G85GAT), .B(n527), .Z(G1336GAT) );
  NOR2_X1 U593 ( .A1(n528), .A2(n532), .ZN(n529) );
  XOR2_X1 U594 ( .A(G92GAT), .B(n529), .Z(G1337GAT) );
  NOR2_X1 U595 ( .A1(n530), .A2(n532), .ZN(n531) );
  XOR2_X1 U596 ( .A(G99GAT), .B(n531), .Z(G1338GAT) );
  NOR2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n535) );
  XNOR2_X1 U598 ( .A(KEYINPUT112), .B(KEYINPUT44), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U600 ( .A(G106GAT), .B(n536), .Z(G1339GAT) );
  NAND2_X1 U601 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U602 ( .A1(n553), .A2(n539), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n579), .A2(n547), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n540), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U606 ( .A1(n547), .A2(n566), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U608 ( .A(G120GAT), .B(n543), .Z(G1341GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n545) );
  NAND2_X1 U610 ( .A1(n547), .A2(n585), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U612 ( .A(G127GAT), .B(n546), .Z(G1342GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n549) );
  NAND2_X1 U614 ( .A1(n547), .A2(n560), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U616 ( .A(G134GAT), .B(n550), .Z(G1343GAT) );
  OR2_X1 U617 ( .A1(n578), .A2(n551), .ZN(n552) );
  NOR2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n561) );
  AND2_X1 U619 ( .A1(n579), .A2(n561), .ZN(n554) );
  XOR2_X1 U620 ( .A(G141GAT), .B(n554), .Z(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n557) );
  NAND2_X1 U622 ( .A1(n561), .A2(n555), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n585), .A2(n561), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n567), .A2(n579), .ZN(n564) );
  XOR2_X1 U630 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n569) );
  XOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT57), .Z(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n571) );
  XOR2_X1 U636 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  NAND2_X1 U638 ( .A1(n572), .A2(n585), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n574), .B(KEYINPUT124), .ZN(n575) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(n575), .Z(n581) );
  INV_X1 U643 ( .A(n576), .ZN(n577) );
  NOR2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n586) );
  NAND2_X1 U645 ( .A1(n586), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  INV_X1 U648 ( .A(n586), .ZN(n589) );
  OR2_X1 U649 ( .A1(n589), .A2(n582), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  XOR2_X1 U651 ( .A(G211GAT), .B(KEYINPUT125), .Z(n588) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n592) );
  XNOR2_X1 U655 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n592), .B(n591), .ZN(n593) );
  XOR2_X1 U657 ( .A(G218GAT), .B(n593), .Z(G1355GAT) );
endmodule

