//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT76), .ZN(new_n189));
  OR2_X1    g003(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G104), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n190), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G101), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n191), .A2(G104), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G104), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G107), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n194), .A2(new_n195), .A3(new_n197), .A4(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(G101), .B1(new_n199), .B2(new_n196), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT1), .B1(new_n207), .B2(G146), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(G128), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G128), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n206), .B(new_n208), .C1(KEYINPUT1), .C2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n189), .B1(new_n204), .B2(new_n214), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n211), .A2(new_n213), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n216), .A2(KEYINPUT76), .A3(new_n202), .A4(new_n203), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n204), .A2(new_n214), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n215), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G137), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(KEYINPUT11), .A3(G134), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT11), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G137), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT65), .A2(G131), .ZN(new_n225));
  OR2_X1    g039(.A1(KEYINPUT64), .A2(G134), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n220), .A2(KEYINPUT11), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT64), .A2(G134), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n224), .A2(new_n225), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n225), .B1(new_n224), .B2(new_n229), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n219), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT12), .ZN(new_n235));
  XOR2_X1   g049(.A(KEYINPUT77), .B(KEYINPUT10), .Z(new_n236));
  NAND3_X1  g050(.A1(new_n215), .A2(new_n217), .A3(new_n236), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n216), .A2(KEYINPUT10), .A3(new_n202), .A4(new_n203), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT0), .A4(G128), .ZN(new_n239));
  XNOR2_X1  g053(.A(G143), .B(G146), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT0), .B(G128), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n201), .A2(new_n197), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n200), .B1(new_n199), .B2(new_n246), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n244), .B(G101), .C1(new_n245), .C2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n202), .A2(KEYINPUT4), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n196), .B1(new_n200), .B2(new_n199), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n195), .B1(new_n250), .B2(new_n194), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n243), .B(new_n248), .C1(new_n249), .C2(new_n251), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n237), .A2(new_n232), .A3(new_n238), .A4(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(G110), .B(G140), .ZN(new_n254));
  INV_X1    g068(.A(G953), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G227), .ZN(new_n256));
  XOR2_X1   g070(.A(new_n254), .B(new_n256), .Z(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT12), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n219), .A2(new_n259), .A3(new_n233), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n235), .A2(new_n253), .A3(new_n258), .A4(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n215), .A2(new_n217), .A3(new_n236), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n252), .A2(new_n238), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n233), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n258), .B1(new_n265), .B2(new_n253), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n187), .B(new_n188), .C1(new_n262), .C2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n187), .A2(new_n188), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n235), .A2(new_n253), .A3(new_n260), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n257), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n265), .A2(new_n253), .A3(new_n258), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n267), .B(new_n269), .C1(new_n187), .C2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(G214), .B1(G237), .B2(G902), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n275), .B(KEYINPUT78), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT9), .B(G234), .ZN(new_n278));
  OAI21_X1  g092(.A(G221), .B1(new_n278), .B2(G902), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n274), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(G110), .B(G122), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G113), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT2), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT2), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G113), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(G116), .B(G119), .ZN(new_n288));
  OR2_X1    g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n288), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n291), .B(new_n248), .C1(new_n249), .C2(new_n251), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT79), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G116), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(G119), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT5), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n283), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G119), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G116), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n295), .A2(G119), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT5), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n298), .A2(new_n302), .B1(new_n288), .B2(new_n287), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n202), .A3(new_n203), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n304), .B1(new_n292), .B2(KEYINPUT79), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n282), .B1(new_n294), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n251), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(KEYINPUT4), .A3(new_n202), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT79), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n308), .A2(new_n309), .A3(new_n291), .A4(new_n248), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n310), .A2(new_n293), .A3(new_n281), .A4(new_n304), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n306), .A2(KEYINPUT6), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G224), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(G953), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n242), .A2(G125), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(G125), .B1(new_n211), .B2(new_n213), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n314), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n317), .ZN(new_n319));
  INV_X1    g133(.A(new_n314), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(new_n315), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT6), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n323), .B(new_n282), .C1(new_n294), .C2(new_n305), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n312), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT80), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n281), .B(KEYINPUT8), .ZN(new_n327));
  INV_X1    g141(.A(new_n304), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n303), .B1(new_n202), .B2(new_n203), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n319), .A2(new_n315), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n314), .A2(KEYINPUT7), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n332), .B1(new_n318), .B2(new_n321), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n326), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n316), .A2(new_n314), .A3(new_n317), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n320), .B1(new_n319), .B2(new_n315), .ZN(new_n338));
  OAI22_X1  g152(.A1(new_n337), .A2(new_n338), .B1(KEYINPUT7), .B2(new_n314), .ZN(new_n339));
  INV_X1    g153(.A(new_n303), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n204), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n304), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n342), .A2(new_n327), .B1(new_n331), .B2(new_n332), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n339), .A2(new_n343), .A3(KEYINPUT80), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n336), .A2(new_n344), .A3(new_n311), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n325), .A2(new_n188), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(G210), .B1(G237), .B2(G902), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(KEYINPUT81), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT81), .B1(new_n346), .B2(new_n348), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n325), .A2(new_n188), .A3(new_n345), .A4(new_n347), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT82), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n345), .A2(new_n188), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n356), .A2(KEYINPUT82), .A3(new_n325), .A4(new_n347), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n280), .B1(new_n352), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G475), .ZN(new_n360));
  AND3_X1   g174(.A1(KEYINPUT70), .A2(G125), .A3(G140), .ZN(new_n361));
  AOI21_X1  g175(.A(G140), .B1(KEYINPUT70), .B2(G125), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT16), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G140), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G125), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n363), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(G146), .B1(new_n364), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(KEYINPUT70), .A2(G125), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n365), .ZN(new_n371));
  NAND3_X1  g185(.A1(KEYINPUT70), .A2(G125), .A3(G140), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(KEYINPUT16), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n205), .A3(new_n367), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G237), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT66), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT66), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G237), .ZN(new_n381));
  AOI21_X1  g195(.A(G953), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(G143), .A3(G214), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(G143), .B1(new_n382), .B2(G214), .ZN(new_n385));
  OAI211_X1 g199(.A(KEYINPUT17), .B(G131), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n369), .A2(KEYINPUT87), .A3(new_n374), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n377), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(G131), .B1(new_n384), .B2(new_n385), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT17), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n380), .A2(G237), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n378), .A2(KEYINPUT66), .ZN(new_n392));
  OAI211_X1 g206(.A(G214), .B(new_n255), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n207), .ZN(new_n394));
  INV_X1    g208(.A(G131), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(new_n383), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n389), .A2(new_n390), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G125), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G140), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n366), .A2(new_n399), .A3(new_n205), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT71), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT71), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n366), .A2(new_n399), .A3(new_n402), .A4(new_n205), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n371), .A2(G146), .A3(new_n372), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n394), .A2(KEYINPUT83), .A3(new_n383), .ZN(new_n407));
  NAND2_X1  g221(.A1(KEYINPUT18), .A2(G131), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n408), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n394), .A2(KEYINPUT83), .A3(new_n383), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n388), .A2(new_n397), .B1(new_n406), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(G113), .B(G122), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(new_n198), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n413), .B(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n360), .B1(new_n416), .B2(new_n188), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n295), .A2(G122), .ZN(new_n419));
  INV_X1    g233(.A(G122), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n420), .A2(G116), .ZN(new_n421));
  OR3_X1    g235(.A1(new_n419), .A2(new_n421), .A3(G107), .ZN(new_n422));
  OAI21_X1  g236(.A(G107), .B1(new_n419), .B2(new_n421), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n207), .A2(G128), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT13), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n212), .A2(G143), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n425), .A2(new_n426), .ZN(new_n430));
  OAI21_X1  g244(.A(G134), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n226), .A2(new_n228), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n425), .A2(new_n428), .ZN(new_n433));
  OR2_X1    g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n424), .A2(new_n431), .A3(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n432), .B(new_n433), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n422), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT88), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT14), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n438), .B1(new_n421), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(KEYINPUT88), .B(KEYINPUT14), .C1(new_n420), .C2(G116), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n419), .B1(new_n439), .B2(new_n421), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n191), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n435), .B1(new_n437), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G217), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n278), .A2(new_n446), .A3(G953), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n435), .B(new_n447), .C1(new_n437), .C2(new_n444), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n188), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT89), .ZN(new_n453));
  AOI21_X1  g267(.A(G902), .B1(new_n449), .B2(new_n450), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT89), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT15), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n453), .A2(new_n456), .B1(new_n457), .B2(G478), .ZN(new_n458));
  AOI211_X1 g272(.A(KEYINPUT89), .B(G902), .C1(new_n449), .C2(new_n450), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(G478), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G952), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(G953), .ZN(new_n463));
  NAND2_X1  g277(.A1(G234), .A2(G237), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT21), .B(G898), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n464), .A2(G902), .A3(G953), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  XOR2_X1   g283(.A(new_n469), .B(KEYINPUT90), .Z(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n458), .A2(new_n461), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT20), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n394), .A2(new_n395), .A3(new_n383), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n395), .B1(new_n394), .B2(new_n383), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT84), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT84), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n389), .A2(new_n477), .A3(new_n396), .ZN(new_n478));
  INV_X1    g292(.A(new_n369), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n371), .A2(KEYINPUT19), .A3(new_n372), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n366), .A2(new_n399), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n480), .B(KEYINPUT85), .C1(KEYINPUT19), .C2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(KEYINPUT85), .B2(new_n480), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n479), .B1(new_n483), .B2(new_n205), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n476), .A2(new_n478), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n412), .A2(new_n406), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n415), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n487), .A2(KEYINPUT86), .B1(new_n413), .B2(new_n415), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n486), .ZN(new_n489));
  INV_X1    g303(.A(new_n415), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT86), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(G475), .A2(G902), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n473), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n495), .ZN(new_n497));
  AOI211_X1 g311(.A(KEYINPUT20), .B(new_n497), .C1(new_n488), .C2(new_n493), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n418), .B(new_n472), .C1(new_n496), .C2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT91), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n489), .A2(KEYINPUT86), .A3(new_n490), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n413), .A2(new_n415), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n487), .A2(KEYINPUT86), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n495), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT20), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n494), .A2(new_n473), .A3(new_n495), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n417), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(KEYINPUT91), .A3(new_n472), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n501), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n446), .B1(G234), .B2(new_n188), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT23), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n299), .B2(G128), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n212), .A2(KEYINPUT23), .A3(G119), .ZN(new_n515));
  INV_X1    g329(.A(G110), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n299), .A2(G128), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n514), .A2(new_n515), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(G119), .B(G128), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n516), .A2(KEYINPUT24), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT24), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(G110), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n518), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n369), .A2(new_n404), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT72), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n212), .A2(G119), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n517), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT24), .B(G110), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT69), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G110), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT69), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n523), .A2(new_n519), .A3(new_n534), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n531), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n375), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n369), .A2(new_n404), .A3(new_n524), .A4(KEYINPUT72), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n527), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT73), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n527), .A2(new_n537), .A3(KEYINPUT73), .A4(new_n538), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT22), .B(G137), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n255), .A2(G221), .A3(G234), .ZN(new_n544));
  XOR2_X1   g358(.A(new_n543), .B(new_n544), .Z(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n541), .A2(new_n542), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n539), .A2(new_n540), .A3(new_n545), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT25), .B1(new_n549), .B2(new_n188), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT25), .ZN(new_n551));
  AOI211_X1 g365(.A(new_n551), .B(G902), .C1(new_n547), .C2(new_n548), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n512), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n512), .A2(G902), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT74), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n549), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n243), .B1(new_n230), .B2(new_n231), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT30), .ZN(new_n560));
  AOI21_X1  g374(.A(G137), .B1(new_n226), .B2(new_n228), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n220), .A2(G134), .ZN(new_n562));
  OAI21_X1  g376(.A(G131), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n229), .A2(new_n395), .A3(new_n223), .A4(new_n221), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n563), .A2(new_n564), .A3(new_n213), .A4(new_n211), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n559), .A2(new_n560), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n560), .B1(new_n559), .B2(new_n565), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n291), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT26), .B(G101), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n382), .A2(G210), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n569), .B1(new_n382), .B2(G210), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n291), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n559), .A2(new_n576), .A3(new_n565), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n568), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT31), .ZN(new_n579));
  AND4_X1   g393(.A1(new_n563), .A2(new_n564), .A3(new_n213), .A4(new_n211), .ZN(new_n580));
  INV_X1    g394(.A(new_n225), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n221), .A2(new_n223), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n224), .A2(new_n225), .A3(new_n229), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n242), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n580), .A2(new_n586), .A3(new_n291), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT30), .B1(new_n580), .B2(new_n586), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n559), .A2(new_n560), .A3(new_n565), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n587), .B1(new_n590), .B2(new_n291), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT31), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n592), .A3(new_n575), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n576), .B1(new_n559), .B2(new_n565), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT28), .B1(new_n587), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT28), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n577), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n574), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n579), .A2(new_n593), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(G472), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n601), .A3(new_n188), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT32), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT32), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n600), .A2(new_n604), .A3(new_n601), .A4(new_n188), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n595), .A2(new_n575), .A3(new_n597), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n576), .B1(new_n588), .B2(new_n589), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n574), .B1(new_n608), .B2(new_n587), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT29), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n607), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n188), .B1(new_n607), .B2(new_n610), .ZN(new_n612));
  OAI21_X1  g426(.A(G472), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT68), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT68), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n615), .B(G472), .C1(new_n611), .C2(new_n612), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n558), .B1(new_n606), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n359), .A2(new_n511), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT92), .B(G101), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G3));
  INV_X1    g435(.A(KEYINPUT94), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n451), .B(KEYINPUT33), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(G478), .A3(new_n188), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT93), .B(G478), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n452), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n622), .B1(new_n509), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n418), .B1(new_n496), .B2(new_n498), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(KEYINPUT94), .A3(new_n627), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n346), .A2(new_n348), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n353), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n275), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n471), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n274), .A2(new_n279), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n600), .A2(new_n188), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(G472), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n639), .A2(new_n557), .A3(new_n553), .A4(new_n602), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n632), .A2(new_n636), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  INV_X1    g458(.A(KEYINPUT95), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n645), .B1(new_n496), .B2(new_n498), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT95), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n454), .A2(new_n455), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n460), .B1(new_n648), .B2(new_n459), .ZN(new_n649));
  INV_X1    g463(.A(new_n461), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n417), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n646), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n636), .A2(new_n652), .A3(new_n641), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  INV_X1    g469(.A(KEYINPUT97), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT96), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n546), .A2(KEYINPUT36), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n539), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n556), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n553), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n657), .B1(new_n553), .B2(new_n660), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n656), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n553), .A2(new_n660), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT96), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n553), .A2(new_n657), .A3(new_n660), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n665), .A2(KEYINPUT97), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n600), .A2(new_n601), .A3(new_n188), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n601), .B1(new_n600), .B2(new_n188), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n668), .A2(new_n359), .A3(new_n511), .A4(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT37), .B(G110), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  OR2_X1    g488(.A1(new_n468), .A2(G900), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n465), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n652), .A2(KEYINPUT98), .A3(new_n676), .ZN(new_n677));
  AOI22_X1  g491(.A1(new_n603), .A2(new_n605), .B1(new_n614), .B2(new_n616), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n678), .A2(new_n635), .A3(new_n637), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n646), .A2(new_n647), .A3(new_n651), .A4(new_n676), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT98), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n677), .A2(new_n679), .A3(new_n668), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G128), .ZN(G30));
  NAND2_X1  g498(.A1(new_n352), .A2(new_n358), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n676), .B(KEYINPUT39), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n274), .A2(new_n279), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT40), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n650), .A2(new_n649), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n630), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n661), .A2(new_n662), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n591), .A2(new_n574), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n587), .A2(new_n594), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n188), .B1(new_n696), .B2(new_n575), .ZN(new_n697));
  OAI21_X1  g511(.A(G472), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n606), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n693), .A2(new_n275), .A3(new_n694), .A4(new_n699), .ZN(new_n700));
  OR3_X1    g514(.A1(new_n687), .A2(new_n690), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G143), .ZN(G45));
  INV_X1    g516(.A(KEYINPUT100), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n630), .A2(new_n627), .A3(new_n676), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n703), .B1(new_n704), .B2(new_n635), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n509), .A2(new_n628), .ZN(new_n706));
  INV_X1    g520(.A(new_n275), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n707), .B1(new_n633), .B2(new_n353), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n706), .A2(KEYINPUT100), .A3(new_n708), .A4(new_n676), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n678), .A2(new_n637), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n705), .A2(new_n668), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G146), .ZN(G48));
  INV_X1    g526(.A(new_n266), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n261), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n188), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(G469), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n279), .A3(new_n267), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n678), .A2(new_n558), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n636), .A3(new_n632), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  NAND3_X1  g535(.A1(new_n718), .A2(new_n636), .A3(new_n652), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  INV_X1    g537(.A(new_n678), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n635), .A2(new_n717), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n668), .A2(new_n724), .A3(new_n511), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT101), .B(G119), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G21));
  INV_X1    g542(.A(KEYINPUT102), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n592), .B1(new_n591), .B2(new_n575), .ZN(new_n730));
  NOR4_X1   g544(.A1(new_n608), .A2(KEYINPUT31), .A3(new_n574), .A4(new_n587), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n575), .B1(new_n595), .B2(new_n597), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n729), .B1(new_n733), .B2(G902), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n734), .B1(new_n669), .B2(new_n670), .ZN(new_n735));
  INV_X1    g549(.A(new_n558), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n638), .A2(new_n729), .A3(new_n601), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT103), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n735), .A2(new_n736), .A3(KEYINPUT103), .A4(new_n737), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR4_X1   g556(.A1(new_n692), .A2(new_n635), .A3(new_n471), .A4(new_n717), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT104), .B(G122), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G24));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n704), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n630), .A2(KEYINPUT105), .A3(new_n627), .A4(new_n676), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n735), .A2(new_n737), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n694), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n750), .A2(KEYINPUT106), .A3(new_n725), .A4(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n752), .A2(new_n725), .A3(new_n748), .A4(new_n749), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT106), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G125), .ZN(G27));
  INV_X1    g572(.A(new_n279), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT107), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n760), .B1(new_n271), .B2(new_n272), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n272), .A2(new_n760), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n761), .A2(new_n187), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n267), .A2(new_n269), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT108), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n273), .A2(KEYINPUT107), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(G469), .A3(new_n762), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n769));
  AOI21_X1  g583(.A(G902), .B1(new_n713), .B2(new_n261), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n268), .B1(new_n770), .B2(new_n187), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n759), .B1(new_n766), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT81), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n633), .A2(new_n774), .ZN(new_n775));
  AND4_X1   g589(.A1(new_n358), .A2(new_n775), .A3(new_n349), .A4(new_n275), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n773), .A2(new_n776), .A3(new_n618), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n750), .A3(KEYINPUT42), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT42), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n773), .A2(new_n776), .A3(new_n618), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n748), .A2(new_n749), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G131), .ZN(G33));
  XNOR2_X1  g598(.A(new_n680), .B(KEYINPUT98), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n777), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G134), .ZN(G36));
  INV_X1    g601(.A(KEYINPUT110), .ZN(new_n788));
  OR3_X1    g602(.A1(new_n630), .A2(KEYINPUT43), .A3(new_n628), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n509), .A2(new_n627), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT43), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT109), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n694), .A2(new_n793), .A3(new_n671), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n793), .B1(new_n694), .B2(new_n671), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n792), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n788), .B1(new_n797), .B2(KEYINPUT44), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n767), .A2(KEYINPUT45), .A3(new_n762), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT45), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n187), .B1(new_n273), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n268), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n802), .A2(KEYINPUT46), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n267), .B1(new_n802), .B2(KEYINPUT46), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n279), .A3(new_n688), .ZN(new_n806));
  INV_X1    g620(.A(new_n776), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT44), .ZN(new_n809));
  INV_X1    g623(.A(new_n796), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n794), .ZN(new_n811));
  OAI211_X1 g625(.A(KEYINPUT110), .B(new_n809), .C1(new_n811), .C2(new_n792), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n797), .A2(KEYINPUT44), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n798), .A2(new_n808), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G137), .ZN(G39));
  NOR3_X1   g629(.A1(new_n724), .A2(new_n736), .A3(new_n704), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n805), .A2(KEYINPUT47), .A3(new_n279), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT47), .B1(new_n805), .B2(new_n279), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n776), .B(new_n816), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G140), .ZN(G42));
  NAND2_X1  g634(.A1(new_n462), .A2(new_n255), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT117), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n717), .A2(new_n275), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n687), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n792), .A2(new_n465), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n742), .ZN(new_n826));
  OR4_X1    g640(.A1(KEYINPUT116), .A2(new_n824), .A3(new_n826), .A4(KEYINPUT50), .ZN(new_n827));
  INV_X1    g641(.A(new_n716), .ZN(new_n828));
  INV_X1    g642(.A(new_n267), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n776), .A2(new_n279), .A3(new_n830), .ZN(new_n831));
  NOR4_X1   g645(.A1(new_n831), .A2(new_n558), .A3(new_n465), .A4(new_n699), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n630), .A2(new_n627), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n831), .A2(new_n792), .A3(new_n465), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n832), .A2(new_n833), .B1(new_n834), .B2(new_n752), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n827), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n817), .A2(new_n818), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n830), .A2(new_n759), .ZN(new_n838));
  AOI211_X1 g652(.A(new_n807), .B(new_n826), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  XOR2_X1   g654(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n841));
  OAI21_X1  g655(.A(new_n841), .B1(new_n824), .B2(new_n826), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n836), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT51), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n836), .A2(new_n840), .A3(KEYINPUT51), .A4(new_n842), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n832), .A2(new_n632), .ZN(new_n847));
  INV_X1    g661(.A(new_n725), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n847), .B(new_n463), .C1(new_n848), .C2(new_n826), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n834), .A2(new_n618), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n850), .A2(KEYINPUT48), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(KEYINPUT48), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n849), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n845), .A2(new_n846), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n754), .B(KEYINPUT106), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n692), .A2(new_n635), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n676), .B(KEYINPUT113), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n553), .A2(new_n660), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT114), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n857), .A2(new_n773), .A3(new_n860), .A4(new_n699), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n683), .A2(new_n711), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n855), .B1(new_n856), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n862), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n757), .A3(KEYINPUT52), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n752), .A2(new_n748), .A3(new_n749), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n773), .A2(new_n776), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n867), .A2(new_n868), .B1(new_n785), .B2(new_n777), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n630), .A2(new_n627), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n691), .A2(KEYINPUT111), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT111), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n650), .A2(new_n649), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n509), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n471), .A2(new_n276), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n876), .A2(new_n685), .A3(new_n641), .A4(new_n877), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n672), .A2(new_n619), .A3(new_n878), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n646), .A2(new_n647), .ZN(new_n880));
  INV_X1    g694(.A(new_n676), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n874), .A2(new_n417), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n776), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT112), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n668), .A2(new_n710), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n776), .A2(KEYINPUT112), .A3(new_n880), .A4(new_n882), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n869), .A2(new_n879), .A3(new_n888), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n718), .B(new_n636), .C1(new_n632), .C2(new_n652), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n744), .A2(new_n890), .A3(new_n726), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n783), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n866), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT53), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n683), .A2(new_n711), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n756), .B2(new_n753), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n861), .A2(KEYINPUT52), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n863), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT115), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n869), .A2(new_n879), .A3(new_n903), .A4(new_n888), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n619), .A2(new_n878), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n750), .A2(new_n868), .A3(new_n752), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n905), .A2(new_n906), .A3(new_n786), .A4(new_n672), .ZN(new_n907));
  INV_X1    g721(.A(new_n888), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT115), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n891), .A2(new_n783), .A3(KEYINPUT53), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n902), .A2(new_n904), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n896), .A2(new_n897), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n894), .A2(KEYINPUT53), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n902), .A2(new_n895), .A3(new_n893), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n912), .B1(new_n915), .B2(new_n897), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n822), .B1(new_n854), .B2(new_n916), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n830), .B(KEYINPUT49), .Z(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(new_n790), .ZN(new_n919));
  NOR4_X1   g733(.A1(new_n699), .A2(new_n558), .A3(new_n276), .A4(new_n759), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n919), .A2(new_n687), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n917), .A2(new_n921), .ZN(G75));
  NAND3_X1  g736(.A1(new_n909), .A2(new_n910), .A3(new_n904), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n864), .A2(new_n757), .ZN(new_n924));
  AOI22_X1  g738(.A1(new_n924), .A2(new_n855), .B1(new_n899), .B2(new_n900), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT53), .B1(new_n866), .B2(new_n893), .ZN(new_n927));
  OAI211_X1 g741(.A(G210), .B(G902), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n312), .A2(new_n324), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(new_n322), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT55), .ZN(new_n931));
  NOR2_X1   g745(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n932));
  AND2_X1   g746(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n928), .B(new_n931), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n255), .A2(G952), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT118), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n188), .B1(new_n896), .B2(new_n911), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT56), .B1(new_n939), .B2(G210), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n938), .B1(new_n940), .B2(new_n931), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT56), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n931), .B1(new_n928), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(KEYINPUT118), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n937), .B1(new_n941), .B2(new_n944), .ZN(G51));
  XNOR2_X1  g759(.A(new_n268), .B(KEYINPUT57), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n926), .A2(new_n927), .A3(KEYINPUT54), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n897), .B1(new_n896), .B2(new_n911), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n714), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n939), .A2(new_n799), .A3(new_n801), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n935), .B1(new_n950), .B2(new_n951), .ZN(G54));
  NAND2_X1  g766(.A1(KEYINPUT58), .A2(G475), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n939), .A2(new_n494), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n494), .B1(new_n939), .B2(new_n954), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n955), .A2(new_n956), .A3(new_n935), .ZN(G60));
  NAND2_X1  g771(.A1(G478), .A2(G902), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT59), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n623), .B1(new_n916), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n623), .A2(new_n959), .ZN(new_n961));
  INV_X1    g775(.A(new_n948), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n961), .B1(new_n962), .B2(new_n912), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n960), .A2(new_n963), .A3(new_n935), .ZN(G63));
  NAND2_X1  g778(.A1(G217), .A2(G902), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT121), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT60), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n926), .B2(new_n927), .ZN(new_n968));
  INV_X1    g782(.A(new_n549), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n935), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n896), .A2(new_n911), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT122), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n971), .A2(new_n972), .A3(new_n659), .A4(new_n967), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n659), .B(new_n967), .C1(new_n926), .C2(new_n927), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(KEYINPUT122), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n970), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  XNOR2_X1  g790(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n970), .A2(KEYINPUT61), .A3(new_n974), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(G66));
  OAI21_X1  g794(.A(G953), .B1(new_n466), .B2(new_n313), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n891), .A2(new_n879), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n981), .B1(new_n983), .B2(G953), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n929), .B1(G898), .B2(new_n255), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n984), .B(new_n985), .ZN(G69));
  XNOR2_X1  g800(.A(new_n590), .B(new_n483), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT124), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n899), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(KEYINPUT124), .B1(new_n856), .B2(new_n898), .ZN(new_n990));
  AND4_X1   g804(.A1(new_n814), .A2(new_n989), .A3(new_n990), .A4(new_n819), .ZN(new_n991));
  INV_X1    g805(.A(new_n618), .ZN(new_n992));
  NOR4_X1   g806(.A1(new_n806), .A2(new_n992), .A3(new_n635), .A4(new_n692), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n783), .A2(new_n786), .ZN(new_n994));
  OR2_X1    g808(.A1(new_n994), .A2(KEYINPUT126), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(KEYINPUT126), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n993), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(G953), .B1(new_n991), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n255), .A2(G900), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT125), .Z(new_n1000));
  OAI21_X1  g814(.A(new_n987), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n987), .B(KEYINPUT123), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n992), .A2(new_n689), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1003), .A2(new_n776), .A3(new_n876), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n814), .A2(new_n819), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n989), .A2(new_n990), .A3(new_n701), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT62), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n989), .A2(new_n990), .A3(KEYINPUT62), .A4(new_n701), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1005), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1002), .B1(new_n1010), .B2(G953), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n255), .B1(G227), .B2(G900), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n1001), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1012), .B1(new_n1001), .B2(new_n1011), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1013), .A2(new_n1014), .ZN(G72));
  NAND3_X1  g829(.A1(new_n991), .A2(new_n997), .A3(new_n983), .ZN(new_n1016));
  NAND2_X1  g830(.A1(G472), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT63), .Z(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1019), .A2(new_n574), .A3(new_n591), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n609), .B(KEYINPUT127), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(new_n578), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(new_n1018), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n1020), .B(new_n936), .C1(new_n915), .C2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1010), .A2(new_n983), .ZN(new_n1025));
  AOI211_X1 g839(.A(new_n574), .B(new_n591), .C1(new_n1025), .C2(new_n1018), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1024), .A2(new_n1026), .ZN(G57));
endmodule


