//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  INV_X1    g000(.A(KEYINPUT31), .ZN(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n189), .B(KEYINPUT27), .Z(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(G101), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT11), .A3(G134), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G137), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  OAI211_X1 g012(.A(KEYINPUT64), .B(new_n198), .C1(new_n195), .C2(G137), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n193), .A2(G134), .ZN(new_n201));
  AOI21_X1  g015(.A(KEYINPUT64), .B1(new_n201), .B2(new_n198), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n197), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G131), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n194), .A2(new_n196), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n198), .B1(new_n195), .B2(G137), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n205), .B1(new_n208), .B2(new_n199), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n204), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT0), .A2(G128), .ZN(new_n218));
  OR2_X1    g032(.A1(KEYINPUT0), .A2(G128), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(G143), .B(G146), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(KEYINPUT0), .A3(G128), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n225), .A3(G128), .ZN(new_n226));
  INV_X1    g040(.A(G128), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n227), .B1(new_n214), .B2(KEYINPUT1), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n229));
  NOR3_X1   g043(.A1(new_n228), .A2(new_n221), .A3(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT1), .B1(new_n215), .B2(G146), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G128), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT65), .B1(new_n232), .B2(new_n217), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n226), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n210), .B1(new_n196), .B2(new_n201), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n235), .B1(new_n209), .B2(new_n210), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n212), .A2(new_n224), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  OR2_X1    g051(.A1(KEYINPUT67), .A2(G119), .ZN(new_n238));
  NAND2_X1  g052(.A1(KEYINPUT67), .A2(G119), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(G116), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G116), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G119), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT2), .B(G113), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n240), .A2(new_n242), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n244), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n192), .B1(new_n237), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n250), .B1(new_n237), .B2(KEYINPUT30), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n234), .A2(new_n236), .ZN(new_n253));
  AOI211_X1 g067(.A(G131), .B(new_n205), .C1(new_n208), .C2(new_n199), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n208), .A2(new_n199), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n210), .B1(new_n255), .B2(new_n197), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n224), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT30), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT66), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n261));
  AOI211_X1 g075(.A(new_n261), .B(KEYINPUT30), .C1(new_n253), .C2(new_n257), .ZN(new_n262));
  OAI211_X1 g076(.A(KEYINPUT68), .B(new_n252), .C1(new_n260), .C2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n261), .B1(new_n237), .B2(KEYINPUT30), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n258), .A2(KEYINPUT66), .A3(new_n259), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT68), .B1(new_n267), .B2(new_n252), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n187), .B(new_n251), .C1(new_n264), .C2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT70), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n252), .B1(new_n260), .B2(new_n262), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n263), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n274), .A2(new_n275), .A3(new_n187), .A4(new_n251), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n251), .B1(new_n264), .B2(new_n268), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT69), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n274), .A2(new_n280), .A3(new_n251), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(KEYINPUT31), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n192), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n237), .A2(new_n250), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n258), .A2(new_n249), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT28), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT28), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n283), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n277), .A2(new_n282), .A3(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(G472), .A2(G902), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT32), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n274), .A2(new_n284), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n192), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n287), .A2(new_n283), .A3(new_n289), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n300), .A2(KEYINPUT29), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(G902), .B1(new_n300), .B2(KEYINPUT29), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G472), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n297), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n292), .A2(new_n293), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT71), .B(KEYINPUT32), .Z(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n307), .A2(KEYINPUT72), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT72), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n290), .B1(new_n270), .B2(new_n276), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n294), .B1(new_n312), .B2(new_n282), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n311), .B1(new_n313), .B2(new_n308), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n306), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G217), .ZN(new_n316));
  INV_X1    g130(.A(G902), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n316), .B1(G234), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n320));
  XOR2_X1   g134(.A(KEYINPUT67), .B(G119), .Z(new_n321));
  OAI21_X1  g135(.A(new_n320), .B1(new_n321), .B2(G128), .ZN(new_n322));
  OR2_X1    g136(.A1(G119), .A2(G128), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n321), .B2(new_n227), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n322), .B1(new_n324), .B2(new_n320), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT24), .B(G110), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  OAI22_X1  g141(.A1(new_n325), .A2(G110), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT16), .ZN(new_n329));
  INV_X1    g143(.A(G140), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(G125), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(G125), .ZN(new_n332));
  INV_X1    g146(.A(G125), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G140), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n331), .B1(new_n335), .B2(new_n329), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(new_n213), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n332), .A2(new_n334), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n337), .B1(new_n213), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n328), .A2(new_n339), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n336), .A2(new_n213), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n213), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n341), .A2(new_n342), .B1(new_n324), .B2(new_n327), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n325), .A2(G110), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT73), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT73), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n340), .A2(new_n345), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT22), .B(G137), .ZN(new_n351));
  INV_X1    g165(.A(G953), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n352), .A2(G221), .A3(G234), .ZN(new_n353));
  XOR2_X1   g167(.A(new_n351), .B(new_n353), .Z(new_n354));
  NAND2_X1  g168(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n354), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n355), .A2(new_n317), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT25), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n357), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(new_n350), .B2(new_n354), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(KEYINPUT25), .A3(new_n317), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n319), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n318), .A2(G902), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n366), .B(KEYINPUT74), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n315), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(G214), .B1(G237), .B2(G902), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(KEYINPUT81), .ZN(new_n373));
  INV_X1    g187(.A(G104), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(G107), .ZN(new_n375));
  AND2_X1   g189(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n376));
  NOR2_X1   g190(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI22_X1  g192(.A1(new_n374), .A2(G107), .B1(KEYINPUT75), .B2(KEYINPUT3), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n374), .A2(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G101), .ZN(new_n382));
  INV_X1    g196(.A(G101), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n378), .A2(new_n383), .A3(new_n379), .A4(new_n380), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(KEYINPUT4), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n381), .A2(new_n386), .A3(G101), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n249), .A3(new_n387), .ZN(new_n388));
  XOR2_X1   g202(.A(KEYINPUT82), .B(KEYINPUT5), .Z(new_n389));
  NAND4_X1  g203(.A1(new_n321), .A2(new_n389), .A3(KEYINPUT83), .A4(G116), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT83), .ZN(new_n391));
  XNOR2_X1  g205(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n391), .B1(new_n240), .B2(new_n392), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(G113), .B1(new_n247), .B2(new_n389), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n246), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT77), .ZN(new_n397));
  INV_X1    g211(.A(G107), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(G104), .ZN(new_n399));
  OAI21_X1  g213(.A(G101), .B1(new_n375), .B2(new_n399), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n384), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n397), .B1(new_n384), .B2(new_n400), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n388), .B1(new_n396), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G110), .B(G122), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n405), .B(new_n388), .C1(new_n396), .C2(new_n403), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(KEYINPUT6), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(KEYINPUT84), .B1(new_n223), .B2(G125), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n229), .B1(new_n228), .B2(new_n221), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n232), .A2(KEYINPUT65), .A3(new_n217), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(new_n333), .A3(new_n226), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n223), .A2(KEYINPUT84), .A3(G125), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n411), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n352), .A2(G224), .ZN(new_n418));
  XOR2_X1   g232(.A(new_n417), .B(new_n418), .Z(new_n419));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n404), .A2(new_n420), .A3(new_n406), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n409), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  XOR2_X1   g236(.A(new_n405), .B(KEYINPUT8), .Z(new_n423));
  INV_X1    g237(.A(G113), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n424), .B1(new_n243), .B2(new_n392), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n390), .A2(new_n393), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n425), .A2(new_n426), .B1(new_n243), .B2(new_n245), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n384), .A2(new_n400), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n423), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n243), .A2(KEYINPUT5), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n426), .A2(new_n430), .A3(G113), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n246), .ZN(new_n432));
  INV_X1    g246(.A(new_n428), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n418), .A2(KEYINPUT7), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n429), .A2(new_n434), .B1(new_n417), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(KEYINPUT7), .B1(new_n418), .B2(KEYINPUT85), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n437), .B1(KEYINPUT85), .B2(new_n418), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n411), .A2(new_n415), .A3(new_n416), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT86), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT84), .ZN(new_n441));
  AOI211_X1 g255(.A(new_n441), .B(new_n333), .C1(new_n220), .C2(new_n222), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n410), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT86), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n443), .A2(new_n444), .A3(new_n415), .A4(new_n438), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT87), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n436), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n408), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n447), .B1(new_n436), .B2(new_n446), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n317), .B(new_n422), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G210), .B1(G237), .B2(G902), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n436), .A2(new_n446), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT87), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(new_n408), .A3(new_n448), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n457), .A2(new_n317), .A3(new_n452), .A4(new_n422), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n373), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G952), .ZN(new_n460));
  AOI211_X1 g274(.A(G953), .B(new_n460), .C1(G234), .C2(G237), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT21), .B(G898), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT95), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI211_X1 g278(.A(new_n317), .B(new_n352), .C1(G234), .C2(G237), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(G113), .B(G122), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(new_n374), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT90), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n338), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n335), .A2(KEYINPUT90), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(G146), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n338), .A2(new_n213), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n188), .A2(G214), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n215), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(KEYINPUT18), .A2(G131), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI211_X1 g296(.A(KEYINPUT89), .B(new_n481), .C1(new_n477), .C2(new_n478), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT89), .ZN(new_n484));
  INV_X1    g298(.A(new_n481), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n484), .B1(new_n479), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n475), .B(new_n482), .C1(new_n483), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n479), .A2(G131), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT17), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n477), .A2(new_n210), .A3(new_n478), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n479), .A2(KEYINPUT17), .A3(G131), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n491), .A2(new_n342), .A3(new_n341), .A4(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n469), .B1(new_n487), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(G902), .B1(new_n494), .B2(KEYINPUT92), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n487), .A2(new_n493), .A3(new_n469), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT92), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n495), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n499), .A2(G475), .ZN(new_n500));
  INV_X1    g314(.A(new_n496), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n337), .B1(new_n488), .B2(new_n490), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n471), .A2(KEYINPUT19), .A3(new_n472), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n503), .B(new_n213), .C1(KEYINPUT19), .C2(new_n335), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n469), .B1(new_n505), .B2(new_n487), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT91), .B1(new_n501), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT91), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n505), .A2(new_n487), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n508), .B(new_n496), .C1(new_n509), .C2(new_n469), .ZN(new_n510));
  NOR2_X1   g324(.A1(G475), .A2(G902), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n507), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT20), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n516), .B(new_n511), .C1(new_n501), .C2(new_n506), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n500), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(G128), .B(G143), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n195), .ZN(new_n520));
  XNOR2_X1  g334(.A(G116), .B(G122), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n522), .A2(G107), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n521), .A2(new_n398), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n520), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT13), .B1(new_n215), .B2(G128), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n526), .A2(KEYINPUT93), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n227), .A2(G143), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(KEYINPUT93), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT94), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT94), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n527), .A2(new_n532), .A3(new_n528), .A4(new_n529), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n215), .A2(KEYINPUT13), .A3(G128), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n525), .B1(new_n535), .B2(G134), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n241), .A2(KEYINPUT14), .A3(G122), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(G107), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT14), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n538), .B1(new_n539), .B2(new_n521), .ZN(new_n540));
  OR2_X1    g354(.A1(new_n519), .A2(new_n195), .ZN(new_n541));
  AOI211_X1 g355(.A(new_n523), .B(new_n540), .C1(new_n520), .C2(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT9), .B(G234), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n543), .A2(new_n316), .A3(G953), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  OR3_X1    g359(.A1(new_n536), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n545), .B1(new_n536), .B2(new_n542), .ZN(new_n547));
  AOI21_X1  g361(.A(G902), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(G478), .ZN(new_n549));
  OR2_X1    g363(.A1(new_n549), .A2(KEYINPUT15), .ZN(new_n550));
  XOR2_X1   g364(.A(new_n548), .B(new_n550), .Z(new_n551));
  NAND4_X1  g365(.A1(new_n459), .A2(new_n467), .A3(new_n518), .A4(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT80), .ZN(new_n553));
  OAI211_X1 g367(.A(KEYINPUT10), .B(new_n234), .C1(new_n401), .C2(new_n402), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT10), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n225), .B1(G143), .B2(new_n213), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT76), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n227), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n231), .A2(KEYINPUT76), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n221), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n226), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n555), .B1(new_n562), .B2(new_n428), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n385), .A2(new_n224), .A3(new_n387), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n254), .A2(new_n256), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n554), .A2(new_n563), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n433), .B1(new_n561), .B2(new_n560), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n428), .A2(new_n414), .A3(new_n226), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(KEYINPUT12), .B1(new_n569), .B2(new_n212), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT12), .ZN(new_n571));
  AOI211_X1 g385(.A(new_n571), .B(new_n565), .C1(new_n567), .C2(new_n568), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n566), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(G110), .B(G140), .ZN(new_n574));
  INV_X1    g388(.A(G227), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(G953), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n574), .B(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n566), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n554), .A2(new_n563), .A3(new_n564), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n212), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n573), .A2(new_n577), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(G469), .B1(new_n583), .B2(G902), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT78), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n570), .A2(new_n572), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT79), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(new_n566), .B2(new_n578), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n580), .A2(new_n588), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n578), .B1(new_n582), .B2(new_n566), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(G469), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(new_n596), .A3(new_n317), .ZN(new_n597));
  OAI211_X1 g411(.A(KEYINPUT78), .B(G469), .C1(new_n583), .C2(G902), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n586), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(G221), .ZN(new_n600));
  INV_X1    g414(.A(new_n543), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n600), .B1(new_n601), .B2(new_n317), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n553), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n599), .A2(new_n553), .A3(new_n603), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n552), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n371), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G101), .ZN(G3));
  AOI21_X1  g423(.A(new_n370), .B1(new_n605), .B2(new_n606), .ZN(new_n610));
  INV_X1    g424(.A(G472), .ZN(new_n611));
  AOI21_X1  g425(.A(G902), .B1(new_n312), .B2(new_n282), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n307), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n546), .A2(new_n547), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n547), .B2(KEYINPUT96), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n546), .B(new_n547), .C1(KEYINPUT96), .C2(new_n617), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(G478), .A3(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n549), .A2(new_n317), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n548), .B2(new_n549), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n518), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n615), .A2(new_n467), .A3(new_n459), .A4(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT34), .B(G104), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  NAND2_X1  g442(.A1(new_n459), .A2(new_n467), .ZN(new_n629));
  AOI21_X1  g443(.A(KEYINPUT97), .B1(new_n512), .B2(new_n514), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n512), .B2(new_n514), .ZN(new_n631));
  INV_X1    g445(.A(new_n512), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n632), .A2(KEYINPUT97), .A3(new_n513), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NOR4_X1   g448(.A1(new_n629), .A2(new_n500), .A3(new_n551), .A4(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n615), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT35), .B(G107), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  NOR2_X1   g452(.A1(new_n356), .A2(KEYINPUT36), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n346), .B(new_n639), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n640), .A2(new_n367), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n364), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n607), .A2(new_n614), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT37), .B(G110), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G12));
  INV_X1    g460(.A(new_n551), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT98), .B(G900), .Z(new_n648));
  AOI21_X1  g462(.A(new_n461), .B1(new_n465), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n500), .A2(new_n649), .ZN(new_n650));
  AND4_X1   g464(.A1(new_n647), .A2(new_n631), .A3(new_n633), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n454), .A2(new_n458), .ZN(new_n652));
  INV_X1    g466(.A(new_n373), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n642), .ZN(new_n655));
  INV_X1    g469(.A(new_n606), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n651), .B(new_n655), .C1(new_n656), .C2(new_n604), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n315), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(new_n227), .ZN(G30));
  NAND2_X1  g473(.A1(new_n286), .A2(new_n192), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n279), .A2(new_n281), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n317), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(G472), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n297), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(KEYINPUT72), .B1(new_n307), .B2(new_n309), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n313), .A2(new_n311), .A3(new_n308), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n652), .B(KEYINPUT38), .Z(new_n669));
  NOR2_X1   g483(.A1(new_n518), .A2(new_n551), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n642), .A2(new_n653), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n673), .A2(KEYINPUT99), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(KEYINPUT99), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n649), .B(KEYINPUT39), .Z(new_n676));
  OAI21_X1  g490(.A(new_n676), .B1(new_n656), .B2(new_n604), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT40), .Z(new_n678));
  NAND3_X1  g492(.A1(new_n674), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT100), .B(G143), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G45));
  NOR3_X1   g495(.A1(new_n518), .A2(new_n624), .A3(new_n649), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n655), .B(new_n682), .C1(new_n656), .C2(new_n604), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n611), .B1(new_n302), .B2(new_n303), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n292), .B2(new_n296), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(new_n666), .B2(new_n667), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  NOR2_X1   g503(.A1(new_n596), .A2(KEYINPUT101), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n593), .B1(new_n590), .B2(new_n591), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n690), .B1(new_n691), .B2(G902), .ZN(new_n692));
  INV_X1    g506(.A(new_n690), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n579), .A2(KEYINPUT79), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n694), .A2(new_n587), .A3(new_n589), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n317), .B(new_n693), .C1(new_n695), .C2(new_n593), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n692), .A2(new_n696), .A3(new_n603), .ZN(new_n697));
  NOR4_X1   g511(.A1(new_n629), .A2(new_n518), .A3(new_n624), .A4(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n371), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G15));
  INV_X1    g515(.A(new_n370), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n692), .A2(new_n696), .A3(new_n603), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n687), .A2(new_n702), .A3(new_n635), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  NAND2_X1  g519(.A1(new_n518), .A2(new_n551), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n466), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n687), .A2(new_n655), .A3(new_n703), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  AND2_X1   g523(.A1(new_n370), .A2(KEYINPUT103), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n370), .A2(KEYINPUT103), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n611), .B1(new_n292), .B2(new_n317), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n293), .B(KEYINPUT102), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n312), .B2(new_n282), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n670), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n629), .A2(new_n718), .A3(new_n697), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n712), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  NAND3_X1  g535(.A1(new_n703), .A2(new_n682), .A3(new_n459), .ZN(new_n722));
  NOR4_X1   g536(.A1(new_n713), .A2(new_n722), .A3(new_n716), .A4(new_n642), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n333), .ZN(G27));
  OAI21_X1  g538(.A(new_n305), .B1(new_n313), .B2(KEYINPUT32), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n292), .A2(KEYINPUT104), .A3(new_n296), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT104), .B1(new_n292), .B2(new_n296), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n710), .A2(new_n711), .ZN(new_n729));
  OAI21_X1  g543(.A(KEYINPUT105), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n726), .A2(new_n727), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n685), .B1(new_n307), .B2(new_n295), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT105), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n734), .A3(new_n712), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n652), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n653), .ZN(new_n738));
  INV_X1    g552(.A(new_n682), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n597), .A2(new_n584), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n603), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT42), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n736), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT42), .B1(new_n371), .B2(new_n742), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G131), .ZN(G33));
  INV_X1    g563(.A(new_n738), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(new_n603), .A3(new_n651), .A4(new_n740), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n315), .A2(new_n370), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n195), .ZN(G36));
  OR2_X1    g567(.A1(new_n583), .A2(KEYINPUT45), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n583), .A2(KEYINPUT45), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(G469), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(G469), .A2(G902), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT46), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n757), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n597), .A3(new_n761), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n762), .A2(new_n603), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n763), .A2(new_n676), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n518), .A2(KEYINPUT43), .A3(new_n621), .A4(new_n623), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT107), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n624), .A2(KEYINPUT106), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n624), .A2(KEYINPUT106), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n515), .A2(new_n517), .ZN(new_n769));
  INV_X1    g583(.A(new_n500), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n767), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n766), .B1(KEYINPUT43), .B2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n773), .A2(KEYINPUT44), .A3(new_n613), .A4(new_n643), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n764), .A2(new_n750), .A3(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(new_n613), .A3(new_n643), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n776), .A2(new_n778), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT108), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n775), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G137), .ZN(G39));
  XOR2_X1   g597(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n763), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n763), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n702), .A2(new_n738), .A3(new_n739), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n315), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G140), .ZN(G42));
  NAND2_X1  g606(.A1(new_n692), .A2(new_n696), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT49), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n771), .A2(new_n624), .A3(new_n602), .A4(new_n373), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n712), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n796), .B(KEYINPUT110), .Z(new_n797));
  AOI21_X1  g611(.A(new_n664), .B1(new_n310), .B2(new_n314), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n793), .A2(KEYINPUT49), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n797), .A2(new_n798), .A3(new_n669), .A4(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n773), .A2(new_n461), .ZN(new_n802));
  NOR4_X1   g616(.A1(new_n802), .A2(new_n713), .A3(new_n729), .A4(new_n716), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n669), .A2(new_n373), .A3(new_n703), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n802), .A2(new_n697), .A3(new_n738), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n713), .A2(new_n642), .A3(new_n716), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n702), .A2(new_n461), .ZN(new_n813));
  NOR4_X1   g627(.A1(new_n668), .A2(new_n697), .A3(new_n738), .A4(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n518), .A3(new_n624), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n809), .A2(new_n812), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n803), .A2(new_n750), .ZN(new_n817));
  XOR2_X1   g631(.A(new_n789), .B(KEYINPUT114), .Z(new_n818));
  NAND3_X1  g632(.A1(new_n692), .A2(new_n602), .A3(new_n696), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n819), .B(KEYINPUT115), .Z(new_n820));
  AOI21_X1  g634(.A(new_n817), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n801), .B1(new_n816), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n803), .A2(new_n459), .A3(new_n703), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(G952), .A3(new_n352), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n625), .B2(new_n814), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n736), .A2(new_n810), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT48), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n789), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n817), .B1(new_n829), .B2(new_n819), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n830), .A2(new_n801), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n822), .B(new_n828), .C1(new_n816), .C2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n643), .A2(new_n741), .A3(new_n649), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n654), .A2(new_n718), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI22_X1  g651(.A1(new_n315), .A2(new_n683), .B1(new_n798), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n722), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n717), .A2(new_n643), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n840), .B1(new_n315), .B2(new_n657), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n834), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n651), .A2(new_n643), .A3(new_n459), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n605), .B2(new_n606), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n723), .B1(new_n687), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n835), .A2(new_n836), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n668), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n845), .A2(KEYINPUT52), .A3(new_n688), .A4(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n842), .A2(KEYINPUT112), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT112), .B1(new_n842), .B2(new_n848), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n771), .A2(new_n624), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n706), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n629), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n610), .A2(new_n614), .A3(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n708), .A2(new_n644), .A3(new_n720), .A4(new_n855), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n687), .B(new_n702), .C1(new_n698), .C2(new_n607), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n704), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n811), .A2(new_n742), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n551), .A2(new_n650), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n642), .A2(new_n634), .A3(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n750), .B(new_n862), .C1(new_n656), .C2(new_n604), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n860), .B1(new_n863), .B2(new_n315), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n752), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n748), .A2(new_n859), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n833), .B1(new_n851), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n743), .B1(new_n730), .B2(new_n735), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n865), .B1(new_n869), .B2(new_n746), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n720), .A2(new_n644), .A3(new_n855), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(new_n704), .A3(new_n708), .A4(new_n857), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT111), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n845), .A2(new_n688), .A3(new_n847), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n874), .B1(new_n875), .B2(new_n834), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT111), .B1(new_n842), .B2(new_n848), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n873), .B(KEYINPUT53), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n867), .A2(new_n868), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n877), .A2(new_n876), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n833), .B1(new_n880), .B2(new_n866), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n873), .B(KEYINPUT53), .C1(new_n850), .C2(new_n849), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g697(.A(KEYINPUT113), .B(new_n879), .C1(new_n883), .C2(new_n868), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n881), .A2(new_n882), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT113), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT54), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n832), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(G952), .A2(G953), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n800), .B1(new_n888), .B2(new_n889), .ZN(G75));
  NAND2_X1  g704(.A1(new_n460), .A2(G953), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT118), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT119), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n867), .A2(new_n878), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(G902), .ZN(new_n897));
  INV_X1    g711(.A(G210), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n409), .A2(new_n421), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT117), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n419), .B(KEYINPUT55), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n901), .B(new_n902), .Z(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n895), .B(new_n903), .C1(new_n897), .C2(new_n898), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n894), .B1(new_n905), .B2(new_n906), .ZN(G51));
  INV_X1    g721(.A(new_n892), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n317), .B1(new_n867), .B2(new_n878), .ZN(new_n909));
  INV_X1    g723(.A(new_n756), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n909), .A2(KEYINPUT120), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT120), .B1(new_n909), .B2(new_n910), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n757), .B(KEYINPUT57), .Z(new_n914));
  AND3_X1   g728(.A1(new_n867), .A2(new_n868), .A3(new_n878), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n868), .B1(new_n867), .B2(new_n878), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n595), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n908), .B1(new_n913), .B2(new_n918), .ZN(G54));
  AND2_X1   g733(.A1(new_n507), .A2(new_n510), .ZN(new_n920));
  NAND2_X1  g734(.A1(KEYINPUT58), .A2(G475), .ZN(new_n921));
  OR3_X1    g735(.A1(new_n897), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n920), .B1(new_n897), .B2(new_n921), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n908), .B1(new_n922), .B2(new_n923), .ZN(G60));
  AND2_X1   g738(.A1(new_n619), .A2(new_n620), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n622), .B(KEYINPUT59), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(new_n915), .B2(new_n916), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n893), .ZN(new_n929));
  INV_X1    g743(.A(new_n926), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n884), .A2(new_n887), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n929), .B1(new_n925), .B2(new_n931), .ZN(G63));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n933));
  NAND2_X1  g747(.A1(G217), .A2(G902), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT60), .Z(new_n935));
  NAND3_X1  g749(.A1(new_n896), .A2(new_n640), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n893), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n362), .B(KEYINPUT121), .Z(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n896), .B2(new_n935), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n933), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n940), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n942), .A2(KEYINPUT61), .A3(new_n893), .A4(new_n936), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n943), .ZN(G66));
  AOI21_X1  g758(.A(new_n352), .B1(new_n463), .B2(G224), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT122), .Z(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n859), .B2(G953), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n901), .B1(G898), .B2(new_n352), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT123), .Z(new_n949));
  XNOR2_X1  g763(.A(new_n947), .B(new_n949), .ZN(G69));
  OR2_X1    g764(.A1(new_n738), .A2(new_n853), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n677), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n953), .A2(KEYINPUT124), .A3(new_n371), .ZN(new_n954));
  AOI21_X1  g768(.A(KEYINPUT124), .B1(new_n953), .B2(new_n371), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n782), .B(new_n791), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n845), .A2(new_n688), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n679), .A2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n679), .A2(KEYINPUT62), .A3(new_n957), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(G953), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n267), .B1(new_n259), .B2(new_n258), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n503), .B1(KEYINPUT19), .B2(new_n335), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(G900), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n966), .B1(new_n968), .B2(new_n352), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n748), .A2(new_n782), .A3(new_n791), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n736), .A2(new_n764), .A3(new_n836), .ZN(new_n971));
  INV_X1    g785(.A(new_n752), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n971), .A2(new_n972), .A3(new_n957), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n969), .B1(new_n974), .B2(new_n352), .ZN(new_n975));
  OAI21_X1  g789(.A(G953), .B1(new_n575), .B2(new_n968), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n966), .B2(KEYINPUT125), .ZN(new_n977));
  OR3_X1    g791(.A1(new_n967), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n977), .B1(new_n967), .B2(new_n975), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(G72));
  INV_X1    g794(.A(new_n298), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n192), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT126), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n981), .A2(new_n192), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(G472), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT63), .Z(new_n987));
  OAI21_X1  g801(.A(new_n892), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n962), .A2(new_n984), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n974), .A2(new_n983), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n988), .B1(new_n991), .B2(new_n859), .ZN(new_n992));
  INV_X1    g806(.A(new_n987), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n279), .A2(new_n281), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n993), .B1(new_n994), .B2(new_n299), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n992), .B(KEYINPUT127), .C1(new_n883), .C2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT127), .ZN(new_n998));
  INV_X1    g812(.A(new_n988), .ZN(new_n999));
  AOI22_X1  g813(.A1(new_n962), .A2(new_n984), .B1(new_n974), .B2(new_n983), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n999), .B1(new_n1000), .B2(new_n872), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n883), .A2(new_n996), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n997), .A2(new_n1003), .ZN(G57));
endmodule


