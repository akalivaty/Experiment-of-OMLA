//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n555, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1105, new_n1106;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT67), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G221), .A3(G219), .A4(G220), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  OR4_X1    g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT68), .Z(new_n456));
  AOI21_X1  g031(.A(new_n456), .B1(G567), .B2(new_n452), .ZN(G319));
  NAND2_X1  g032(.A1(G113), .A2(G2104), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n458), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT3), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n469), .A2(G137), .A3(new_n470), .A4(new_n460), .ZN(new_n471));
  NOR3_X1   g046(.A1(new_n467), .A2(new_n468), .A3(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n466), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n469), .A2(new_n470), .A3(new_n460), .ZN(new_n478));
  INV_X1    g053(.A(G136), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n469), .A2(G2105), .A3(new_n460), .ZN(new_n481));
  OAI221_X1 g056(.A(new_n477), .B1(new_n478), .B2(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT70), .ZN(G162));
  NAND4_X1  g058(.A1(new_n469), .A2(G138), .A3(new_n470), .A4(new_n460), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  AND4_X1   g063(.A1(new_n486), .A2(new_n488), .A3(new_n460), .A4(new_n462), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n469), .A2(G126), .A3(G2105), .A4(new_n460), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT71), .B(G114), .ZN(new_n494));
  OAI211_X1 g069(.A(G2104), .B(new_n493), .C1(new_n494), .C2(new_n470), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT72), .B1(new_n500), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n500), .A2(G543), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT74), .A3(G62), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT74), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n505), .A2(new_n506), .ZN(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n508), .A2(new_n509), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G50), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n505), .A2(G88), .A3(new_n506), .A4(new_n516), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n518), .A2(KEYINPUT73), .A3(new_n519), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n515), .A2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND3_X1  g101(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n517), .A2(G51), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n507), .A2(new_n516), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n527), .B(new_n528), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT75), .ZN(new_n533));
  XOR2_X1   g108(.A(new_n533), .B(KEYINPUT7), .Z(new_n534));
  OR2_X1    g109(.A1(new_n531), .A2(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  AOI22_X1  g111(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G651), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n517), .A2(G52), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n529), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G171));
  AOI22_X1  g118(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n538), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  INV_X1    g121(.A(new_n517), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT76), .B(G43), .Z(new_n548));
  OAI22_X1  g123(.A1(new_n529), .A2(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT77), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT78), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  NAND2_X1  g134(.A1(KEYINPUT79), .A2(KEYINPUT9), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n517), .A2(G53), .A3(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(KEYINPUT79), .A2(KEYINPUT9), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n561), .B(new_n562), .Z(new_n563));
  AOI22_X1  g138(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n538), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n507), .A2(new_n516), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G91), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n563), .A2(new_n565), .A3(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  OAI21_X1  g144(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n507), .A2(G87), .A3(new_n516), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n517), .A2(G49), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  AOI22_X1  g148(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(new_n538), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n517), .A2(G48), .ZN(new_n576));
  INV_X1    g151(.A(G86), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n529), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G305));
  XOR2_X1   g155(.A(KEYINPUT80), .B(G85), .Z(new_n581));
  AOI22_X1  g156(.A1(new_n566), .A2(new_n581), .B1(G47), .B2(new_n517), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n538), .B2(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n566), .A2(G92), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT81), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT10), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n586), .B(KEYINPUT81), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n511), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(G54), .B2(new_n517), .ZN(new_n596));
  AND3_X1   g171(.A1(new_n589), .A2(new_n592), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n585), .B1(new_n597), .B2(G868), .ZN(G284));
  OAI21_X1  g173(.A(new_n585), .B1(new_n597), .B2(G868), .ZN(G321));
  NAND2_X1  g174(.A1(G286), .A2(G868), .ZN(new_n600));
  INV_X1    g175(.A(G299), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G297));
  OAI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n597), .B1(new_n604), .B2(G860), .ZN(G148));
  NAND2_X1  g180(.A1(new_n597), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g184(.A1(G99), .A2(G2105), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n610), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n611));
  INV_X1    g186(.A(G135), .ZN(new_n612));
  INV_X1    g187(.A(G123), .ZN(new_n613));
  OAI221_X1 g188(.A(new_n611), .B1(new_n478), .B2(new_n612), .C1(new_n613), .C2(new_n481), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(G2096), .Z(new_n615));
  INV_X1    g190(.A(new_n463), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(new_n472), .ZN(new_n617));
  XOR2_X1   g192(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT83), .B(G2100), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(KEYINPUT84), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT13), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n619), .B(new_n622), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n615), .B(new_n623), .C1(KEYINPUT84), .C2(new_n620), .ZN(G156));
  XNOR2_X1  g199(.A(G2427), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2430), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT15), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2435), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(KEYINPUT14), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n629), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G1341), .B(G1348), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(G14), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n637), .A2(new_n638), .ZN(G401));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2067), .B(G2678), .Z(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(new_n644), .A3(KEYINPUT17), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT18), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2072), .B(G2078), .Z(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(new_n643), .B2(KEYINPUT18), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2096), .B(G2100), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT86), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G227));
  XOR2_X1   g229(.A(G1956), .B(G2474), .Z(new_n655));
  XOR2_X1   g230(.A(G1961), .B(G1966), .Z(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1971), .B(G1976), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n655), .A2(new_n656), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT20), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n658), .A2(new_n660), .A3(new_n662), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n665), .B(new_n666), .C1(new_n664), .C2(new_n663), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  INV_X1    g245(.A(G1981), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G1986), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n669), .B(new_n673), .ZN(G229));
  INV_X1    g249(.A(G16), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n675), .A2(G22), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(G303), .B2(G16), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1971), .ZN(new_n678));
  NOR2_X1   g253(.A1(G16), .A2(G23), .ZN(new_n679));
  INV_X1    g254(.A(G288), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(G16), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT33), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(G6), .A2(G16), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n579), .B2(G16), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT32), .B(G1981), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n678), .A2(new_n683), .A3(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT34), .Z(new_n689));
  MUX2_X1   g264(.A(G24), .B(G290), .S(G16), .Z(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(G1986), .Z(new_n691));
  INV_X1    g266(.A(new_n481), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G119), .ZN(new_n693));
  INV_X1    g268(.A(new_n478), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G131), .ZN(new_n695));
  OAI21_X1  g270(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n470), .A2(G107), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n693), .B(new_n695), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G25), .B(new_n698), .S(G29), .Z(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT35), .B(G1991), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n699), .B(new_n700), .Z(new_n701));
  NAND3_X1  g276(.A1(new_n689), .A2(new_n691), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT36), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n614), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n552), .A2(new_n675), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n675), .B2(G19), .ZN(new_n707));
  INV_X1    g282(.A(G1341), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT25), .Z(new_n711));
  INV_X1    g286(.A(G139), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n616), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n713));
  OAI221_X1 g288(.A(new_n711), .B1(new_n478), .B2(new_n712), .C1(new_n713), .C2(new_n470), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n704), .A2(G33), .ZN(new_n716));
  INV_X1    g291(.A(G2072), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n715), .B(new_n716), .C1(KEYINPUT87), .C2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(KEYINPUT87), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n718), .B(new_n719), .Z(new_n720));
  INV_X1    g295(.A(G2084), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT88), .B(KEYINPUT24), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G34), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(new_n704), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n474), .B2(new_n704), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT27), .B(G1996), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n692), .A2(G129), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n694), .A2(G141), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n472), .A2(G105), .ZN(new_n729));
  NAND3_X1  g304(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT26), .Z(new_n731));
  NAND4_X1  g306(.A1(new_n727), .A2(new_n728), .A3(new_n729), .A4(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n732), .A2(new_n704), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(KEYINPUT89), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G29), .B2(G32), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n734), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  OAI221_X1 g312(.A(new_n720), .B1(new_n721), .B2(new_n725), .C1(new_n726), .C2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT90), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n738), .A2(new_n739), .ZN(new_n741));
  OAI22_X1  g316(.A1(new_n740), .A2(new_n741), .B1(new_n708), .B2(new_n707), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT91), .ZN(new_n743));
  INV_X1    g318(.A(G35), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(G29), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n704), .A2(KEYINPUT91), .A3(G35), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n745), .B(new_n746), .C1(G162), .C2(new_n704), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT29), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(G2090), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n675), .A2(G20), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT92), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT23), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G299), .B2(G16), .ZN(new_n753));
  INV_X1    g328(.A(G1956), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n749), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n737), .A2(new_n726), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n675), .A2(G21), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G168), .B2(new_n675), .ZN(new_n759));
  INV_X1    g334(.A(G1966), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n748), .A2(G2090), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n756), .A2(new_n757), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n704), .A2(G26), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n692), .A2(G128), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n694), .A2(G140), .ZN(new_n766));
  OAI21_X1  g341(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n470), .A2(G116), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n765), .B(new_n766), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n764), .B1(new_n769), .B2(G29), .ZN(new_n770));
  MUX2_X1   g345(.A(new_n764), .B(new_n770), .S(KEYINPUT28), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G2067), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n704), .A2(G27), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G164), .B2(new_n704), .ZN(new_n774));
  INV_X1    g349(.A(G2078), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT31), .B(G11), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT30), .B(G28), .Z(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(G29), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n725), .B2(new_n721), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n772), .A2(new_n776), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n675), .A2(G5), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G171), .B2(new_n675), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1961), .ZN(new_n784));
  NOR4_X1   g359(.A1(new_n742), .A2(new_n763), .A3(new_n781), .A4(new_n784), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n703), .A2(new_n705), .A3(new_n709), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n675), .A2(G4), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n597), .B2(new_n675), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1348), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n786), .A2(new_n789), .ZN(G311));
  AND3_X1   g365(.A1(new_n703), .A2(new_n709), .A3(new_n785), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT93), .ZN(new_n792));
  INV_X1    g367(.A(new_n789), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n791), .A2(new_n792), .A3(new_n793), .A4(new_n705), .ZN(new_n794));
  OAI21_X1  g369(.A(KEYINPUT93), .B1(new_n786), .B2(new_n789), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(G150));
  NAND2_X1  g371(.A1(new_n517), .A2(G55), .ZN(new_n797));
  INV_X1    g372(.A(G93), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n529), .B2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT94), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n803));
  OAI22_X1  g378(.A1(new_n801), .A2(new_n802), .B1(new_n538), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(G860), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT37), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n597), .A2(G559), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n552), .A2(new_n804), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n550), .B2(new_n804), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n807), .B(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n806), .B1(new_n812), .B2(G860), .ZN(G145));
  NAND3_X1  g388(.A1(new_n694), .A2(KEYINPUT97), .A3(G142), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n692), .A2(G130), .ZN(new_n815));
  OR2_X1    g390(.A1(G106), .A2(G2105), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n816), .B(G2104), .C1(G118), .C2(new_n470), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT97), .ZN(new_n818));
  INV_X1    g393(.A(G142), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n478), .B2(new_n819), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n814), .A2(new_n815), .A3(new_n817), .A4(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(new_n619), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n698), .B(KEYINPUT98), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT99), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n732), .B(new_n498), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n769), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n714), .A2(KEYINPUT96), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n714), .B(KEYINPUT96), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(new_n827), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n825), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(G162), .B(KEYINPUT95), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G160), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(new_n614), .Z(new_n835));
  AND2_X1   g410(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  MUX2_X1   g411(.A(new_n824), .B(new_n825), .S(new_n831), .Z(new_n837));
  NOR2_X1   g412(.A1(new_n837), .A2(new_n835), .ZN(new_n838));
  NOR3_X1   g413(.A1(new_n836), .A2(new_n838), .A3(G37), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT40), .Z(G395));
  INV_X1    g415(.A(KEYINPUT102), .ZN(new_n841));
  XNOR2_X1  g416(.A(G303), .B(KEYINPUT100), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G305), .ZN(new_n843));
  XNOR2_X1  g418(.A(G290), .B(G288), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n841), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT102), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n843), .A2(new_n844), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT101), .B1(new_n843), .B2(new_n844), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n845), .B(new_n847), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n597), .A2(G299), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n589), .A2(new_n592), .A3(new_n596), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(new_n601), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT41), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n606), .B(new_n809), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n859), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(new_n856), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT42), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n863), .B1(new_n860), .B2(new_n862), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n852), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n860), .A2(new_n862), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT42), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n850), .A2(new_n851), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n847), .A2(new_n845), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .A4(new_n864), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n867), .A2(new_n872), .A3(G868), .ZN(new_n873));
  INV_X1    g448(.A(G868), .ZN(new_n874));
  AOI21_X1  g449(.A(KEYINPUT103), .B1(new_n804), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n867), .A2(new_n872), .A3(KEYINPUT103), .A4(G868), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(G295));
  AND2_X1   g453(.A1(new_n876), .A2(new_n877), .ZN(G331));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n880));
  AOI21_X1  g455(.A(G286), .B1(new_n880), .B2(G171), .ZN(new_n881));
  NAND2_X1  g456(.A1(G301), .A2(KEYINPUT104), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n809), .B(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n856), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n856), .B(KEYINPUT41), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n885), .B1(new_n886), .B2(new_n884), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n887), .A2(new_n870), .A3(new_n871), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n809), .A2(new_n883), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n809), .A2(new_n883), .ZN(new_n892));
  AOI22_X1  g467(.A1(new_n891), .A2(new_n892), .B1(new_n855), .B2(new_n853), .ZN(new_n893));
  INV_X1    g468(.A(new_n884), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n893), .B1(new_n858), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(G37), .B1(new_n895), .B2(new_n852), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n887), .A2(KEYINPUT105), .A3(new_n870), .A4(new_n871), .ZN(new_n897));
  AND4_X1   g472(.A1(KEYINPUT43), .A2(new_n890), .A3(new_n896), .A4(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT43), .B1(new_n896), .B2(new_n888), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT44), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n890), .A2(new_n901), .A3(new_n896), .A4(new_n897), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n896), .A2(new_n888), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT43), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n900), .A2(new_n907), .ZN(G397));
  INV_X1    g483(.A(G1384), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n489), .B1(new_n484), .B2(KEYINPUT4), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n909), .B1(new_n910), .B2(new_n496), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT45), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n466), .A2(G40), .A3(new_n471), .A4(new_n473), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G2067), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n769), .B(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n732), .B(G1996), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n915), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT106), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n698), .B(new_n700), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n921), .B1(new_n915), .B2(new_n922), .ZN(new_n923));
  AND2_X1   g498(.A1(G290), .A2(G1986), .ZN(new_n924));
  NOR2_X1   g499(.A1(G290), .A2(G1986), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n915), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT107), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n911), .A2(KEYINPUT50), .ZN(new_n929));
  INV_X1    g504(.A(new_n914), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT50), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n931), .B(new_n909), .C1(new_n910), .C2(new_n496), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(G1348), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(G1384), .B1(new_n491), .B2(new_n497), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(new_n916), .A3(new_n930), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT121), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n911), .A2(new_n914), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT121), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n941), .A3(new_n916), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT60), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n935), .A2(KEYINPUT60), .A3(new_n942), .A4(new_n938), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT123), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n597), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n854), .A2(new_n944), .A3(KEYINPUT123), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OR2_X1    g523(.A1(new_n944), .A2(KEYINPUT123), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n943), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT57), .ZN(new_n951));
  NAND2_X1  g526(.A1(G299), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n563), .A2(KEYINPUT57), .A3(new_n565), .A4(new_n567), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT117), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n956), .B(new_n930), .C1(new_n936), .C2(new_n931), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n932), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n914), .B1(new_n911), .B2(KEYINPUT50), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(new_n956), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n754), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT120), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT120), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n963), .B(new_n754), .C1(new_n958), .C2(new_n960), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n936), .A2(KEYINPUT45), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n966), .A2(new_n930), .A3(new_n913), .ZN(new_n967));
  XNOR2_X1  g542(.A(KEYINPUT56), .B(G2072), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n955), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n969), .ZN(new_n971));
  AOI211_X1 g546(.A(new_n954), .B(new_n971), .C1(new_n962), .C2(new_n964), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n950), .B1(new_n973), .B2(KEYINPUT61), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT61), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n975), .B1(new_n970), .B2(new_n972), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT122), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g553(.A(KEYINPUT122), .B(new_n975), .C1(new_n970), .C2(new_n972), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n966), .A2(new_n930), .A3(new_n913), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT58), .B(G1341), .ZN(new_n981));
  OAI22_X1  g556(.A1(new_n980), .A2(G1996), .B1(new_n940), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n552), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT59), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n974), .A2(new_n978), .A3(new_n979), .A4(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n972), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n854), .B1(new_n942), .B2(new_n939), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n986), .B1(new_n987), .B2(new_n970), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n985), .A2(KEYINPUT124), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT124), .B1(new_n985), .B2(new_n988), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n967), .A2(new_n775), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT126), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n991), .B(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n992), .A2(KEYINPUT126), .ZN(new_n995));
  INV_X1    g570(.A(G1961), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n995), .B1(new_n933), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(G171), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n994), .A2(G301), .A3(new_n997), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1001), .B(KEYINPUT54), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n579), .A2(new_n671), .ZN(new_n1003));
  OAI21_X1  g578(.A(G1981), .B1(new_n575), .B2(new_n578), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(KEYINPUT49), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT115), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1003), .A2(new_n1004), .A3(new_n1007), .A4(KEYINPUT49), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G8), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n940), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT114), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1012), .A2(KEYINPUT114), .A3(new_n1013), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1009), .B(new_n1011), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n1017));
  INV_X1    g592(.A(G1976), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1011), .B(new_n1017), .C1(new_n1018), .C2(G288), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n680), .A2(G1976), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(new_n1011), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1019), .B(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1016), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G303), .A2(G8), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1010), .B1(new_n515), .B2(new_n524), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(KEYINPUT110), .A3(KEYINPUT55), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1026), .A2(KEYINPUT111), .A3(new_n1027), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1033), .B1(new_n1029), .B2(KEYINPUT55), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1024), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1037), .A2(KEYINPUT112), .A3(new_n1034), .A4(new_n1032), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  OR2_X1    g614(.A1(new_n933), .A2(G2090), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT109), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT108), .B(G1971), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n980), .A2(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1041), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1044), .A2(new_n1045), .A3(new_n1010), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1023), .B1(new_n1039), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n958), .A2(KEYINPUT118), .A3(new_n960), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(G2090), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT118), .B1(new_n958), .B2(new_n960), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1050), .A2(new_n1051), .B1(new_n1042), .B2(new_n980), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1048), .B1(new_n1052), .B2(new_n1010), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1047), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n980), .A2(new_n760), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n959), .A2(new_n721), .A3(new_n932), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(G8), .ZN(new_n1059));
  NAND2_X1  g634(.A1(G286), .A2(G8), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT125), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT51), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  OR2_X1    g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1064), .B(new_n1065), .C1(G168), .C2(new_n1059), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1002), .A2(new_n1055), .A3(new_n1066), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n989), .A2(new_n990), .A3(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1059), .A2(G286), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1047), .A2(new_n1053), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT63), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT119), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1070), .A2(new_n1074), .A3(new_n1071), .ZN(new_n1075));
  OR3_X1    g650(.A1(new_n1046), .A2(new_n1031), .A3(new_n1035), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1047), .A2(new_n1076), .A3(KEYINPUT63), .A4(new_n1069), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1073), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1039), .A2(new_n1046), .A3(new_n1016), .A4(new_n1022), .ZN(new_n1079));
  XOR2_X1   g654(.A(new_n1011), .B(KEYINPUT116), .Z(new_n1080));
  NAND3_X1  g655(.A1(new_n1016), .A2(new_n1018), .A3(new_n680), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(new_n1003), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1054), .B1(KEYINPUT62), .B2(new_n1066), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1066), .A2(KEYINPUT62), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(new_n999), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1082), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1078), .A2(new_n1079), .A3(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n928), .B1(new_n1068), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n915), .B1(new_n918), .B2(new_n732), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n913), .A2(G1996), .A3(new_n914), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1090), .A2(KEYINPUT46), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(KEYINPUT46), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1089), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1093), .B(KEYINPUT127), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1094), .B(KEYINPUT47), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n921), .A2(new_n700), .A3(new_n698), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n769), .A2(G2067), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n915), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n925), .A2(new_n915), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1099), .B(KEYINPUT48), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n923), .A2(new_n1100), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1095), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1088), .A2(new_n1102), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g678(.A1(new_n839), .A2(G401), .A3(G227), .ZN(new_n1105));
  INV_X1    g679(.A(G229), .ZN(new_n1106));
  NAND4_X1  g680(.A1(new_n905), .A2(new_n1105), .A3(G319), .A4(new_n1106), .ZN(G225));
  INV_X1    g681(.A(G225), .ZN(G308));
endmodule


