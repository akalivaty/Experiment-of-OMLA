//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n552,
    new_n554, new_n555, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1179, new_n1180, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n463), .A3(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n461), .A2(new_n463), .A3(G137), .ZN(new_n467));
  NAND2_X1  g042(.A1(G101), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n470), .B(KEYINPUT66), .ZN(G160));
  OR2_X1    g046(.A1(G100), .A2(G2105), .ZN(new_n472));
  OAI211_X1 g047(.A(new_n472), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n461), .A2(new_n463), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n461), .A2(new_n463), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(KEYINPUT67), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n476), .A2(G2105), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  INV_X1    g055(.A(G136), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n476), .A2(new_n459), .A3(new_n478), .ZN(new_n482));
  OAI221_X1 g057(.A(new_n473), .B1(new_n479), .B2(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  OR2_X1    g059(.A1(new_n459), .A2(G114), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(G126), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n477), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n492), .A2(new_n461), .A3(new_n463), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n490), .B1(new_n495), .B2(new_n496), .ZN(G164));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(KEYINPUT6), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT68), .B1(new_n500), .B2(G651), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(new_n498), .A3(KEYINPUT6), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G88), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  AOI211_X1 g084(.A(new_n509), .B(new_n499), .C1(new_n501), .C2(new_n503), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G50), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n512), .A2(new_n498), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n508), .A2(new_n511), .A3(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  NAND3_X1  g090(.A1(new_n504), .A2(G51), .A3(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(G63), .A2(G651), .ZN(new_n521));
  OR3_X1    g096(.A1(new_n520), .A2(KEYINPUT69), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(KEYINPUT69), .B1(new_n520), .B2(new_n521), .ZN(new_n523));
  AND3_X1   g098(.A1(new_n516), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT70), .B(G89), .Z(new_n525));
  NAND3_X1  g100(.A1(new_n504), .A2(new_n505), .A3(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n527), .B1(new_n526), .B2(new_n529), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n524), .B1(new_n531), .B2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n520), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n504), .A2(G52), .A3(G543), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n538), .B(new_n539), .C1(new_n540), .C2(new_n506), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  NAND2_X1  g117(.A1(new_n510), .A2(G43), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n504), .A2(G81), .A3(new_n505), .ZN(new_n544));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n520), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G651), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n543), .A2(new_n544), .A3(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n552), .A2(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(new_n501), .A2(new_n503), .ZN(new_n557));
  INV_X1    g132(.A(new_n499), .ZN(new_n558));
  AND4_X1   g133(.A1(G91), .A2(new_n557), .A3(new_n558), .A4(new_n505), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n517), .A2(new_n519), .A3(G65), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n498), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n560), .A2(KEYINPUT74), .A3(new_n561), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n559), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n557), .A2(G53), .A3(G543), .A4(new_n558), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  XNOR2_X1  g143(.A(KEYINPUT72), .B(KEYINPUT9), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n504), .A2(G53), .A3(G543), .A4(new_n569), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n568), .B1(KEYINPUT73), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n570), .A2(KEYINPUT73), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n566), .B1(new_n571), .B2(new_n572), .ZN(G299));
  NAND2_X1  g148(.A1(new_n507), .A2(G87), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n510), .A2(G49), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(new_n507), .A2(G86), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n510), .A2(G48), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n505), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(new_n498), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(new_n507), .A2(G85), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(new_n498), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n510), .A2(G47), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n557), .A2(G92), .A3(new_n558), .A4(new_n505), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n504), .A2(KEYINPUT10), .A3(G92), .A4(new_n505), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT75), .ZN(new_n594));
  INV_X1    g169(.A(G79), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(new_n509), .ZN(new_n596));
  NAND3_X1  g171(.A1(KEYINPUT75), .A2(G79), .A3(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI211_X1 g173(.A(new_n596), .B(new_n597), .C1(new_n520), .C2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n510), .A2(G54), .B1(new_n599), .B2(G651), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n593), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n588), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n588), .B1(new_n601), .B2(G868), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT73), .ZN(new_n605));
  NAND4_X1  g180(.A1(new_n510), .A2(new_n605), .A3(G53), .A4(new_n569), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n570), .A2(KEYINPUT73), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n606), .A2(new_n607), .A3(new_n568), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n608), .A2(new_n566), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n604), .B1(new_n609), .B2(G868), .ZN(G297));
  OAI21_X1  g185(.A(new_n604), .B1(new_n609), .B2(G868), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n601), .B1(new_n612), .B2(G860), .ZN(G148));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n549), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n593), .A2(new_n600), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n616), .A2(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n615), .B1(new_n617), .B2(new_n614), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g194(.A1(new_n460), .A2(G2105), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n474), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT13), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n622), .A2(new_n623), .B1(KEYINPUT76), .B2(G2100), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n623), .B2(new_n622), .ZN(new_n625));
  NOR2_X1   g200(.A1(KEYINPUT76), .A2(G2100), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(G99), .A2(G2105), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n628), .B(G2104), .C1(G111), .C2(new_n459), .ZN(new_n629));
  INV_X1    g204(.A(G123), .ZN(new_n630));
  INV_X1    g205(.A(G135), .ZN(new_n631));
  OAI221_X1 g206(.A(new_n629), .B1(new_n479), .B2(new_n630), .C1(new_n631), .C2(new_n482), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2096), .Z(new_n633));
  NAND2_X1  g208(.A1(new_n627), .A2(new_n633), .ZN(G156));
  INV_X1    g209(.A(G14), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2435), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(KEYINPUT14), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G1341), .B(G1348), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT78), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n635), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n647), .A2(new_n649), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n651), .A2(KEYINPUT79), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT79), .ZN(new_n653));
  NOR3_X1   g228(.A1(new_n647), .A2(new_n653), .A3(new_n649), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n650), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT80), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g232(.A(KEYINPUT80), .B(new_n650), .C1(new_n652), .C2(new_n654), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G401));
  XNOR2_X1  g235(.A(G2072), .B(G2078), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT81), .Z(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT17), .Z(new_n663));
  XOR2_X1   g238(.A(G2067), .B(G2678), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n663), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n662), .A2(new_n666), .A3(new_n665), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT18), .Z(new_n672));
  AOI21_X1  g247(.A(new_n668), .B1(new_n662), .B2(KEYINPUT82), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n673), .B1(KEYINPUT82), .B2(new_n662), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n670), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2096), .B(G2100), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n681), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n679), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n679), .A2(new_n684), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n683), .B(new_n685), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n687), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1991), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G1996), .ZN(new_n691));
  INV_X1    g266(.A(G1991), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n689), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G1996), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  INV_X1    g274(.A(new_n697), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n691), .A2(new_n695), .A3(new_n700), .ZN(new_n701));
  AND3_X1   g276(.A1(new_n698), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n699), .B1(new_n698), .B2(new_n701), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(G229));
  INV_X1    g279(.A(KEYINPUT94), .ZN(new_n705));
  INV_X1    g280(.A(new_n482), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n706), .A2(G141), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT93), .ZN(new_n708));
  INV_X1    g283(.A(new_n479), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G129), .ZN(new_n710));
  NAND3_X1  g285(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT26), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n713), .A2(new_n714), .B1(G105), .B2(new_n620), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n710), .A2(new_n715), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n708), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n705), .B1(new_n717), .B2(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n708), .A2(new_n716), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  NOR3_X1   g295(.A1(new_n719), .A2(KEYINPUT94), .A3(new_n720), .ZN(new_n721));
  OAI22_X1  g296(.A1(new_n718), .A2(new_n721), .B1(G29), .B2(G32), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT27), .B(G1996), .Z(new_n723));
  XOR2_X1   g298(.A(new_n722), .B(new_n723), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n720), .A2(G35), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G162), .B2(new_n720), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT29), .Z(new_n727));
  INV_X1    g302(.A(G2090), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G34), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n730), .A2(KEYINPUT24), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(KEYINPUT24), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n720), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G160), .B2(new_n720), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT92), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n729), .B1(G2084), .B2(new_n736), .ZN(new_n737));
  AND3_X1   g312(.A1(G168), .A2(KEYINPUT95), .A3(G16), .ZN(new_n738));
  AOI21_X1  g313(.A(KEYINPUT95), .B1(G168), .B2(G16), .ZN(new_n739));
  OAI22_X1  g314(.A1(new_n738), .A2(new_n739), .B1(G16), .B2(G21), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT96), .B(G1966), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G2084), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n727), .A2(new_n728), .B1(new_n744), .B2(new_n735), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n737), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n740), .A2(new_n742), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT98), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n720), .A2(G26), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT28), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n709), .A2(G128), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n706), .A2(G140), .ZN(new_n752));
  NOR3_X1   g327(.A1(KEYINPUT89), .A2(G104), .A3(G2105), .ZN(new_n753));
  OAI21_X1  g328(.A(KEYINPUT89), .B1(G104), .B2(G2105), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n754), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n751), .B(new_n752), .C1(new_n753), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G29), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n757), .A2(KEYINPUT90), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n757), .A2(KEYINPUT90), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n750), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G2067), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n720), .A2(G33), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(new_n459), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n620), .A2(G103), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT25), .Z(new_n767));
  INV_X1    g342(.A(G139), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n482), .B2(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(KEYINPUT91), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(KEYINPUT91), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n765), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n763), .B1(new_n772), .B2(new_n720), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(G2072), .Z(new_n774));
  NOR2_X1   g349(.A1(new_n632), .A2(new_n720), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT31), .B(G11), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT97), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n720), .B1(new_n778), .B2(G28), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n778), .B2(G28), .ZN(new_n780));
  NOR3_X1   g355(.A1(new_n775), .A2(new_n777), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(G171), .A2(G16), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G5), .B2(G16), .ZN(new_n783));
  INV_X1    g358(.A(G1961), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(G27), .A2(G29), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G164), .B2(G29), .ZN(new_n787));
  INV_X1    g362(.A(G2078), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n781), .A2(new_n785), .A3(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G16), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(G4), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n601), .B2(new_n791), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1348), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n783), .A2(new_n784), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n790), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n791), .A2(G19), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n550), .B2(new_n791), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT88), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1341), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n762), .A2(new_n774), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  NOR4_X1   g376(.A1(new_n724), .A2(new_n746), .A3(new_n748), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n791), .A2(G20), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n609), .B2(new_n791), .ZN(new_n804));
  MUX2_X1   g379(.A(new_n803), .B(new_n804), .S(KEYINPUT23), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT100), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT99), .B(G1956), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n720), .A2(G25), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n709), .A2(G119), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n706), .A2(G131), .ZN(new_n811));
  OR2_X1    g386(.A1(G95), .A2(G2105), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n812), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT83), .Z(new_n814));
  NAND3_X1  g389(.A1(new_n810), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(KEYINPUT84), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(KEYINPUT84), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n809), .B1(new_n819), .B2(new_n720), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT35), .B(G1991), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n791), .A2(G24), .ZN(new_n824));
  INV_X1    g399(.A(G290), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n825), .B2(new_n791), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(G1986), .Z(new_n827));
  NAND4_X1  g402(.A1(new_n822), .A2(KEYINPUT87), .A3(new_n823), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n791), .A2(G22), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(G166), .B2(new_n791), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(G1971), .Z(new_n831));
  MUX2_X1   g406(.A(G6), .B(G305), .S(G16), .Z(new_n832));
  XOR2_X1   g407(.A(KEYINPUT32), .B(G1981), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(G16), .A2(G23), .ZN(new_n835));
  INV_X1    g410(.A(G288), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n835), .B1(new_n836), .B2(G16), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT33), .B(G1976), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n831), .A2(new_n834), .A3(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT85), .B(KEYINPUT34), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n828), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n840), .A2(new_n841), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT86), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT36), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n843), .A2(new_n845), .A3(KEYINPUT36), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n802), .A2(new_n808), .A3(new_n848), .A4(new_n849), .ZN(G150));
  INV_X1    g425(.A(G150), .ZN(G311));
  INV_X1    g426(.A(KEYINPUT101), .ZN(new_n852));
  NAND2_X1  g427(.A1(G80), .A2(G543), .ZN(new_n853));
  INV_X1    g428(.A(G67), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n520), .B2(new_n854), .ZN(new_n855));
  AOI22_X1  g430(.A1(new_n510), .A2(G55), .B1(new_n855), .B2(G651), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n504), .A2(G93), .A3(new_n505), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n852), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(G651), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n504), .A2(G55), .A3(G543), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n857), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n861), .A2(KEYINPUT101), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(G860), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT37), .Z(new_n865));
  NAND2_X1  g440(.A1(new_n861), .A2(KEYINPUT101), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n856), .A2(new_n852), .A3(new_n857), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n550), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n549), .B1(new_n857), .B2(new_n856), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT39), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n616), .A2(new_n612), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT38), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n874), .A2(G860), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n871), .A2(new_n873), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n865), .B1(new_n875), .B2(new_n876), .ZN(G145));
  INV_X1    g452(.A(new_n489), .ZN(new_n878));
  AOI22_X1  g453(.A1(new_n474), .A2(new_n878), .B1(new_n485), .B2(new_n487), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n879), .B1(new_n880), .B2(new_n494), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n818), .B(new_n881), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n772), .B(new_n622), .Z(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n483), .B(new_n632), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n756), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(G160), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n887), .A2(G160), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n709), .A2(KEYINPUT102), .A3(G130), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n706), .A2(G142), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT102), .ZN(new_n893));
  INV_X1    g468(.A(G130), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n893), .B1(new_n479), .B2(new_n894), .ZN(new_n895));
  OR2_X1    g470(.A1(G106), .A2(G2105), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n896), .B(G2104), .C1(G118), .C2(new_n459), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n891), .A2(new_n892), .A3(new_n895), .A4(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n719), .B(new_n898), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n889), .A2(new_n890), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n887), .A2(G160), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n901), .B1(new_n902), .B2(new_n888), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n885), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(G37), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n899), .B1(new_n889), .B2(new_n890), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n902), .A2(new_n888), .A3(new_n901), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n884), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n904), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g485(.A(KEYINPUT103), .B1(G299), .B2(new_n601), .ZN(new_n911));
  NAND2_X1  g486(.A1(G299), .A2(new_n601), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n616), .A2(new_n608), .A3(new_n913), .A4(new_n566), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT105), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n913), .B1(new_n609), .B2(new_n616), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n912), .A2(new_n914), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n911), .A2(KEYINPUT41), .A3(new_n912), .A4(new_n914), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n917), .B1(new_n922), .B2(KEYINPUT105), .ZN(new_n923));
  INV_X1    g498(.A(new_n869), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n549), .B1(new_n858), .B2(new_n862), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(new_n617), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n915), .B(KEYINPUT104), .Z(new_n929));
  AOI21_X1  g504(.A(new_n928), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(G303), .B(G288), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n933));
  XNOR2_X1  g508(.A(G305), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n825), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n934), .A2(new_n825), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n932), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n934), .A2(new_n825), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(new_n931), .A3(new_n935), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(KEYINPUT42), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT107), .B1(new_n930), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n930), .A2(new_n942), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n930), .A2(KEYINPUT107), .A3(new_n942), .ZN(new_n946));
  OAI21_X1  g521(.A(G868), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n863), .A2(new_n614), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(G295));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n948), .ZN(G331));
  OAI211_X1 g525(.A(new_n524), .B(G301), .C1(new_n531), .C2(new_n532), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n526), .A2(new_n529), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT71), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n530), .ZN(new_n955));
  AOI21_X1  g530(.A(G301), .B1(new_n955), .B2(new_n524), .ZN(new_n956));
  OAI22_X1  g531(.A1(new_n952), .A2(new_n956), .B1(new_n868), .B2(new_n869), .ZN(new_n957));
  NAND2_X1  g532(.A1(G286), .A2(G171), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n924), .A2(new_n925), .A3(new_n958), .A4(new_n951), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n957), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n926), .B(KEYINPUT109), .C1(new_n952), .C2(new_n956), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n915), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n957), .A2(new_n959), .A3(new_n965), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n870), .A2(KEYINPUT108), .A3(new_n951), .A4(new_n958), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n941), .B(new_n964), .C1(new_n923), .C2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT110), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT105), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n971), .B1(new_n920), .B2(new_n921), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n967), .B(new_n966), .C1(new_n972), .C2(new_n917), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n973), .A2(new_n974), .A3(new_n941), .A4(new_n964), .ZN(new_n975));
  INV_X1    g550(.A(new_n941), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n912), .A2(new_n914), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT41), .B1(new_n977), .B2(new_n911), .ZN(new_n978));
  INV_X1    g553(.A(new_n921), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT105), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n917), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n968), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n963), .A2(new_n915), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n976), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n970), .A2(new_n905), .A3(new_n975), .A4(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(G37), .B1(new_n969), .B2(KEYINPUT110), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n929), .A2(new_n968), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n963), .B1(new_n920), .B2(new_n921), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n976), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AND4_X1   g566(.A1(KEYINPUT43), .A2(new_n988), .A3(new_n975), .A4(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT44), .B1(new_n987), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n988), .A2(new_n986), .A3(new_n975), .A4(new_n991), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n993), .A2(new_n998), .ZN(G397));
  XOR2_X1   g574(.A(KEYINPUT111), .B(G1384), .Z(new_n1000));
  NAND2_X1  g575(.A1(new_n881), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(KEYINPUT112), .B(G40), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n470), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n694), .ZN(new_n1007));
  XOR2_X1   g582(.A(new_n1007), .B(KEYINPUT46), .Z(new_n1008));
  INV_X1    g583(.A(new_n1006), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n756), .B(new_n761), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1009), .B1(new_n717), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g587(.A(new_n1012), .B(KEYINPUT47), .Z(new_n1013));
  NOR3_X1   g588(.A1(new_n1009), .A2(G1986), .A3(G290), .ZN(new_n1014));
  XOR2_X1   g589(.A(new_n1014), .B(KEYINPUT48), .Z(new_n1015));
  NOR2_X1   g590(.A1(new_n717), .A2(G1996), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n719), .A2(new_n694), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1010), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n818), .B(new_n821), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1015), .B1(new_n1020), .B2(new_n1009), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n818), .A2(new_n821), .ZN(new_n1022));
  OAI22_X1  g597(.A1(new_n1018), .A2(new_n1022), .B1(G2067), .B2(new_n756), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n1006), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1013), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(G305), .A2(G1981), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1026), .B(KEYINPUT117), .ZN(new_n1027));
  AND2_X1   g602(.A1(G305), .A2(G1981), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1028), .A2(new_n1026), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT49), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(KEYINPUT116), .A3(KEYINPUT49), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1029), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1005), .ZN(new_n1037));
  INV_X1    g612(.A(G1384), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n881), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G8), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1034), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G1976), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n836), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1027), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n881), .A2(new_n1038), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1046), .A2(new_n1005), .ZN(new_n1047));
  INV_X1    g622(.A(G8), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1005), .B1(new_n1046), .B2(new_n1002), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n881), .A2(KEYINPUT45), .A3(new_n1000), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT113), .B(G1971), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n881), .A2(new_n1056), .A3(new_n1038), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1055), .A2(new_n1057), .A3(new_n1037), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(G2090), .ZN(new_n1059));
  OAI21_X1  g634(.A(G8), .B1(new_n1054), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n1061));
  NAND2_X1  g636(.A1(G303), .A2(G8), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  NAND4_X1  g640(.A1(G303), .A2(KEYINPUT114), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1060), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT52), .B1(G288), .B2(new_n1043), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1049), .B(new_n1070), .C1(new_n1043), .C2(G288), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1040), .B1(G1976), .B2(new_n836), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1071), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1074), .B1(new_n1034), .B2(new_n1041), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1045), .A2(new_n1049), .B1(new_n1069), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1060), .A2(new_n1067), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1075), .A2(new_n1068), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(new_n1046), .B2(new_n1002), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n881), .A2(KEYINPUT118), .A3(KEYINPUT45), .A4(new_n1038), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(new_n1050), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n742), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1058), .A2(G2084), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1085), .A2(G8), .A3(G168), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT63), .B1(new_n1078), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1075), .A2(new_n1068), .A3(new_n1077), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT63), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1089), .A2(new_n1090), .A3(new_n1086), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1076), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1052), .A2(new_n788), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1093), .A2(new_n1094), .B1(new_n784), .B2(new_n1058), .ZN(new_n1095));
  OR3_X1    g670(.A1(new_n1082), .A2(new_n1094), .A3(G2078), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(G171), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1098), .A2(KEYINPUT62), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1085), .A2(G8), .ZN(new_n1100));
  NAND2_X1  g675(.A1(G286), .A2(G8), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT51), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(G168), .A2(new_n1048), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n1103), .B2(new_n1085), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1100), .A2(KEYINPUT51), .A3(new_n1101), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1099), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n1107));
  NAND3_X1  g682(.A1(G299), .A2(new_n1107), .A3(KEYINPUT57), .ZN(new_n1108));
  NAND2_X1  g683(.A1(G299), .A2(new_n1107), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(G1956), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1058), .A2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT56), .B(G2072), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1050), .A2(new_n1051), .A3(new_n1114), .ZN(new_n1115));
  AND4_X1   g690(.A1(new_n1108), .A2(new_n1111), .A3(new_n1113), .A4(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1111), .A2(new_n1108), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1111), .A2(KEYINPUT121), .A3(new_n1108), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1113), .A2(KEYINPUT120), .A3(new_n1115), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT120), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1119), .B(new_n1120), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(G1348), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1058), .A2(new_n1124), .B1(new_n1047), .B2(new_n761), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1125), .A2(new_n616), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1116), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1116), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1123), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1058), .A2(new_n1124), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1047), .A2(new_n761), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1131), .A2(KEYINPUT60), .A3(new_n616), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(KEYINPUT124), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1131), .A2(KEYINPUT60), .A3(new_n1132), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n601), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1125), .A2(new_n1137), .A3(KEYINPUT60), .A4(new_n616), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1134), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n1125), .A2(KEYINPUT60), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  XOR2_X1   g716(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1142));
  NAND2_X1  g717(.A1(new_n1052), .A2(new_n694), .ZN(new_n1143));
  XOR2_X1   g718(.A(KEYINPUT58), .B(G1341), .Z(new_n1144));
  NAND2_X1  g719(.A1(new_n1039), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1142), .B1(new_n1146), .B2(new_n550), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1142), .ZN(new_n1148));
  AOI211_X1 g723(.A(new_n549), .B(new_n1148), .C1(new_n1143), .C2(new_n1145), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1130), .A2(new_n1141), .A3(new_n1150), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1111), .A2(new_n1108), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1128), .B1(new_n1116), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT123), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1127), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(KEYINPUT125), .B(G2078), .ZN(new_n1157));
  AND4_X1   g732(.A1(KEYINPUT53), .A2(new_n470), .A3(G40), .A4(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1003), .A2(new_n1158), .A3(new_n1051), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1095), .A2(G301), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT126), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT54), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1095), .A2(new_n1163), .A3(G301), .A4(new_n1159), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1161), .A2(new_n1098), .A3(new_n1162), .A4(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1097), .A2(G301), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1095), .A2(G171), .A3(new_n1159), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1166), .A2(KEYINPUT54), .A3(new_n1167), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1106), .B1(new_n1156), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1104), .B(new_n1105), .C1(new_n1171), .C2(new_n1098), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1172), .A2(new_n1078), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1092), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  XOR2_X1   g749(.A(G290), .B(G1986), .Z(new_n1175));
  AOI21_X1  g750(.A(new_n1009), .B1(new_n1020), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1025), .B1(new_n1174), .B2(new_n1176), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g752(.A(G319), .ZN(new_n1179));
  OR2_X1    g753(.A1(G227), .A2(new_n1179), .ZN(new_n1180));
  NOR3_X1   g754(.A1(new_n702), .A2(new_n703), .A3(new_n1180), .ZN(new_n1181));
  NAND3_X1  g755(.A1(new_n909), .A2(new_n659), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g756(.A(new_n1182), .B1(new_n994), .B2(new_n995), .ZN(G308));
  NAND4_X1  g757(.A1(new_n996), .A2(new_n659), .A3(new_n909), .A4(new_n1181), .ZN(G225));
endmodule


