//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1283, new_n1284, new_n1285, new_n1286;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n207), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OR2_X1    g0009(.A1(new_n207), .A2(KEYINPUT66), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n207), .A2(KEYINPUT66), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n210), .A2(G50), .A3(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G1), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n215), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT0), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n218), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT67), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  INV_X1    g0027(.A(G238), .ZN(new_n228));
  INV_X1    g0028(.A(G87), .ZN(new_n229));
  INV_X1    g0029(.A(G250), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n227), .B1(new_n202), .B2(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n232));
  AOI22_X1  g0032(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n221), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT1), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n226), .A2(new_n236), .ZN(G361));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G226), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(KEYINPUT72), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  INV_X1    g0055(.A(G45), .ZN(new_n256));
  AOI21_X1  g0056(.A(G1), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G1), .A3(G13), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(new_n259), .A3(G274), .ZN(new_n260));
  INV_X1    g0060(.A(G226), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n219), .B1(G41), .B2(G45), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT3), .B(G33), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G223), .A3(G1698), .ZN(new_n266));
  INV_X1    g0066(.A(G77), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G222), .ZN(new_n270));
  OAI221_X1 g0070(.A(new_n266), .B1(new_n267), .B2(new_n265), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n259), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n264), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G200), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n254), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT10), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(G190), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT73), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n273), .A2(new_n274), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT72), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n214), .ZN(new_n284));
  INV_X1    g0084(.A(G50), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n215), .B1(new_n206), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n215), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(G150), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI22_X1  g0091(.A1(new_n287), .A2(new_n288), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n284), .B1(new_n286), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G13), .ZN(new_n294));
  NOR3_X1   g0094(.A1(new_n294), .A2(new_n215), .A3(G1), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(new_n284), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n285), .B1(new_n219), .B2(G20), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n296), .A2(new_n297), .B1(new_n285), .B2(new_n295), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT9), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n279), .A2(new_n280), .A3(new_n282), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n282), .A2(new_n300), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT73), .B1(new_n302), .B2(new_n278), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n300), .B(new_n277), .C1(new_n274), .C2(new_n273), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n273), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT69), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n299), .B1(new_n273), .B2(G169), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n287), .B1(new_n219), .B2(G20), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n315), .A2(new_n296), .B1(new_n295), .B2(new_n287), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n284), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G58), .A2(G68), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n203), .A2(new_n205), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G20), .ZN(new_n321));
  INV_X1    g0121(.A(G159), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n322), .A2(G20), .A3(G33), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT77), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT77), .ZN(new_n326));
  AOI211_X1 g0126(.A(new_n326), .B(new_n323), .C1(new_n320), .C2(G20), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT7), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(new_n265), .B2(G20), .ZN(new_n330));
  INV_X1    g0130(.A(G33), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT3), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT3), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G33), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(KEYINPUT7), .A3(new_n215), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n202), .B1(new_n330), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT16), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n318), .B1(new_n328), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n321), .A2(new_n324), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n326), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n321), .A2(KEYINPUT77), .A3(new_n324), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT7), .B1(new_n335), .B2(new_n215), .ZN(new_n344));
  AOI211_X1 g0144(.A(new_n329), .B(G20), .C1(new_n332), .C2(new_n334), .ZN(new_n345));
  OAI21_X1  g0145(.A(G68), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n342), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n338), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n317), .B1(new_n340), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G232), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n260), .B1(new_n350), .B2(new_n263), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n265), .A2(G226), .A3(G1698), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n265), .A2(G223), .A3(new_n268), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G87), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n351), .B1(new_n355), .B2(new_n272), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n308), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(G169), .B2(new_n356), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT18), .B1(new_n349), .B2(new_n358), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n342), .A2(KEYINPUT16), .A3(new_n343), .A4(new_n346), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n284), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT16), .B1(new_n328), .B2(new_n346), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n316), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT18), .ZN(new_n364));
  INV_X1    g0164(.A(new_n358), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n359), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT78), .B(KEYINPUT17), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n355), .A2(new_n272), .ZN(new_n369));
  INV_X1    g0169(.A(G190), .ZN(new_n370));
  INV_X1    g0170(.A(new_n351), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(G200), .B2(new_n356), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n368), .B1(new_n349), .B2(new_n373), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n325), .A2(new_n327), .A3(new_n337), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n284), .B(new_n360), .C1(new_n375), .C2(KEYINPUT16), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT17), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n377), .A2(KEYINPUT78), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  AND4_X1   g0179(.A1(new_n376), .A2(new_n316), .A3(new_n373), .A4(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n374), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n260), .ZN(new_n382));
  INV_X1    g0182(.A(new_n263), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n382), .B1(G244), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n265), .A2(G238), .A3(G1698), .ZN(new_n385));
  INV_X1    g0185(.A(G107), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n385), .B1(new_n386), .B2(new_n265), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT70), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n265), .A2(new_n388), .A3(G232), .A4(new_n268), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT70), .B1(new_n269), .B2(new_n350), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n387), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n384), .B1(new_n391), .B2(new_n259), .ZN(new_n392));
  INV_X1    g0192(.A(G169), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n229), .A2(KEYINPUT15), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT15), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G87), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n398), .A2(new_n288), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n287), .A2(new_n291), .B1(new_n215), .B2(new_n267), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n284), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n219), .A2(G20), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n296), .A2(G77), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n294), .A2(G1), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G20), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n401), .B(new_n403), .C1(G77), .C2(new_n405), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n308), .B(new_n384), .C1(new_n391), .C2(new_n259), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n394), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n406), .B1(new_n392), .B2(G200), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT71), .ZN(new_n410));
  OAI22_X1  g0210(.A1(new_n409), .A2(new_n410), .B1(new_n370), .B2(new_n392), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n409), .A2(new_n410), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NOR4_X1   g0213(.A1(new_n314), .A2(new_n367), .A3(new_n381), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n295), .A2(new_n202), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n415), .B(KEYINPUT12), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n290), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n267), .B2(new_n288), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n418), .A2(KEYINPUT11), .A3(new_n284), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n296), .A2(G68), .A3(new_n402), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n416), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT11), .B1(new_n418), .B2(new_n284), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(KEYINPUT76), .A2(KEYINPUT14), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n332), .A2(new_n334), .A3(G226), .A4(new_n268), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT74), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n265), .A2(KEYINPUT74), .A3(G226), .A4(new_n268), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G97), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n265), .A2(G232), .A3(G1698), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n427), .A2(new_n428), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n272), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n260), .B1(new_n228), .B2(new_n263), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT13), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT13), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n432), .A2(new_n437), .A3(new_n434), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n424), .B1(new_n439), .B2(G169), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n437), .B1(new_n432), .B2(new_n434), .ZN(new_n441));
  AOI211_X1 g0241(.A(KEYINPUT13), .B(new_n433), .C1(new_n431), .C2(new_n272), .ZN(new_n442));
  OAI211_X1 g0242(.A(G169), .B(new_n424), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n436), .A2(G179), .A3(new_n438), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n423), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n441), .A2(new_n442), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n423), .B1(new_n447), .B2(G190), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT75), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n449), .B1(new_n439), .B2(G200), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n449), .B(G200), .C1(new_n441), .C2(new_n442), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n448), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n446), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n414), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G116), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n405), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n219), .A2(G33), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n318), .A2(new_n405), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n458), .B1(new_n461), .B2(new_n457), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G283), .ZN(new_n463));
  INV_X1    g0263(.A(G97), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n463), .B(new_n215), .C1(G33), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n457), .A2(G20), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(new_n284), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT20), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n465), .A2(KEYINPUT20), .A3(new_n284), .A4(new_n466), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(KEYINPUT85), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT85), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n467), .A2(new_n472), .A3(new_n468), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n462), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n256), .A2(G1), .ZN(new_n476));
  AND2_X1   g0276(.A1(KEYINPUT5), .A2(G41), .ZN(new_n477));
  NOR2_X1   g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(G270), .A3(new_n259), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT5), .B(G41), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n481), .A2(G274), .A3(new_n259), .A4(new_n476), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n332), .A2(new_n334), .A3(G264), .A4(G1698), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n332), .A2(new_n334), .A3(G257), .A4(new_n268), .ZN(new_n485));
  INV_X1    g0285(.A(G303), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n484), .B(new_n485), .C1(new_n486), .C2(new_n265), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n483), .B1(new_n272), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G190), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n475), .B(new_n489), .C1(new_n274), .C2(new_n488), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT21), .ZN(new_n491));
  INV_X1    g0291(.A(new_n483), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n487), .A2(new_n272), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G169), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n491), .B1(new_n475), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n474), .A2(G179), .A3(new_n488), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n474), .A2(KEYINPUT21), .A3(G169), .A4(new_n494), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n490), .A2(new_n496), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n405), .A2(G97), .ZN(new_n500));
  XNOR2_X1  g0300(.A(new_n500), .B(KEYINPUT80), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n501), .B1(new_n461), .B2(G97), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n291), .A2(new_n267), .ZN(new_n503));
  XNOR2_X1  g0303(.A(G97), .B(G107), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n505), .A2(new_n464), .A3(G107), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n503), .B1(new_n509), .B2(G20), .ZN(new_n510));
  OAI21_X1  g0310(.A(G107), .B1(new_n344), .B2(new_n345), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT79), .B1(new_n512), .B2(new_n284), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT79), .ZN(new_n514));
  AOI211_X1 g0314(.A(new_n514), .B(new_n318), .C1(new_n510), .C2(new_n511), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n502), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n479), .A2(G257), .A3(new_n259), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n332), .A2(new_n334), .A3(G250), .A4(G1698), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT81), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT81), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n265), .A2(new_n521), .A3(G250), .A4(G1698), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n265), .A2(KEYINPUT4), .A3(G244), .A4(new_n268), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n332), .A2(new_n334), .A3(G244), .A4(new_n268), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT4), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n523), .A2(new_n463), .A3(new_n524), .A4(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n518), .B1(new_n528), .B2(new_n272), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n393), .B1(new_n529), .B2(new_n482), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n520), .A2(new_n522), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n527), .A2(new_n524), .A3(new_n463), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n272), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(new_n482), .A3(new_n517), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(new_n308), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n516), .B1(new_n530), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n507), .B1(new_n505), .B2(new_n504), .ZN(new_n537));
  OAI22_X1  g0337(.A1(new_n537), .A2(new_n215), .B1(new_n267), .B2(new_n291), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n386), .B1(new_n330), .B2(new_n336), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n284), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g0340(.A(new_n540), .B(new_n514), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n529), .A2(G190), .A3(new_n482), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n534), .A2(G200), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .A4(new_n502), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n536), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT19), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n215), .B1(new_n429), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n229), .A2(new_n464), .A3(new_n386), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n332), .A2(new_n334), .A3(new_n215), .A4(G68), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n546), .B1(new_n288), .B2(new_n464), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n284), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n395), .A2(new_n397), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n405), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT83), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT83), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n553), .A2(new_n559), .A3(new_n556), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n558), .A2(new_n560), .B1(G87), .B2(new_n461), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n259), .A2(G274), .A3(new_n476), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT82), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n259), .A2(KEYINPUT82), .A3(G274), .A4(new_n476), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n476), .A2(new_n230), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n259), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n332), .A2(new_n334), .A3(G238), .A4(new_n268), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n332), .A2(new_n334), .A3(G244), .A4(G1698), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G33), .A2(G116), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n568), .B1(new_n272), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n573), .A2(KEYINPUT84), .A3(G190), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT84), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n572), .A2(new_n272), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n562), .A2(new_n563), .B1(new_n566), .B2(new_n259), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n576), .A2(G190), .A3(new_n565), .A4(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n565), .A3(new_n577), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n575), .A2(new_n578), .B1(new_n579), .B2(G200), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n561), .A2(new_n574), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n479), .A2(G264), .A3(new_n259), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n582), .A2(new_n482), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n332), .A2(new_n334), .A3(G257), .A4(G1698), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n332), .A2(new_n334), .A3(G250), .A4(new_n268), .ZN(new_n585));
  NAND2_X1  g0385(.A1(G33), .A2(G294), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n272), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n583), .A2(new_n308), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(G169), .B1(new_n583), .B2(new_n588), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT23), .B1(new_n215), .B2(G107), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT23), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(new_n386), .A3(G20), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n215), .A2(G33), .A3(G116), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT86), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT86), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n592), .A2(new_n594), .A3(new_n595), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n332), .A2(new_n334), .A3(new_n215), .A4(G87), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT22), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT22), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n265), .A2(new_n603), .A3(new_n215), .A4(G87), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT24), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT24), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n600), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n318), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n295), .A2(new_n386), .ZN(new_n611));
  NOR2_X1   g0411(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n611), .B2(new_n612), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n613), .A2(new_n615), .B1(new_n461), .B2(G107), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n591), .B1(new_n610), .B2(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n583), .A2(G190), .A3(new_n588), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n274), .B1(new_n583), .B2(new_n588), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n609), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n608), .B1(new_n600), .B2(new_n605), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n284), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n621), .A2(new_n624), .A3(new_n616), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n559), .B1(new_n553), .B2(new_n556), .ZN(new_n626));
  AOI211_X1 g0426(.A(KEYINPUT83), .B(new_n555), .C1(new_n552), .C2(new_n284), .ZN(new_n627));
  OAI22_X1  g0427(.A1(new_n626), .A2(new_n627), .B1(new_n398), .B2(new_n460), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n579), .A2(new_n393), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n573), .A2(new_n308), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n581), .A2(new_n618), .A3(new_n625), .A4(new_n631), .ZN(new_n632));
  NOR4_X1   g0432(.A1(new_n456), .A2(new_n499), .A3(new_n545), .A4(new_n632), .ZN(G372));
  NAND2_X1  g0433(.A1(new_n408), .A2(KEYINPUT91), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT91), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n394), .A2(new_n635), .A3(new_n406), .A4(new_n407), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n453), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n381), .B1(new_n637), .B2(new_n446), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n307), .B1(new_n638), .B2(new_n367), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n313), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n534), .A2(G169), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(new_n308), .B2(new_n534), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n643), .A2(new_n516), .A3(new_n581), .A4(new_n631), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT26), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n572), .A2(KEYINPUT88), .A3(new_n272), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(KEYINPUT88), .B1(new_n572), .B2(new_n272), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(G200), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n561), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT89), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT89), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n561), .A2(new_n651), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n653), .A2(new_n578), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT90), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n536), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n628), .A2(new_n630), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n650), .A2(new_n393), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n643), .A2(KEYINPUT90), .A3(new_n516), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n656), .A2(new_n658), .A3(new_n661), .A4(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n645), .B1(new_n663), .B2(KEYINPUT26), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n498), .A2(new_n497), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(new_n496), .A3(new_n618), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n666), .A2(new_n536), .A3(new_n544), .A4(new_n625), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n656), .A2(new_n661), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n661), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n641), .B1(new_n456), .B2(new_n670), .ZN(G369));
  NAND2_X1  g0471(.A1(new_n665), .A2(new_n496), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n404), .A2(new_n215), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G343), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n618), .A2(new_n625), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n618), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n678), .B(KEYINPUT92), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n475), .A2(new_n678), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n672), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n499), .B2(new_n685), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G330), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n678), .B1(new_n624), .B2(new_n616), .ZN(new_n692));
  OAI22_X1  g0492(.A1(new_n680), .A2(new_n692), .B1(new_n618), .B2(new_n678), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n684), .B1(new_n691), .B2(new_n694), .ZN(G399));
  NAND3_X1  g0495(.A1(new_n222), .A2(KEYINPUT93), .A3(new_n255), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT93), .B1(new_n222), .B2(new_n255), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n548), .A2(G116), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G1), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n212), .B2(new_n700), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  INV_X1    g0504(.A(new_n678), .ZN(new_n705));
  INV_X1    g0505(.A(new_n669), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n644), .A2(KEYINPUT26), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n663), .B2(KEYINPUT26), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n705), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT95), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(new_n710), .A3(KEYINPUT29), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n663), .A2(KEYINPUT26), .ZN(new_n712));
  INV_X1    g0512(.A(new_n707), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI211_X1 g0514(.A(KEYINPUT29), .B(new_n678), .C1(new_n714), .C2(new_n669), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT95), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n683), .B1(new_n664), .B2(new_n669), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT29), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n711), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n582), .A2(new_n482), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n722), .B1(new_n272), .B2(new_n587), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n573), .A2(new_n488), .A3(new_n723), .A4(G179), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n533), .A2(new_n517), .ZN(new_n725));
  OAI21_X1  g0525(.A(KEYINPUT30), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n646), .A2(new_n588), .A3(new_n583), .A4(new_n576), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n492), .A2(new_n493), .A3(G179), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n729), .A2(new_n730), .A3(new_n529), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n583), .A2(new_n588), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n494), .A2(new_n732), .A3(new_n308), .ZN(new_n733));
  INV_X1    g0533(.A(new_n649), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n568), .B1(new_n734), .B2(new_n647), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n726), .A2(new_n731), .B1(new_n534), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n678), .ZN(new_n738));
  XOR2_X1   g0538(.A(KEYINPUT94), .B(KEYINPUT31), .Z(new_n739));
  OR2_X1    g0539(.A1(new_n683), .A2(new_n739), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n738), .A2(KEYINPUT31), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n683), .ZN(new_n742));
  NOR4_X1   g0542(.A1(new_n545), .A2(new_n632), .A3(new_n499), .A4(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(G330), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n721), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n704), .B1(new_n745), .B2(G1), .ZN(G364));
  NOR2_X1   g0546(.A1(new_n294), .A2(G20), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n219), .B1(new_n747), .B2(G45), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n699), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G13), .A2(G33), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n688), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n214), .B1(G20), .B2(new_n393), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G179), .A2(G200), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(G20), .A3(new_n370), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G159), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(KEYINPUT32), .ZN(new_n761));
  AND2_X1   g0561(.A1(new_n760), .A2(KEYINPUT32), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n215), .B1(new_n757), .B2(G190), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n761), .B(new_n762), .C1(G97), .C2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n215), .A2(new_n308), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G200), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT99), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n370), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n768), .A2(G190), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n765), .B1(new_n770), .B2(new_n285), .C1(new_n202), .C2(new_n772), .ZN(new_n773));
  NOR4_X1   g0573(.A1(new_n215), .A2(new_n274), .A3(G179), .A4(G190), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n775), .A2(KEYINPUT100), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(KEYINPUT100), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G107), .ZN(new_n780));
  INV_X1    g0580(.A(new_n766), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n781), .A2(new_n370), .A3(G200), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n265), .B1(new_n783), .B2(new_n201), .ZN(new_n784));
  NOR4_X1   g0584(.A1(new_n215), .A2(new_n370), .A3(new_n274), .A4(G179), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n784), .B1(G87), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G190), .A2(G200), .ZN(new_n787));
  AND3_X1   g0587(.A1(new_n766), .A2(KEYINPUT98), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(KEYINPUT98), .B1(new_n766), .B2(new_n787), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n780), .B(new_n786), .C1(new_n267), .C2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n790), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n779), .A2(G283), .B1(G311), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n764), .A2(G294), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n265), .B1(new_n782), .B2(G322), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n785), .A2(G303), .B1(new_n759), .B2(G329), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n793), .A2(new_n794), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n769), .A2(G326), .ZN(new_n798));
  XOR2_X1   g0598(.A(KEYINPUT33), .B(G317), .Z(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n772), .B2(new_n799), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n773), .A2(new_n791), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n213), .A2(new_n256), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n222), .A2(new_n335), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT96), .Z(new_n804));
  OAI211_X1 g0604(.A(new_n802), .B(new_n804), .C1(new_n256), .C2(new_n249), .ZN(new_n805));
  INV_X1    g0605(.A(G355), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n222), .A2(new_n265), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n805), .B1(G116), .B2(new_n222), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n754), .A2(new_n756), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT97), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n756), .A2(new_n801), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n751), .B1(new_n755), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n687), .B(G330), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n813), .B1(new_n814), .B2(new_n751), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT101), .ZN(G396));
  OR2_X1    g0616(.A1(new_n756), .A2(new_n752), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n750), .B1(G77), .B2(new_n817), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n792), .A2(G159), .B1(G143), .B2(new_n782), .ZN(new_n819));
  INV_X1    g0619(.A(G137), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n819), .B1(new_n770), .B2(new_n820), .C1(new_n289), .C2(new_n772), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT34), .ZN(new_n822));
  INV_X1    g0622(.A(G132), .ZN(new_n823));
  INV_X1    g0623(.A(new_n785), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n265), .B1(new_n758), .B2(new_n823), .C1(new_n824), .C2(new_n285), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G58), .B2(new_n764), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n822), .B(new_n826), .C1(new_n202), .C2(new_n778), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n785), .A2(G107), .B1(new_n759), .B2(G311), .ZN(new_n828));
  INV_X1    g0628(.A(G294), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n828), .B(new_n335), .C1(new_n783), .C2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G97), .B2(new_n764), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n779), .A2(G87), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n831), .B(new_n832), .C1(new_n457), .C2(new_n790), .ZN(new_n833));
  INV_X1    g0633(.A(G283), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n834), .A2(new_n772), .B1(new_n770), .B2(new_n486), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n827), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n818), .B1(new_n836), .B2(new_n756), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n705), .A2(new_n406), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n634), .A2(new_n636), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n413), .B2(new_n838), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n837), .B1(new_n753), .B2(new_n840), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n683), .B(new_n840), .C1(new_n664), .C2(new_n669), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(KEYINPUT102), .ZN(new_n843));
  INV_X1    g0643(.A(new_n840), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n717), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n843), .B(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n744), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n751), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n846), .A2(new_n744), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n841), .B1(new_n848), .B2(new_n849), .ZN(G384));
  OR2_X1    g0650(.A1(new_n509), .A2(KEYINPUT35), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n509), .A2(KEYINPUT35), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n851), .A2(G116), .A3(new_n217), .A4(new_n852), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT36), .Z(new_n854));
  NAND3_X1  g0654(.A1(new_n213), .A2(G77), .A3(new_n319), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(G50), .B2(new_n202), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n219), .A2(G13), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n854), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OR2_X1    g0658(.A1(new_n408), .A2(new_n705), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n842), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n349), .A2(new_n676), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n381), .B2(new_n367), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n316), .B(new_n373), .C1(new_n361), .C2(new_n362), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n349), .B2(new_n358), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT37), .B1(new_n864), .B2(new_n861), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n363), .A2(new_n365), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n363), .A2(new_n677), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n866), .A2(new_n867), .A3(new_n868), .A4(new_n863), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n862), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n862), .A2(new_n870), .A3(KEYINPUT38), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n423), .A2(new_n705), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n454), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n446), .A2(new_n453), .A3(new_n876), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n860), .A2(new_n875), .A3(new_n880), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n446), .A2(new_n705), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT103), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n883), .A2(KEYINPUT39), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(KEYINPUT39), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n873), .B(new_n874), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n862), .A2(new_n870), .A3(KEYINPUT38), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT38), .B1(new_n862), .B2(new_n870), .ZN(new_n888));
  OAI22_X1  g0688(.A1(new_n887), .A2(new_n888), .B1(new_n883), .B2(KEYINPUT39), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n882), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n367), .A2(new_n676), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n881), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n456), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n720), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n641), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n894), .B(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT40), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n887), .A2(new_n888), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n536), .A2(new_n544), .ZN(new_n901));
  INV_X1    g0701(.A(new_n499), .ZN(new_n902));
  INV_X1    g0702(.A(new_n632), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n901), .A2(new_n902), .A3(new_n903), .A4(new_n683), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n736), .A2(new_n534), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n730), .B1(new_n729), .B2(new_n529), .ZN(new_n906));
  NOR4_X1   g0706(.A1(new_n725), .A2(new_n727), .A3(new_n728), .A4(KEYINPUT30), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(KEYINPUT31), .A3(new_n705), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n739), .B1(new_n737), .B2(new_n678), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n904), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(new_n880), .A3(new_n840), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n899), .B1(new_n900), .B2(new_n912), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n446), .A2(new_n453), .A3(new_n876), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n876), .B1(new_n446), .B2(new_n453), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n840), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n910), .A2(new_n909), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n743), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n875), .A2(new_n919), .A3(KEYINPUT40), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n913), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n456), .B2(new_n918), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n895), .A2(new_n913), .A3(new_n911), .A4(new_n920), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n923), .A3(G330), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n898), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n219), .B2(new_n747), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n898), .A2(new_n924), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n858), .B1(new_n926), .B2(new_n927), .ZN(G367));
  OAI21_X1  g0728(.A(new_n809), .B1(new_n222), .B2(new_n398), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n804), .B2(new_n245), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n785), .A2(G116), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT46), .ZN(new_n932));
  OAI221_X1 g0732(.A(new_n932), .B1(new_n386), .B2(new_n763), .C1(new_n772), .C2(new_n829), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n783), .A2(new_n486), .ZN(new_n934));
  AOI211_X1 g0734(.A(new_n265), .B(new_n934), .C1(G317), .C2(new_n759), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n779), .A2(G97), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n935), .B(new_n936), .C1(new_n834), .C2(new_n790), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n933), .B(new_n937), .C1(G311), .C2(new_n769), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n779), .A2(G77), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n285), .B2(new_n790), .ZN(new_n940));
  INV_X1    g0740(.A(G143), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n941), .A2(new_n770), .B1(new_n772), .B2(new_n322), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n782), .A2(G150), .B1(G137), .B2(new_n759), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n335), .B1(new_n785), .B2(G58), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n943), .B(new_n944), .C1(new_n202), .C2(new_n763), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n940), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n938), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT47), .Z(new_n948));
  AOI211_X1 g0748(.A(new_n751), .B(new_n930), .C1(new_n948), .C2(new_n756), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n561), .A2(new_n678), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n656), .A2(new_n661), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n661), .B2(new_n950), .ZN(new_n952));
  INV_X1    g0752(.A(new_n754), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n536), .A2(new_n683), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT104), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n742), .A2(new_n516), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n901), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n681), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT42), .Z(new_n961));
  AOI21_X1  g0761(.A(new_n618), .B1(new_n956), .B2(new_n958), .ZN(new_n962));
  INV_X1    g0762(.A(new_n536), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n683), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n961), .A2(new_n964), .B1(KEYINPUT43), .B2(new_n952), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n965), .B(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n691), .A2(new_n694), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n959), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n967), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n959), .A2(new_n684), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT45), .Z(new_n972));
  NOR2_X1   g0772(.A1(new_n959), .A2(new_n684), .ZN(new_n973));
  XNOR2_X1  g0773(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(new_n968), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n694), .A2(new_n679), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n680), .B2(new_n679), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n690), .B(new_n979), .Z(new_n980));
  OAI21_X1  g0780(.A(new_n745), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n699), .B(KEYINPUT41), .Z(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n749), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n954), .B1(new_n970), .B2(new_n984), .ZN(G387));
  INV_X1    g0785(.A(new_n980), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n694), .A2(new_n754), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n807), .A2(new_n701), .B1(G107), .B2(new_n222), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n242), .A2(G45), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT106), .ZN(new_n990));
  INV_X1    g0790(.A(new_n804), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n287), .A2(G50), .ZN(new_n992));
  XNOR2_X1  g0792(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n992), .B(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n701), .ZN(new_n995));
  AOI211_X1 g0795(.A(G45), .B(new_n995), .C1(G68), .C2(G77), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n991), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n988), .B1(new_n990), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n750), .B1(new_n998), .B2(new_n810), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT108), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n335), .B1(new_n759), .B2(G150), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n936), .B(new_n1001), .C1(new_n267), .C2(new_n824), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT109), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n782), .A2(G50), .B1(new_n554), .B2(new_n764), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n202), .B2(new_n790), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G159), .B2(new_n769), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1003), .B(new_n1006), .C1(new_n287), .C2(new_n772), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n265), .B1(new_n759), .B2(G326), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n824), .A2(new_n829), .B1(new_n763), .B2(new_n834), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n771), .A2(G311), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n792), .A2(G303), .B1(G317), .B2(new_n782), .ZN(new_n1011));
  INV_X1    g0811(.A(G322), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1010), .B(new_n1011), .C1(new_n770), .C2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT48), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1009), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n1014), .B2(new_n1013), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT49), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1008), .B1(new_n457), .B2(new_n778), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1007), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1000), .B1(new_n756), .B2(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n986), .A2(new_n749), .B1(new_n987), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n745), .A2(new_n986), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n699), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n745), .A2(new_n986), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1022), .B1(new_n1024), .B2(new_n1025), .ZN(G393));
  AND2_X1   g0826(.A1(new_n977), .A2(new_n1023), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n699), .B1(new_n977), .B2(new_n1023), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n809), .B1(new_n464), .B2(new_n222), .C1(new_n991), .C2(new_n252), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n750), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT110), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n335), .B1(new_n758), .B2(new_n1012), .C1(new_n824), .C2(new_n834), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n780), .B1(new_n829), .B2(new_n790), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1033), .B(new_n1034), .C1(G116), .C2(new_n764), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n769), .A2(G317), .B1(G311), .B2(new_n782), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT52), .Z(new_n1037));
  OAI211_X1 g0837(.A(new_n1035), .B(new_n1037), .C1(new_n486), .C2(new_n772), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n265), .B1(new_n758), .B2(new_n941), .C1(new_n824), .C2(new_n202), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n832), .B1(new_n287), .B2(new_n790), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(G77), .C2(new_n764), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n770), .A2(new_n289), .B1(new_n322), .B2(new_n783), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1041), .B(new_n1044), .C1(new_n285), .C2(new_n772), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1038), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(KEYINPUT112), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n756), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1047), .A2(KEYINPUT112), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1032), .B1(new_n953), .B2(new_n959), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n977), .B2(new_n748), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1029), .A2(new_n1052), .ZN(G390));
  NAND3_X1  g0853(.A1(new_n886), .A2(new_n752), .A3(new_n889), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n287), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n750), .B1(new_n1055), .B2(new_n817), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n785), .A2(G150), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1057), .B(new_n1058), .Z(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G159), .B2(new_n764), .ZN(new_n1060));
  INV_X1    g0860(.A(G128), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1060), .B1(new_n770), .B2(new_n1061), .C1(new_n820), .C2(new_n772), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n265), .B1(new_n783), .B2(new_n823), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G125), .B2(new_n759), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(KEYINPUT54), .B(G143), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1064), .B1(new_n285), .B2(new_n778), .C1(new_n790), .C2(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n783), .A2(new_n457), .B1(new_n829), .B2(new_n758), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n265), .B(new_n1067), .C1(G87), .C2(new_n785), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n779), .A2(G68), .B1(G97), .B2(new_n792), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n267), .C2(new_n763), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n386), .A2(new_n772), .B1(new_n770), .B2(new_n834), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n1062), .A2(new_n1066), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1056), .B1(new_n1072), .B2(new_n756), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1054), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n709), .A2(new_n840), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1075), .A2(new_n859), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n880), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n875), .B(new_n882), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1077), .B1(new_n842), .B2(new_n859), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n882), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n886), .B(new_n889), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n744), .A2(new_n844), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n880), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n919), .A2(G330), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1074), .B1(new_n1090), .B2(new_n748), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n911), .A2(G330), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n456), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n896), .A2(new_n641), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1087), .B1(new_n880), .B2(new_n1084), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n860), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1077), .B1(new_n1092), .B2(new_n844), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1085), .A2(new_n1075), .A3(new_n1098), .A4(new_n859), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1095), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1090), .A2(KEYINPUT113), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(KEYINPUT113), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1088), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n700), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1091), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(G378));
  OAI21_X1  g0907(.A(new_n750), .B1(G50), .B2(new_n817), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n265), .A2(G41), .ZN(new_n1109));
  AOI211_X1 g0909(.A(G50), .B(new_n1109), .C1(new_n331), .C2(new_n255), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n782), .A2(G107), .B1(G283), .B2(new_n759), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1111), .B(new_n1109), .C1(new_n267), .C2(new_n824), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G68), .B2(new_n764), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G97), .A2(new_n771), .B1(new_n769), .B2(G116), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n792), .A2(new_n554), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n779), .A2(G58), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT58), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1110), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(KEYINPUT116), .B(G124), .ZN(new_n1120));
  AOI211_X1 g0920(.A(G33), .B(G41), .C1(new_n759), .C2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n824), .A2(new_n1065), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT115), .Z(new_n1123));
  AOI22_X1  g0923(.A1(new_n782), .A2(G128), .B1(G150), .B2(new_n764), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1123), .B(new_n1124), .C1(new_n820), .C2(new_n790), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n772), .A2(new_n823), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1125), .B(new_n1126), .C1(G125), .C2(new_n769), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT59), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1121), .B1(new_n322), .B2(new_n778), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1127), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1130), .A2(KEYINPUT59), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1119), .B1(new_n1118), .B2(new_n1117), .C1(new_n1129), .C2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1108), .B1(new_n1132), .B2(new_n756), .ZN(new_n1133));
  XOR2_X1   g0933(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n307), .A2(new_n313), .A3(new_n1135), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n301), .A2(new_n303), .B1(KEYINPUT10), .B2(new_n305), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1134), .B1(new_n1137), .B2(new_n312), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n299), .A2(new_n677), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT117), .Z(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1136), .A2(new_n1138), .A3(new_n1141), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1143), .A2(new_n752), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1133), .A2(new_n1145), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT118), .Z(new_n1147));
  NAND3_X1  g0947(.A1(new_n913), .A2(G330), .A3(new_n920), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT119), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1136), .A2(new_n1138), .A3(new_n1141), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1141), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1143), .A2(KEYINPUT119), .A3(new_n1144), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1148), .A2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n913), .A2(new_n1153), .A3(new_n920), .A4(G330), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n893), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT122), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n893), .A2(KEYINPUT122), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT120), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1155), .A2(KEYINPUT120), .A3(new_n1156), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(KEYINPUT121), .B1(new_n1167), .B2(new_n894), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1155), .A2(KEYINPUT120), .A3(new_n1156), .ZN(new_n1169));
  AOI21_X1  g0969(.A(KEYINPUT120), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1170));
  OAI211_X1 g0970(.A(KEYINPUT121), .B(new_n894), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1162), .B1(new_n1168), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1147), .B1(new_n1173), .B2(new_n749), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT57), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n894), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT121), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1161), .B1(new_n1178), .B2(new_n1171), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1094), .B1(new_n1104), .B2(new_n1100), .ZN(new_n1180));
  OAI211_X1 g0980(.A(KEYINPUT123), .B(new_n1175), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1100), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1095), .B1(new_n1090), .B2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1163), .B(new_n893), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1184), .A2(new_n1175), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n700), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1181), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1173), .A2(new_n1183), .ZN(new_n1188));
  AOI21_X1  g0988(.A(KEYINPUT123), .B1(new_n1188), .B2(new_n1175), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1174), .B1(new_n1187), .B2(new_n1189), .ZN(G375));
  NAND2_X1  g0990(.A1(new_n1094), .A2(new_n1182), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1101), .A2(new_n983), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1077), .A2(new_n752), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n750), .B1(G68), .B2(new_n817), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(G116), .A2(new_n771), .B1(new_n769), .B2(G294), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n785), .A2(G97), .B1(new_n759), .B2(G303), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1196), .B(new_n335), .C1(new_n783), .C2(new_n834), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n554), .B2(new_n764), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n792), .A2(G107), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1195), .A2(new_n1198), .A3(new_n939), .A4(new_n1199), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n824), .A2(new_n322), .B1(new_n1061), .B2(new_n758), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n265), .B1(new_n783), .B2(new_n820), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(G50), .C2(new_n764), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1203), .B(new_n1116), .C1(new_n289), .C2(new_n790), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n823), .A2(new_n770), .B1(new_n772), .B2(new_n1065), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1200), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1194), .B1(new_n1206), .B2(new_n756), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1100), .A2(new_n749), .B1(new_n1193), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1192), .A2(new_n1208), .ZN(G381));
  NOR2_X1   g1009(.A1(new_n1029), .A2(new_n1052), .ZN(new_n1210));
  INV_X1    g1010(.A(G384), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NOR4_X1   g1012(.A1(new_n1212), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n984), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n969), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n967), .B(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1213), .A2(new_n1217), .A3(new_n954), .ZN(new_n1218));
  OR3_X1    g1018(.A1(new_n1218), .A2(G375), .A3(G378), .ZN(G407));
  INV_X1    g1019(.A(G343), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(G213), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1106), .A2(new_n1222), .ZN(new_n1223));
  OAI211_X1 g1023(.A(G407), .B(G213), .C1(G375), .C2(new_n1223), .ZN(G409));
  OAI211_X1 g1024(.A(G378), .B(new_n1174), .C1(new_n1187), .C2(new_n1189), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1188), .A2(new_n982), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1147), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1184), .B2(new_n748), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1106), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1222), .B1(new_n1225), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT62), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n699), .B1(new_n1094), .B2(new_n1182), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT60), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1232), .B1(new_n1233), .B2(new_n1191), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1094), .A2(KEYINPUT60), .A3(new_n1182), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(KEYINPUT124), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT124), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1094), .A2(new_n1182), .A3(new_n1237), .A4(KEYINPUT60), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1236), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1234), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(KEYINPUT125), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT125), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1234), .A2(new_n1239), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1241), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(G384), .B1(new_n1244), .B2(new_n1208), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1234), .A2(new_n1239), .A3(new_n1242), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1242), .B1(new_n1234), .B2(new_n1239), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G384), .B(new_n1208), .C1(new_n1246), .C2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1245), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1230), .A2(new_n1231), .A3(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1222), .A2(G2897), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n1245), .B2(new_n1249), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1208), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1211), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(new_n1248), .A3(new_n1253), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1255), .A2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1251), .B(new_n1252), .C1(new_n1230), .C2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1231), .B1(new_n1230), .B2(new_n1250), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1217), .A2(G390), .A3(new_n954), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G387), .A2(new_n1210), .ZN(new_n1263));
  XOR2_X1   g1063(.A(G393), .B(G396), .Z(new_n1264));
  AND3_X1   g1064(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1264), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n1260), .A2(new_n1261), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1265), .A2(new_n1266), .A3(KEYINPUT61), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n1230), .B2(new_n1259), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT63), .B1(new_n1230), .B2(new_n1250), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1225), .A2(new_n1229), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1257), .A2(KEYINPUT63), .A3(new_n1248), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(new_n1221), .A3(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT126), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1230), .A2(KEYINPUT126), .A3(new_n1273), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT127), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1271), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1279), .B1(new_n1271), .B2(new_n1278), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1267), .B1(new_n1280), .B2(new_n1281), .ZN(G405));
  NAND2_X1  g1082(.A1(G375), .A2(new_n1106), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1225), .ZN(new_n1284));
  XOR2_X1   g1084(.A(new_n1284), .B(new_n1250), .Z(new_n1285));
  NOR2_X1   g1085(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1285), .B(new_n1286), .ZN(G402));
endmodule


