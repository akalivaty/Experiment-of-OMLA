//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  AOI22_X1  g0007(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G116), .ZN(new_n209));
  INV_X1    g0009(.A(G270), .ZN(new_n210));
  OAI21_X1  g0010(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G68), .A2(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n212), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n211), .B(new_n216), .C1(G97), .C2(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G1), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n202), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(new_n219), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G13), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n220), .A2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT0), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n222), .A2(new_n227), .A3(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT64), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G68), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT65), .ZN(new_n244));
  XOR2_X1   g0044(.A(G50), .B(G58), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n225), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT66), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n218), .A2(G13), .A3(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n218), .A2(G20), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n254), .A2(G50), .A3(new_n255), .A4(new_n256), .ZN(new_n257));
  OR2_X1    g0057(.A1(new_n255), .A2(G50), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(KEYINPUT70), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(KEYINPUT70), .B1(new_n257), .B2(new_n258), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n263));
  INV_X1    g0063(.A(G150), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G58), .ZN(new_n267));
  OR3_X1    g0067(.A1(new_n267), .A2(KEYINPUT68), .A3(KEYINPUT8), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT68), .B1(new_n267), .B2(KEYINPUT8), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT67), .B(G58), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT8), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n268), .B(new_n269), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  OAI21_X1  g0074(.A(KEYINPUT69), .B1(new_n274), .B2(G20), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT69), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(new_n219), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  OAI221_X1 g0078(.A(new_n263), .B1(new_n264), .B2(new_n266), .C1(new_n273), .C2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n254), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT9), .B1(new_n262), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n261), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n259), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT9), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(new_n286), .A3(new_n281), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n274), .ZN(new_n290));
  NAND2_X1  g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G223), .A2(G1698), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G222), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n292), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G41), .ZN(new_n297));
  OAI211_X1 g0097(.A(G1), .B(G13), .C1(new_n274), .C2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n296), .B(new_n299), .C1(G77), .C2(new_n292), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n218), .B1(G41), .B2(G45), .ZN(new_n301));
  INV_X1    g0101(.A(G274), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n298), .A2(new_n301), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n300), .B(new_n303), .C1(new_n215), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G200), .ZN(new_n306));
  INV_X1    g0106(.A(G190), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n306), .B1(new_n307), .B2(new_n305), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n288), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n288), .A2(KEYINPUT74), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n309), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT74), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n283), .A2(new_n314), .A3(new_n287), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT10), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT75), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n313), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n317), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n308), .B1(new_n288), .B2(KEYINPUT74), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT75), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n311), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n305), .A2(G179), .ZN(new_n324));
  XOR2_X1   g0124(.A(new_n324), .B(KEYINPUT71), .Z(new_n325));
  NAND2_X1  g0125(.A1(new_n285), .A2(new_n281), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n305), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n325), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G238), .A2(G1698), .ZN(new_n330));
  INV_X1    g0130(.A(G232), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n292), .B(new_n330), .C1(new_n331), .C2(G1698), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n332), .B(new_n299), .C1(G107), .C2(new_n292), .ZN(new_n333));
  INV_X1    g0133(.A(new_n304), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G244), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n303), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT72), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT72), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n333), .A2(new_n338), .A3(new_n303), .A4(new_n335), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G179), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G20), .A2(G77), .ZN(new_n343));
  XNOR2_X1  g0143(.A(KEYINPUT8), .B(G58), .ZN(new_n344));
  XOR2_X1   g0144(.A(KEYINPUT15), .B(G87), .Z(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  OAI221_X1 g0146(.A(new_n343), .B1(new_n266), .B2(new_n344), .C1(new_n346), .C2(new_n278), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n347), .A2(new_n252), .ZN(new_n348));
  INV_X1    g0148(.A(new_n252), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n349), .A2(G77), .A3(new_n256), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT73), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n255), .A2(G77), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n348), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n342), .B(new_n354), .C1(G169), .C2(new_n340), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n340), .A2(G190), .ZN(new_n356));
  INV_X1    g0156(.A(G200), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n356), .B(new_n353), .C1(new_n357), .C2(new_n340), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n323), .A2(new_n329), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n270), .A2(G68), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n202), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n362), .A2(G20), .B1(G159), .B2(new_n265), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n290), .A2(new_n219), .A3(new_n291), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT7), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g0166(.A1(KEYINPUT3), .A2(G33), .ZN(new_n367));
  NOR2_X1   g0167(.A1(KEYINPUT3), .A2(G33), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n367), .A2(new_n368), .A3(G20), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT79), .B1(new_n369), .B2(KEYINPUT7), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT79), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n364), .A2(new_n371), .A3(new_n365), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n366), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G68), .ZN(new_n374));
  OAI211_X1 g0174(.A(KEYINPUT16), .B(new_n363), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n252), .ZN(new_n376));
  XOR2_X1   g0176(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n377));
  NAND2_X1  g0177(.A1(new_n364), .A2(new_n365), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n367), .A2(new_n368), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n379), .A2(KEYINPUT7), .A3(new_n219), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(new_n380), .A3(KEYINPUT81), .ZN(new_n381));
  OR3_X1    g0181(.A1(new_n364), .A2(KEYINPUT81), .A3(new_n365), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(new_n382), .A3(G68), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n377), .B1(new_n383), .B2(new_n363), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT82), .B1(new_n376), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT84), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n304), .B2(new_n331), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n298), .A2(KEYINPUT84), .A3(G232), .A4(new_n301), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n387), .A2(new_n303), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n215), .A2(G1698), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n292), .B(new_n390), .C1(G223), .C2(G1698), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G87), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n298), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n357), .B1(new_n389), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT85), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n389), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n393), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n387), .A2(KEYINPUT85), .A3(new_n303), .A4(new_n388), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n394), .B1(new_n399), .B2(G190), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n383), .A2(new_n363), .ZN(new_n401));
  INV_X1    g0201(.A(new_n377), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT82), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n403), .A2(new_n404), .A3(new_n252), .A4(new_n375), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n254), .A2(new_n255), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n272), .A2(new_n256), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n406), .A2(new_n407), .B1(new_n255), .B2(new_n272), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT83), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n408), .B(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n385), .A2(new_n400), .A3(new_n405), .A4(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT17), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n385), .A2(new_n405), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n414), .A2(KEYINPUT17), .A3(new_n400), .A4(new_n410), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n385), .A2(new_n410), .A3(new_n405), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n396), .A2(new_n341), .A3(new_n397), .A4(new_n398), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n327), .B1(new_n389), .B2(new_n393), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n416), .A2(KEYINPUT18), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT18), .B1(new_n416), .B2(new_n420), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n413), .B(new_n415), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(G33), .A2(G97), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n292), .B1(G232), .B2(new_n294), .ZN(new_n426));
  NOR2_X1   g0226(.A1(G226), .A2(G1698), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n428), .A2(new_n299), .B1(G238), .B2(new_n334), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT13), .ZN(new_n430));
  XOR2_X1   g0230(.A(new_n303), .B(KEYINPUT76), .Z(new_n431));
  NAND3_X1  g0231(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT77), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n430), .B1(new_n429), .B2(new_n431), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI211_X1 g0236(.A(KEYINPUT77), .B(new_n430), .C1(new_n429), .C2(new_n431), .ZN(new_n437));
  OAI21_X1  g0237(.A(G179), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(G169), .B1(new_n433), .B2(new_n435), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT78), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n439), .B1(new_n440), .B2(KEYINPUT14), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(KEYINPUT14), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n440), .A2(KEYINPUT14), .ZN(new_n443));
  OAI211_X1 g0243(.A(G169), .B(new_n443), .C1(new_n433), .C2(new_n435), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n438), .A2(new_n441), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(G77), .ZN(new_n446));
  OAI22_X1  g0246(.A1(new_n278), .A2(new_n446), .B1(new_n214), .B2(new_n266), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n219), .A2(G68), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n280), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT11), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n349), .A2(G68), .A3(new_n256), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n449), .B2(new_n450), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n448), .A2(new_n218), .A3(G13), .ZN(new_n454));
  XOR2_X1   g0254(.A(new_n454), .B(KEYINPUT12), .Z(new_n455));
  NOR3_X1   g0255(.A1(new_n451), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n445), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(G190), .B1(new_n436), .B2(new_n437), .ZN(new_n459));
  OAI21_X1  g0259(.A(G200), .B1(new_n433), .B2(new_n435), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n460), .A3(new_n456), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n424), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n360), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n218), .A2(new_n209), .A3(G13), .A4(G20), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n218), .A2(G33), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n349), .A2(G116), .A3(new_n255), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G283), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n467), .B(new_n219), .C1(G33), .C2(new_n204), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n468), .B(new_n252), .C1(new_n219), .C2(G116), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT20), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n469), .A2(new_n470), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n464), .B(new_n466), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT5), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT87), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n475), .B1(new_n476), .B2(G41), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n297), .A2(KEYINPUT87), .A3(KEYINPUT5), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n477), .A2(new_n478), .A3(new_n218), .A4(G45), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(new_n302), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n292), .A2(G257), .A3(new_n294), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT89), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n379), .A2(G303), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n292), .A2(KEYINPUT89), .A3(G257), .A4(new_n294), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n292), .A2(G264), .A3(G1698), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n483), .A2(new_n484), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n480), .B1(new_n487), .B2(new_n299), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n479), .A2(new_n298), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G270), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n474), .B1(new_n491), .B2(new_n307), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n357), .B1(new_n488), .B2(new_n490), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n252), .A2(new_n253), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT66), .B1(new_n251), .B2(new_n225), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n255), .B(new_n465), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(new_n205), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT24), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n219), .B(G87), .C1(new_n367), .C2(new_n368), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT22), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT22), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n292), .A2(new_n503), .A3(new_n219), .A4(G87), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n274), .A2(new_n209), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n219), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n219), .A2(G107), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n508), .B(KEYINPUT23), .ZN(new_n509));
  AND4_X1   g0309(.A1(new_n500), .A2(new_n505), .A3(new_n507), .A4(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n502), .A2(new_n504), .B1(new_n219), .B2(new_n506), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n500), .B1(new_n511), .B2(new_n509), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n252), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n499), .B1(new_n513), .B2(KEYINPUT90), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n255), .A2(G107), .ZN(new_n515));
  XNOR2_X1  g0315(.A(KEYINPUT91), .B(KEYINPUT25), .ZN(new_n516));
  XNOR2_X1  g0316(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT90), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n518), .B(new_n252), .C1(new_n510), .C2(new_n512), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n514), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n292), .A2(G257), .A3(G1698), .ZN(new_n521));
  INV_X1    g0321(.A(G294), .ZN(new_n522));
  OAI21_X1  g0322(.A(G250), .B1(new_n367), .B2(new_n368), .ZN(new_n523));
  OAI221_X1 g0323(.A(new_n521), .B1(new_n274), .B2(new_n522), .C1(G1698), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n299), .ZN(new_n525));
  INV_X1    g0325(.A(new_n480), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n489), .A2(G264), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n327), .ZN(new_n529));
  INV_X1    g0329(.A(new_n528), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n341), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n520), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n491), .A2(KEYINPUT21), .A3(G169), .A4(new_n473), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n488), .A2(G179), .A3(new_n473), .A4(new_n490), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n327), .B1(new_n488), .B2(new_n490), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT21), .B1(new_n536), .B2(new_n473), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n532), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n345), .A2(new_n255), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n275), .A2(new_n277), .A3(G97), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT19), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n219), .B1(new_n425), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(G87), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n544), .A2(new_n204), .A3(new_n205), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n541), .A2(new_n542), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n292), .A2(new_n219), .A3(G68), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n540), .B1(new_n548), .B2(new_n252), .ZN(new_n549));
  OR2_X1    g0349(.A1(new_n498), .A2(new_n346), .ZN(new_n550));
  OR2_X1    g0350(.A1(G238), .A2(G1698), .ZN(new_n551));
  OAI221_X1 g0351(.A(new_n551), .B1(G244), .B2(new_n294), .C1(new_n367), .C2(new_n368), .ZN(new_n552));
  INV_X1    g0352(.A(new_n506), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n299), .ZN(new_n555));
  AOI21_X1  g0355(.A(G274), .B1(KEYINPUT88), .B2(G250), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n218), .A2(G45), .ZN(new_n557));
  OR2_X1    g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT88), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n559), .A3(G250), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n299), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n549), .A2(new_n550), .B1(new_n563), .B2(new_n327), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n555), .A2(new_n341), .A3(new_n562), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n357), .B1(new_n555), .B2(new_n562), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n298), .B1(new_n552), .B2(new_n553), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n567), .A2(new_n561), .A3(new_n307), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n349), .B1(new_n546), .B2(new_n547), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n498), .A2(new_n544), .ZN(new_n571));
  NOR3_X1   g0371(.A1(new_n570), .A2(new_n571), .A3(new_n540), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n564), .A2(new_n565), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n528), .A2(G200), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n514), .A2(new_n517), .A3(new_n519), .A4(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n528), .A2(new_n307), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n573), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n255), .A2(G97), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n381), .A2(new_n382), .A3(G107), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n205), .A2(KEYINPUT6), .A3(G97), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G97), .A2(G107), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n206), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n580), .B1(new_n582), .B2(KEYINPUT6), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G20), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n265), .A2(G77), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n579), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n578), .B1(new_n586), .B2(new_n252), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n498), .A2(new_n204), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n489), .A2(G257), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT4), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n292), .A2(G244), .A3(new_n294), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n591), .B1(new_n592), .B2(KEYINPUT86), .ZN(new_n593));
  INV_X1    g0393(.A(new_n467), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n591), .A2(KEYINPUT86), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n294), .B1(new_n523), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n595), .B1(new_n292), .B2(G244), .ZN(new_n597));
  NOR4_X1   g0397(.A1(new_n593), .A2(new_n594), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n526), .B(new_n590), .C1(new_n598), .C2(new_n298), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n587), .A2(new_n589), .B1(new_n599), .B2(new_n327), .ZN(new_n600));
  INV_X1    g0400(.A(new_n593), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n596), .A2(new_n594), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n299), .B1(new_n603), .B2(new_n597), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n604), .A2(new_n341), .A3(new_n526), .A4(new_n590), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n599), .A2(G200), .ZN(new_n607));
  AOI211_X1 g0407(.A(new_n578), .B(new_n588), .C1(new_n586), .C2(new_n252), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n607), .B(new_n608), .C1(new_n307), .C2(new_n599), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n577), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n463), .A2(new_n495), .A3(new_n539), .A4(new_n611), .ZN(new_n612));
  XNOR2_X1  g0412(.A(new_n612), .B(KEYINPUT92), .ZN(G372));
  OAI21_X1  g0413(.A(KEYINPUT93), .B1(new_n535), .B2(new_n537), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n491), .A2(G169), .A3(new_n473), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT21), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT93), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n617), .A2(new_n618), .A3(new_n534), .A4(new_n533), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n532), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n611), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n564), .A2(new_n565), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n587), .A2(new_n589), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n599), .A2(new_n327), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n573), .A2(new_n624), .A3(new_n625), .A4(new_n605), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n600), .A2(KEYINPUT26), .A3(new_n605), .A4(new_n573), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n623), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n622), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n463), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n329), .ZN(new_n633));
  INV_X1    g0433(.A(new_n355), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n445), .A2(new_n457), .B1(new_n461), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n415), .A2(new_n413), .ZN(new_n636));
  OAI22_X1  g0436(.A1(new_n635), .A2(new_n636), .B1(new_n422), .B2(new_n421), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n633), .B1(new_n323), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n632), .A2(new_n638), .ZN(G369));
  NOR2_X1   g0439(.A1(new_n228), .A2(G20), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n218), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(G213), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(G343), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n538), .B(new_n495), .C1(new_n474), .C2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n474), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n614), .A2(new_n619), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT94), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n532), .A2(new_n646), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n520), .A2(new_n646), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n576), .B2(new_n575), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n654), .B1(new_n656), .B2(new_n532), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n653), .A2(G330), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g0458(.A(new_n658), .B(KEYINPUT95), .Z(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n538), .A2(new_n646), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n654), .B1(new_n657), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n660), .A2(new_n662), .ZN(G399));
  NOR2_X1   g0463(.A1(new_n229), .A2(G41), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n545), .A2(G116), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G1), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n223), .B2(new_n665), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT28), .ZN(new_n669));
  AOI211_X1 g0469(.A(KEYINPUT29), .B(new_n646), .C1(new_n622), .C2(new_n630), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT96), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n630), .A2(new_n671), .ZN(new_n672));
  AOI211_X1 g0472(.A(KEYINPUT96), .B(new_n623), .C1(new_n628), .C2(new_n629), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n539), .A2(KEYINPUT97), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n532), .A2(new_n538), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT97), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n675), .A2(new_n611), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n646), .B1(new_n674), .B2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n670), .B1(new_n681), .B2(KEYINPUT29), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n611), .A2(new_n539), .A3(new_n495), .A4(new_n647), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n491), .A2(new_n341), .A3(new_n563), .ZN(new_n684));
  INV_X1    g0484(.A(new_n599), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n684), .A2(new_n685), .A3(new_n527), .A4(new_n525), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT30), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n685), .A2(new_n530), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(new_n341), .A3(new_n491), .A4(new_n563), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n686), .A2(new_n687), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n646), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n683), .A2(KEYINPUT31), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT31), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n692), .A2(new_n695), .A3(new_n646), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n682), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n669), .B1(new_n700), .B2(G1), .ZN(G364));
  NAND2_X1  g0501(.A1(new_n640), .A2(G45), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n665), .A2(G1), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n653), .A2(G330), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n704), .A2(KEYINPUT98), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(KEYINPUT98), .ZN(new_n706));
  OAI221_X1 g0506(.A(new_n703), .B1(G330), .B2(new_n653), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n703), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n219), .A2(new_n341), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT99), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(G190), .A2(G200), .ZN(new_n712));
  OAI21_X1  g0512(.A(KEYINPUT99), .B1(new_n219), .B2(new_n341), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(G311), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n219), .A2(G179), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n712), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G329), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n307), .A2(G200), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n711), .A2(new_n722), .A3(new_n713), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(G322), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n721), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n718), .A2(new_n307), .A3(G200), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI211_X1 g0528(.A(new_n717), .B(new_n726), .C1(G283), .C2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n709), .A2(G200), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n307), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G326), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n718), .A2(G190), .A3(G200), .ZN(new_n733));
  INV_X1    g0533(.A(G303), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n379), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n735), .A2(KEYINPUT101), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n722), .A2(new_n341), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n709), .A2(new_n307), .A3(G200), .ZN(new_n740));
  XOR2_X1   g0540(.A(KEYINPUT33), .B(G317), .Z(new_n741));
  OAI22_X1  g0541(.A1(new_n739), .A2(new_n522), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n742), .B1(KEYINPUT101), .B2(new_n735), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n729), .A2(new_n732), .A3(new_n736), .A4(new_n743), .ZN(new_n744));
  OAI221_X1 g0544(.A(new_n292), .B1(new_n733), .B2(new_n544), .C1(new_n205), .C2(new_n727), .ZN(new_n745));
  XOR2_X1   g0545(.A(new_n745), .B(KEYINPUT100), .Z(new_n746));
  OAI22_X1  g0546(.A1(new_n715), .A2(new_n446), .B1(new_n374), .B2(new_n740), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(new_n270), .B2(new_n723), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n720), .A2(G159), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n749), .A2(KEYINPUT32), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n749), .A2(KEYINPUT32), .B1(new_n738), .B2(G97), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n746), .A2(new_n748), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n731), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n214), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n744), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n225), .B1(G20), .B2(new_n327), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n756), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n229), .A2(new_n292), .ZN(new_n761));
  INV_X1    g0561(.A(G45), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n224), .A2(new_n762), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n761), .B(new_n763), .C1(new_n246), .C2(new_n762), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n230), .A2(G355), .A3(new_n292), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n764), .B(new_n765), .C1(G116), .C2(new_n230), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n755), .A2(new_n756), .B1(new_n760), .B2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n759), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n708), .B(new_n767), .C1(new_n651), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n707), .A2(new_n769), .ZN(G396));
  INV_X1    g0570(.A(new_n270), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n739), .A2(new_n771), .B1(new_n727), .B2(new_n374), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n292), .B1(new_n733), .B2(new_n214), .ZN(new_n773));
  INV_X1    g0573(.A(new_n740), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n723), .A2(G143), .B1(G150), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G137), .ZN(new_n776));
  INV_X1    g0576(.A(G159), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n775), .B1(new_n776), .B2(new_n753), .C1(new_n777), .C2(new_n715), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT104), .Z(new_n779));
  AOI211_X1 g0579(.A(new_n772), .B(new_n773), .C1(new_n779), .C2(KEYINPUT34), .ZN(new_n780));
  INV_X1    g0580(.A(G132), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n780), .B1(KEYINPUT34), .B2(new_n779), .C1(new_n781), .C2(new_n719), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n739), .A2(new_n204), .B1(new_n716), .B2(new_n719), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n209), .A2(new_n715), .B1(new_n724), .B2(new_n522), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n783), .B(new_n784), .C1(G303), .C2(new_n731), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n728), .A2(G87), .ZN(new_n786));
  INV_X1    g0586(.A(G283), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n740), .A2(KEYINPUT102), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n740), .A2(KEYINPUT102), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n785), .B(new_n786), .C1(new_n787), .C2(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n379), .B1(new_n733), .B2(new_n205), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT103), .Z(new_n793));
  OAI21_X1  g0593(.A(new_n782), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n756), .A2(new_n757), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n794), .A2(new_n756), .B1(new_n446), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n354), .A2(new_n646), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n355), .A2(new_n358), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(KEYINPUT105), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT105), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n355), .A2(new_n358), .A3(new_n800), .A4(new_n797), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n799), .A2(new_n801), .B1(new_n634), .B2(new_n646), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n796), .B(new_n708), .C1(new_n758), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n799), .A2(new_n801), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n631), .A2(new_n647), .A3(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n802), .B(KEYINPUT106), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n646), .B1(new_n622), .B2(new_n630), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n699), .B(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n804), .B1(new_n811), .B2(new_n708), .ZN(G384));
  INV_X1    g0612(.A(new_n461), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n457), .B(new_n646), .C1(new_n813), .C2(new_n445), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n457), .A2(new_n646), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n458), .A2(new_n461), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n802), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  AND4_X1   g0617(.A1(KEYINPUT40), .A2(new_n817), .A3(new_n694), .A4(new_n696), .ZN(new_n818));
  INV_X1    g0618(.A(new_n644), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n201), .B1(new_n270), .B2(G68), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n820), .A2(new_n219), .B1(new_n777), .B2(new_n266), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n370), .A2(new_n372), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n380), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n821), .B1(new_n823), .B2(G68), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n280), .B(new_n375), .C1(new_n824), .C2(new_n377), .ZN(new_n825));
  INV_X1    g0625(.A(new_n408), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n421), .A2(new_n422), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n819), .B(new_n827), .C1(new_n828), .C2(new_n636), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n419), .A2(new_n644), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n411), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(KEYINPUT37), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT109), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n416), .A2(new_n420), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n416), .A2(new_n819), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT37), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n835), .A2(new_n836), .A3(new_n837), .A4(new_n411), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT109), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n832), .A2(new_n839), .A3(KEYINPUT37), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n834), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  AND3_X1   g0641(.A1(new_n829), .A2(KEYINPUT38), .A3(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n836), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n423), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n835), .A2(new_n836), .A3(new_n411), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n838), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT38), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(KEYINPUT112), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n829), .A2(new_n841), .A3(KEYINPUT38), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT112), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n423), .A2(new_n843), .B1(new_n846), .B2(new_n838), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n850), .B(new_n851), .C1(KEYINPUT38), .C2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n818), .A2(new_n849), .A3(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT40), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT38), .B1(new_n829), .B2(new_n841), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n842), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n817), .A2(new_n694), .A3(new_n696), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n463), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n861), .A2(new_n697), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n860), .B(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(G330), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT113), .Z(new_n865));
  OAI21_X1  g0665(.A(new_n638), .B1(new_n682), .B2(new_n861), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT111), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n828), .A2(new_n644), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n355), .A2(new_n646), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n869), .A2(KEYINPUT108), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(KEYINPUT108), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n807), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n814), .A2(new_n816), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n874), .A2(new_n857), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT110), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT39), .B1(new_n842), .B2(new_n856), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT39), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n850), .B(new_n879), .C1(KEYINPUT38), .C2(new_n852), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n877), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n829), .A2(new_n841), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n850), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT110), .B1(new_n885), .B2(KEYINPUT39), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n458), .A2(new_n646), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n868), .B(new_n876), .C1(new_n887), .C2(new_n889), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n867), .B(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n865), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n865), .A2(new_n891), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n892), .B1(new_n894), .B2(KEYINPUT114), .ZN(new_n895));
  OAI221_X1 g0695(.A(new_n895), .B1(KEYINPUT114), .B2(new_n894), .C1(new_n218), .C2(new_n640), .ZN(new_n896));
  OAI211_X1 g0696(.A(G116), .B(new_n226), .C1(new_n583), .C2(KEYINPUT35), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n897), .B(KEYINPUT107), .Z(new_n898));
  NAND2_X1  g0698(.A1(new_n583), .A2(KEYINPUT35), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT36), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n224), .A2(new_n361), .A3(G77), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(G50), .B2(new_n374), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(G1), .A3(new_n228), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n896), .A2(new_n901), .A3(new_n904), .ZN(G367));
  NOR2_X1   g0705(.A1(new_n733), .A2(new_n209), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT46), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n724), .B2(new_n734), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(G283), .B2(new_n714), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n731), .A2(G311), .ZN(new_n910));
  INV_X1    g0710(.A(new_n790), .ZN(new_n911));
  INV_X1    g0711(.A(G317), .ZN(new_n912));
  OAI221_X1 g0712(.A(new_n379), .B1(new_n719), .B2(new_n912), .C1(new_n204), .C2(new_n727), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n911), .A2(G294), .B1(new_n914), .B2(KEYINPUT119), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n739), .A2(new_n205), .B1(new_n906), .B2(KEYINPUT46), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT119), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n916), .B1(new_n917), .B2(new_n913), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n909), .A2(new_n910), .A3(new_n915), .A4(new_n918), .ZN(new_n919));
  OAI221_X1 g0719(.A(new_n292), .B1(new_n771), .B2(new_n733), .C1(new_n724), .C2(new_n264), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(G50), .B2(new_n714), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n727), .A2(new_n446), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(G143), .B2(new_n731), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n739), .A2(new_n374), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n911), .B2(G159), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n921), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n719), .A2(new_n776), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n919), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT47), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n703), .B1(new_n929), .B2(new_n756), .ZN(new_n930));
  INV_X1    g0730(.A(new_n761), .ZN(new_n931));
  OAI221_X1 g0731(.A(new_n760), .B1(new_n230), .B2(new_n346), .C1(new_n241), .C2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n572), .A2(new_n647), .ZN(new_n933));
  MUX2_X1   g0733(.A(new_n573), .B(new_n623), .S(new_n933), .Z(new_n934));
  OAI211_X1 g0734(.A(new_n930), .B(new_n932), .C1(new_n768), .C2(new_n934), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n606), .B(new_n609), .C1(new_n608), .C2(new_n647), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n600), .A2(new_n605), .A3(new_n646), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n657), .A2(new_n661), .A3(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT42), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n936), .A2(new_n532), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n941), .A2(new_n606), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n939), .A2(new_n940), .B1(new_n646), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT115), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n939), .A2(new_n940), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n943), .A2(new_n944), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n945), .A2(new_n950), .A3(new_n946), .A4(new_n947), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n953), .A2(KEYINPUT116), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(KEYINPUT116), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n938), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n660), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n956), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n702), .A2(G1), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n657), .B(new_n661), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n705), .B2(new_n706), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT117), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n704), .A2(new_n962), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT118), .Z(new_n966));
  NAND2_X1  g0766(.A1(new_n963), .A2(KEYINPUT117), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n662), .A2(KEYINPUT44), .A3(new_n938), .ZN(new_n969));
  OAI21_X1  g0769(.A(KEYINPUT44), .B1(new_n662), .B2(new_n938), .ZN(new_n970));
  AND3_X1   g0770(.A1(new_n662), .A2(KEYINPUT45), .A3(new_n938), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT45), .B1(new_n662), .B2(new_n938), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n969), .B(new_n970), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n659), .B(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n700), .B1(new_n968), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n664), .B(KEYINPUT41), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n961), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n935), .B1(new_n960), .B2(new_n977), .ZN(G387));
  INV_X1    g0778(.A(new_n700), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n968), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n964), .A2(new_n966), .A3(new_n967), .A4(new_n700), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n980), .A2(new_n664), .A3(new_n981), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G303), .A2(new_n714), .B1(new_n723), .B2(G317), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n983), .B1(new_n725), .B2(new_n753), .C1(new_n716), .C2(new_n790), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT48), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n787), .B2(new_n739), .C1(new_n522), .C2(new_n733), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT49), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n720), .A2(G326), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n292), .B1(new_n728), .B2(G116), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n273), .A2(new_n740), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n715), .A2(new_n374), .B1(new_n204), .B2(new_n727), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n379), .B(new_n992), .C1(G150), .C2(new_n720), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n733), .A2(new_n446), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n739), .A2(new_n346), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(G159), .C2(new_n731), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n993), .B(new_n996), .C1(new_n214), .C2(new_n724), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n990), .B1(new_n991), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT120), .Z(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n756), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n657), .A2(new_n768), .ZN(new_n1001));
  OR3_X1    g0801(.A1(new_n344), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1002));
  OAI21_X1  g0802(.A(KEYINPUT50), .B1(new_n344), .B2(G50), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n1002), .A2(new_n1003), .A3(new_n762), .A4(new_n666), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(G68), .B2(G77), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n761), .B1(new_n238), .B2(new_n762), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n230), .B(new_n292), .C1(G116), .C2(new_n545), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n230), .A2(G107), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n760), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1000), .A2(new_n708), .A3(new_n1001), .A4(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n961), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n982), .B(new_n1011), .C1(new_n1012), .C2(new_n968), .ZN(G393));
  OAI221_X1 g0813(.A(new_n760), .B1(new_n204), .B2(new_n230), .C1(new_n249), .C2(new_n931), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n723), .A2(G311), .B1(G317), .B2(new_n731), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT52), .Z(new_n1016));
  AOI21_X1  g0816(.A(new_n292), .B1(new_n720), .B2(G322), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(new_n522), .C2(new_n715), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n733), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G283), .A2(new_n1019), .B1(new_n738), .B2(G116), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n205), .B2(new_n727), .C1(new_n790), .C2(new_n734), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n723), .A2(G159), .B1(G150), .B2(new_n731), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT51), .Z(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n786), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n733), .A2(new_n374), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n739), .A2(new_n446), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(G143), .C2(new_n720), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n911), .A2(G50), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n715), .A2(new_n344), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1027), .A2(new_n292), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n1018), .A2(new_n1021), .B1(new_n1024), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n703), .B1(new_n1031), .B2(new_n756), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1014), .B(new_n1032), .C1(new_n938), .C2(new_n768), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n974), .B2(new_n1012), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n981), .A2(new_n974), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n665), .B1(new_n981), .B2(new_n974), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(G390));
  INV_X1    g0838(.A(KEYINPUT121), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n888), .B1(new_n872), .B2(new_n873), .ZN(new_n1040));
  NOR3_X1   g0840(.A1(new_n881), .A2(new_n886), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n869), .B1(new_n680), .B2(new_n806), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n873), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n889), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n849), .A2(new_n853), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n698), .A2(G330), .A3(new_n817), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1041), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n880), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n879), .B1(new_n884), .B2(new_n850), .ZN(new_n1051));
  OAI21_X1  g0851(.A(KEYINPUT110), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n878), .A2(new_n877), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n874), .A2(new_n889), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n646), .B(new_n805), .C1(new_n674), .C2(new_n679), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n873), .B1(new_n1056), .B2(new_n869), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1057), .A2(new_n849), .A3(new_n853), .A4(new_n889), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1047), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1039), .B1(new_n1049), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n463), .A2(G330), .A3(new_n698), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1061), .B(new_n638), .C1(new_n682), .C2(new_n861), .ZN(new_n1062));
  AND3_X1   g0862(.A1(new_n698), .A2(G330), .A3(new_n808), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1047), .B(new_n1042), .C1(new_n1063), .C2(new_n873), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n694), .A2(G330), .A3(new_n696), .A4(new_n803), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n1043), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1047), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n872), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1062), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1048), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1055), .A2(new_n1047), .A3(new_n1058), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1071), .A2(new_n1072), .A3(KEYINPUT121), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1060), .A2(new_n1070), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT122), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1071), .A2(new_n1069), .A3(new_n1072), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1060), .A2(KEYINPUT122), .A3(new_n1070), .A4(new_n1073), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1076), .A2(new_n664), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n1049), .A2(new_n1059), .A3(new_n1012), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1026), .B1(new_n911), .B2(G107), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n714), .A2(G97), .B1(G87), .B2(new_n1019), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n379), .B1(new_n719), .B2(new_n522), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n723), .B2(G116), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n731), .A2(G283), .B1(new_n728), .B2(G68), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1081), .A2(new_n1082), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  XOR2_X1   g0886(.A(KEYINPUT54), .B(G143), .Z(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n781), .A2(new_n724), .B1(new_n715), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(G128), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n753), .A2(new_n1090), .B1(new_n739), .B2(new_n777), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n292), .B1(new_n727), .B2(new_n214), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n1089), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(G125), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1093), .B1(new_n1094), .B2(new_n719), .C1(new_n776), .C2(new_n790), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1019), .A2(G150), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT53), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1086), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n756), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n795), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1099), .B1(new_n272), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n887), .B2(new_n757), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1080), .B1(new_n708), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1079), .A2(new_n1103), .ZN(G378));
  NAND2_X1  g0904(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n875), .B1(new_n1105), .B2(new_n888), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n318), .B1(new_n313), .B2(new_n317), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n320), .A2(KEYINPUT75), .A3(new_n321), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1107), .A2(new_n1108), .B1(KEYINPUT10), .B2(new_n310), .ZN(new_n1109));
  OAI21_X1  g0909(.A(KEYINPUT55), .B1(new_n1109), .B2(new_n633), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT55), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n323), .A2(new_n1111), .A3(new_n329), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n326), .A2(new_n819), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT56), .Z(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1110), .A2(new_n1112), .A3(new_n1115), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1119), .A2(G330), .A3(new_n859), .A4(new_n854), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n854), .A2(new_n859), .A3(G330), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1119), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1106), .A2(new_n868), .A3(new_n1120), .A4(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1120), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n890), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1012), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1122), .A2(new_n757), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G132), .A2(new_n774), .B1(new_n738), .B2(G150), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n1094), .B2(new_n753), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT123), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n1088), .B2(new_n733), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1019), .A2(KEYINPUT123), .A3(new_n1087), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1132), .B(new_n1133), .C1(new_n715), .C2(new_n776), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1130), .B(new_n1134), .C1(G128), .C2(new_n723), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT59), .ZN(new_n1136));
  AOI21_X1  g0936(.A(G41), .B1(new_n728), .B2(G159), .ZN(new_n1137));
  AOI21_X1  g0937(.A(G33), .B1(new_n720), .B2(G124), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n214), .B1(new_n367), .B2(G41), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n723), .A2(G107), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n714), .A2(new_n345), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n292), .B1(new_n720), .B2(G283), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1141), .A2(new_n1142), .A3(new_n297), .A4(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n994), .B1(new_n270), .B2(new_n728), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n204), .B2(new_n740), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n753), .A2(new_n209), .ZN(new_n1147));
  NOR4_X1   g0947(.A1(new_n1144), .A2(new_n1146), .A3(new_n924), .A4(new_n1147), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT58), .Z(new_n1149));
  NAND3_X1  g0949(.A1(new_n1139), .A2(new_n1140), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n703), .B1(new_n1150), .B2(new_n756), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1128), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n214), .B2(new_n795), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1127), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1062), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1077), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT57), .ZN(new_n1160));
  AOI21_X1  g0960(.A(KEYINPUT124), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT124), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1162), .B(KEYINPUT57), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1156), .A2(new_n1077), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n665), .B1(new_n1165), .B2(KEYINPUT57), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1155), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(G375));
  OAI221_X1 g0968(.A(new_n379), .B1(new_n734), .B2(new_n719), .C1(new_n724), .C2(new_n787), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n922), .B(new_n1169), .C1(G107), .C2(new_n714), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n733), .A2(new_n204), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n995), .B(new_n1171), .C1(new_n911), .C2(G116), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(new_n522), .C2(new_n753), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n739), .A2(new_n214), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n753), .A2(new_n781), .B1(new_n777), .B2(new_n733), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n911), .B2(new_n1087), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n714), .A2(G150), .B1(new_n270), .B2(new_n728), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n292), .B1(new_n719), .B2(new_n1090), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n723), .B2(G137), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1173), .B1(new_n1174), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n756), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(G68), .B2(new_n1100), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n703), .B(new_n1183), .C1(new_n1043), .C2(new_n757), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1184), .B1(new_n1185), .B2(new_n961), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n976), .B1(new_n1185), .B2(new_n1156), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1186), .B1(new_n1187), .B2(new_n1069), .ZN(G381));
  NOR2_X1   g0988(.A1(G375), .A2(G378), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1190), .A2(G384), .A3(G381), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n935), .B(new_n1037), .C1(new_n960), .C2(new_n977), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1192), .A2(G396), .A3(G393), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1191), .A2(new_n1193), .ZN(G407));
  OAI211_X1 g0994(.A(G407), .B(G213), .C1(G343), .C2(new_n1190), .ZN(G409));
  XNOR2_X1  g0995(.A(G393), .B(G396), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(G387), .A2(G390), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n1192), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1196), .A2(new_n1192), .A3(new_n1198), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT62), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n976), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1154), .B1(new_n1159), .B2(new_n1204), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1079), .A2(new_n1103), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n1167), .B2(G378), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n645), .A2(G213), .ZN(new_n1208));
  OAI21_X1  g1008(.A(KEYINPUT125), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1162), .B1(new_n1165), .B2(KEYINPUT57), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1159), .A2(KEYINPUT124), .A3(new_n1160), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1210), .A2(new_n1166), .A3(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(G378), .A2(new_n1154), .A3(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1079), .A2(new_n1103), .A3(new_n1205), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1208), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT125), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1209), .A2(new_n1217), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1219), .A2(KEYINPUT60), .A3(new_n1062), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1220), .A2(new_n664), .A3(new_n1070), .ZN(new_n1221));
  AOI21_X1  g1021(.A(KEYINPUT60), .B1(new_n1219), .B2(new_n1062), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1186), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(G384), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1203), .B1(new_n1218), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1208), .A2(G2897), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1224), .B(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1209), .A2(new_n1217), .A3(new_n1228), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1223), .B(G384), .Z(new_n1230));
  AOI211_X1 g1030(.A(new_n1208), .B(new_n1230), .C1(new_n1213), .C2(new_n1214), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT61), .B1(new_n1231), .B2(new_n1203), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1202), .B1(new_n1225), .B2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1218), .A2(KEYINPUT63), .A3(new_n1224), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT61), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1231), .ZN(new_n1237));
  OAI21_X1  g1037(.A(KEYINPUT63), .B1(new_n1215), .B2(new_n1227), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1202), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1235), .A2(new_n1236), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1234), .A2(new_n1240), .ZN(G405));
  INV_X1    g1041(.A(new_n1201), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1196), .B1(new_n1198), .B2(new_n1192), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1230), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1200), .A2(new_n1201), .A3(new_n1224), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT126), .B1(new_n1167), .B2(G378), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n1248), .A2(new_n1249), .B1(G378), .B2(new_n1167), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1167), .A2(G378), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1250), .A2(new_n1254), .ZN(G402));
endmodule


