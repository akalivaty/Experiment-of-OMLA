//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n552,
    new_n554, new_n555, new_n556, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1231, new_n1232,
    new_n1233;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT64), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT66), .B(G2104), .ZN(new_n461));
  OAI211_X1 g036(.A(G137), .B(new_n460), .C1(new_n461), .C2(new_n459), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(G101), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  XNOR2_X1  g041(.A(new_n466), .B(KEYINPUT65), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n460), .A2(new_n469), .A3(G125), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n465), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n464), .A2(new_n471), .ZN(G160));
  OAI21_X1  g047(.A(new_n460), .B1(new_n461), .B2(new_n459), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(new_n465), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n477));
  INV_X1    g052(.A(G136), .ZN(new_n478));
  INV_X1    g053(.A(new_n460), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n468), .A2(KEYINPUT66), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n479), .B1(new_n483), .B2(KEYINPUT3), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(new_n465), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n475), .B(new_n477), .C1(new_n478), .C2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NOR2_X1   g062(.A1(new_n481), .A2(G2104), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n468), .A2(KEYINPUT66), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT3), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g065(.A1(KEYINPUT4), .A2(G138), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n490), .A2(new_n465), .A3(new_n460), .A4(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n460), .A2(new_n469), .A3(G138), .A4(new_n465), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n468), .A2(G2105), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n493), .A2(new_n494), .B1(G102), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(G114), .A2(G2104), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n484), .B2(G126), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n492), .B(new_n496), .C1(new_n499), .C2(new_n465), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  XNOR2_X1  g076(.A(KEYINPUT67), .B(G651), .ZN(new_n502));
  INV_X1    g077(.A(G62), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(KEYINPUT68), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT5), .A3(G543), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n503), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(G75), .A2(G543), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n502), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n514), .A2(KEYINPUT67), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT6), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n506), .A2(new_n508), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  XOR2_X1   g094(.A(KEYINPUT69), .B(G88), .Z(new_n520));
  NAND4_X1  g095(.A1(new_n516), .A2(new_n517), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT6), .ZN(new_n523));
  OAI211_X1 g098(.A(G543), .B(new_n519), .C1(new_n502), .C2(new_n523), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n511), .B(new_n521), .C1(new_n522), .C2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  AND3_X1   g101(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G89), .ZN(new_n528));
  INV_X1    g103(.A(new_n524), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G51), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n528), .A2(new_n530), .A3(new_n531), .A4(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  AOI22_X1  g110(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  XOR2_X1   g111(.A(KEYINPUT67), .B(G651), .Z(new_n537));
  OR2_X1    g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n527), .A2(G90), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n529), .A2(G52), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  AOI22_X1  g117(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n537), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n527), .A2(G81), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n529), .A2(G43), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(KEYINPUT70), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(KEYINPUT70), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  XOR2_X1   g128(.A(KEYINPUT71), .B(KEYINPUT8), .Z(new_n554));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(G188));
  INV_X1    g132(.A(KEYINPUT72), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n517), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n506), .A2(KEYINPUT72), .A3(new_n508), .ZN(new_n560));
  XOR2_X1   g135(.A(KEYINPUT73), .B(G65), .Z(new_n561));
  NAND3_X1  g136(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G651), .ZN(new_n565));
  AND4_X1   g140(.A1(G91), .A2(new_n516), .A3(new_n517), .A4(new_n519), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n518), .B1(new_n537), .B2(KEYINPUT6), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n568), .A2(new_n569), .A3(G53), .A4(G543), .ZN(new_n570));
  INV_X1    g145(.A(G53), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT9), .B1(new_n524), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n565), .A2(new_n567), .A3(new_n573), .ZN(G299));
  NAND4_X1  g149(.A1(new_n516), .A2(G49), .A3(G543), .A4(new_n519), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n516), .A2(G87), .A3(new_n517), .A4(new_n519), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT74), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT74), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n575), .A2(new_n576), .A3(new_n580), .A4(new_n577), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(G288));
  NAND4_X1  g157(.A1(new_n516), .A2(G86), .A3(new_n517), .A4(new_n519), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n506), .B2(new_n508), .ZN(new_n585));
  AND2_X1   g160(.A1(G73), .A2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n502), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n516), .A2(G48), .A3(G543), .A4(new_n519), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n583), .A2(new_n587), .A3(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(new_n537), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n527), .A2(G85), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n529), .A2(G47), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(G290));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NOR2_X1   g170(.A1(G171), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n527), .A2(G92), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT76), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(KEYINPUT10), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n598), .B(KEYINPUT76), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n559), .A2(G66), .A3(new_n560), .ZN(new_n605));
  INV_X1    g180(.A(G79), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(new_n504), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G651), .B1(G54), .B2(new_n529), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n601), .A2(new_n604), .A3(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n597), .B1(new_n610), .B2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(KEYINPUT75), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(KEYINPUT75), .B2(new_n596), .ZN(G284));
  OAI21_X1  g188(.A(new_n612), .B1(KEYINPUT75), .B2(new_n596), .ZN(G321));
  NAND2_X1  g189(.A1(G299), .A2(new_n595), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n595), .B2(G168), .ZN(G297));
  OAI21_X1  g191(.A(new_n615), .B1(new_n595), .B2(G168), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n610), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND3_X1  g194(.A1(new_n548), .A2(new_n595), .A3(new_n549), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n609), .A2(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n595), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND4_X1  g198(.A1(new_n461), .A2(new_n465), .A3(new_n460), .A4(new_n469), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  INV_X1    g201(.A(G2100), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n474), .A2(G123), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n473), .A2(G2105), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G135), .ZN(new_n631));
  NOR2_X1   g206(.A1(G99), .A2(G2105), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(new_n465), .B2(G111), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n629), .B(new_n631), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G2096), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n628), .A2(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2435), .ZN(new_n639));
  XOR2_X1   g214(.A(G2427), .B(G2438), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT77), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n648), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(G14), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G401));
  XNOR2_X1  g228(.A(G2072), .B(G2078), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT78), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XOR2_X1   g231(.A(G2067), .B(G2678), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT18), .Z(new_n660));
  INV_X1    g235(.A(new_n656), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(new_n657), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n655), .A2(KEYINPUT17), .A3(new_n662), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n664));
  OAI221_X1 g239(.A(new_n663), .B1(new_n661), .B2(new_n657), .C1(new_n664), .C2(new_n655), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(new_n635), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(new_n627), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT79), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT20), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n672), .A2(new_n673), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n679), .A2(new_n671), .A3(new_n674), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n677), .B(new_n680), .C1(new_n671), .C2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n683), .B(new_n684), .Z(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT22), .B(G1981), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G229));
  MUX2_X1   g263(.A(G23), .B(new_n578), .S(G16), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT80), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT33), .B(G1976), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT80), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n689), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n691), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G22), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G166), .B2(new_n697), .ZN(new_n699));
  INV_X1    g274(.A(G1971), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n697), .A2(G6), .ZN(new_n702));
  INV_X1    g277(.A(G305), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n697), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT32), .B(G1981), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n692), .A2(new_n696), .A3(new_n701), .A4(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT34), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT81), .B(KEYINPUT36), .Z(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n474), .A2(G119), .ZN(new_n714));
  OR2_X1    g289(.A1(G95), .A2(G2105), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n715), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n716));
  INV_X1    g291(.A(G131), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n714), .B(new_n716), .C1(new_n717), .C2(new_n485), .ZN(new_n718));
  MUX2_X1   g293(.A(G25), .B(new_n718), .S(G29), .Z(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT35), .B(G1991), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n697), .A2(G24), .ZN(new_n722));
  INV_X1    g297(.A(G290), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(new_n697), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(G1986), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(G1986), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n719), .A2(new_n720), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n721), .A2(new_n725), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n711), .A2(KEYINPUT82), .A3(new_n713), .A4(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT82), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n711), .A2(new_n729), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(KEYINPUT36), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n712), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n730), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n697), .A2(G4), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n610), .B2(new_n697), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT83), .B(G1348), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G16), .A2(G19), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n550), .B2(G16), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G1341), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G29), .A2(G32), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n484), .A2(G141), .B1(G105), .B2(new_n461), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(G2105), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n474), .A2(G129), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT26), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n746), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n744), .B1(new_n752), .B2(G29), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT27), .B(G1996), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(G162), .A2(G29), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G29), .B2(G35), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT29), .B(G2090), .Z(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  INV_X1    g335(.A(G29), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G27), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G164), .B2(new_n761), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G2078), .ZN(new_n764));
  AND4_X1   g339(.A1(new_n755), .A2(new_n759), .A3(new_n760), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(G171), .A2(G16), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G5), .B2(G16), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G1966), .ZN(new_n769));
  NAND2_X1  g344(.A1(G168), .A2(G16), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G16), .B2(G21), .ZN(new_n771));
  OAI221_X1 g346(.A(new_n765), .B1(G1961), .B2(new_n768), .C1(new_n769), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(G299), .A2(G16), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n697), .A2(KEYINPUT23), .A3(G20), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT23), .ZN(new_n775));
  INV_X1    g350(.A(G20), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(G16), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n773), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1956), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT30), .B(G28), .ZN(new_n780));
  OR2_X1    g355(.A1(KEYINPUT31), .A2(G11), .ZN(new_n781));
  NAND2_X1  g356(.A1(KEYINPUT31), .A2(G11), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n780), .A2(new_n761), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n634), .B2(new_n761), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT84), .Z(new_n785));
  OR2_X1    g360(.A1(new_n779), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n772), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n753), .A2(new_n754), .ZN(new_n788));
  INV_X1    g363(.A(G2078), .ZN(new_n789));
  INV_X1    g364(.A(new_n763), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G2072), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n761), .A2(G33), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n460), .A2(new_n469), .A3(G127), .ZN(new_n794));
  INV_X1    g369(.A(G115), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n468), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n630), .A2(G139), .B1(G2105), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n495), .A2(G103), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT25), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n793), .B1(new_n800), .B2(G29), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n771), .A2(new_n769), .B1(new_n792), .B2(new_n801), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n791), .B(new_n802), .C1(new_n792), .C2(new_n801), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G1961), .B2(new_n768), .ZN(new_n804));
  OR2_X1    g379(.A1(KEYINPUT24), .A2(G34), .ZN(new_n805));
  NAND2_X1  g380(.A1(KEYINPUT24), .A2(G34), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n805), .A2(new_n761), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G160), .B2(new_n761), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(G2084), .Z(new_n809));
  AND3_X1   g384(.A1(new_n787), .A2(new_n804), .A3(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n735), .A2(new_n739), .A3(new_n743), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n761), .A2(G26), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n474), .A2(G128), .ZN(new_n813));
  OR2_X1    g388(.A1(G104), .A2(G2105), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n814), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n815));
  INV_X1    g390(.A(G140), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n813), .B(new_n815), .C1(new_n816), .C2(new_n485), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n812), .B1(new_n818), .B2(new_n761), .ZN(new_n819));
  MUX2_X1   g394(.A(new_n812), .B(new_n819), .S(KEYINPUT28), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G2067), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n811), .A2(new_n821), .ZN(G311));
  AND3_X1   g397(.A1(new_n735), .A2(new_n743), .A3(new_n810), .ZN(new_n823));
  INV_X1    g398(.A(new_n821), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n823), .A2(KEYINPUT85), .A3(new_n824), .A4(new_n739), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT85), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n811), .B2(new_n821), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(G150));
  AND2_X1   g403(.A1(new_n517), .A2(G67), .ZN(new_n829));
  AND2_X1   g404(.A1(G80), .A2(G543), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n502), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT86), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g408(.A(KEYINPUT86), .B(new_n502), .C1(new_n829), .C2(new_n830), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT87), .ZN(new_n836));
  AOI22_X1  g411(.A1(G93), .A2(new_n527), .B1(new_n529), .B2(G55), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n837), .A2(new_n833), .A3(new_n834), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(KEYINPUT87), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(KEYINPUT88), .B(G860), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT37), .Z(new_n845));
  NOR2_X1   g420(.A1(new_n609), .A2(new_n618), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n841), .A2(new_n547), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n548), .A2(new_n549), .B1(new_n837), .B2(new_n835), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n848), .B(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n845), .B1(new_n853), .B2(new_n843), .ZN(G145));
  XNOR2_X1  g429(.A(new_n486), .B(KEYINPUT89), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(G160), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n634), .ZN(new_n857));
  INV_X1    g432(.A(new_n625), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(new_n465), .B2(G118), .ZN(new_n859));
  INV_X1    g434(.A(G106), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n859), .B1(new_n860), .B2(new_n465), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n861), .B1(new_n474), .B2(G130), .ZN(new_n862));
  INV_X1    g437(.A(G142), .ZN(new_n863));
  OAI21_X1  g438(.A(KEYINPUT91), .B1(new_n485), .B2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT91), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n630), .A2(new_n865), .A3(G142), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n862), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(new_n718), .Z(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT92), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n868), .A2(KEYINPUT92), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n858), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n817), .B(new_n500), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT90), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n800), .A2(new_n874), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n873), .A2(new_n875), .ZN(new_n877));
  OR3_X1    g452(.A1(new_n876), .A2(new_n877), .A3(new_n751), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n868), .A2(KEYINPUT92), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n879), .A2(new_n625), .A3(new_n869), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n751), .B1(new_n876), .B2(new_n877), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n872), .A2(new_n878), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT95), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n857), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n878), .A2(new_n881), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n886), .A2(KEYINPUT95), .A3(new_n880), .A4(new_n872), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT93), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n870), .A2(new_n871), .A3(new_n858), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n625), .B1(new_n879), .B2(new_n869), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n872), .A2(new_n880), .A3(KEYINPUT93), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(new_n892), .A3(new_n885), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n884), .A2(new_n887), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT96), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n884), .A2(new_n887), .A3(new_n893), .A4(KEYINPUT96), .ZN(new_n897));
  AOI21_X1  g472(.A(G37), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n891), .A2(new_n892), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n886), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(KEYINPUT94), .A3(new_n893), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n901), .B(new_n857), .C1(KEYINPUT94), .C2(new_n893), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g479(.A(new_n852), .B(new_n621), .Z(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n609), .A2(G299), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n609), .A2(G299), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n609), .A2(G299), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(KEYINPUT41), .A3(new_n907), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n905), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n907), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n913), .B1(new_n914), .B2(new_n905), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n915), .A2(KEYINPUT42), .ZN(new_n916));
  XNOR2_X1  g491(.A(G305), .B(new_n578), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(new_n723), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(G166), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n915), .A2(KEYINPUT42), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n919), .B1(new_n916), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g497(.A(G868), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n842), .A2(new_n595), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(G295));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n924), .ZN(G331));
  INV_X1    g501(.A(G37), .ZN(new_n927));
  NAND2_X1  g502(.A1(G168), .A2(KEYINPUT97), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT97), .ZN(new_n929));
  NAND2_X1  g504(.A1(G286), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(G171), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(G286), .A2(G301), .A3(new_n929), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n849), .A2(new_n851), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n547), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n935), .B1(new_n838), .B2(new_n840), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n932), .B(new_n931), .C1(new_n936), .C2(new_n850), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT98), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n934), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n849), .A2(new_n851), .A3(new_n933), .A4(KEYINPUT98), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n939), .A2(new_n910), .A3(new_n912), .A4(new_n940), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n934), .A2(new_n937), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(new_n907), .A3(new_n911), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g519(.A(KEYINPUT99), .B(new_n927), .C1(new_n944), .C2(new_n919), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n941), .A2(new_n943), .A3(new_n919), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT100), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT100), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n941), .A2(new_n943), .A3(new_n948), .A4(new_n919), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT99), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n919), .B1(new_n941), .B2(new_n943), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(new_n952), .B2(G37), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n945), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n910), .A2(new_n912), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n957), .A2(new_n942), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n914), .B1(new_n939), .B2(new_n940), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n960), .A2(new_n919), .ZN(new_n961));
  AND4_X1   g536(.A1(KEYINPUT43), .A2(new_n961), .A3(new_n950), .A4(new_n927), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT44), .B1(new_n956), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n961), .A2(new_n950), .A3(new_n955), .A4(new_n927), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n963), .A2(new_n968), .ZN(G397));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n492), .A2(new_n496), .ZN(new_n971));
  OAI211_X1 g546(.A(G126), .B(new_n460), .C1(new_n461), .C2(new_n459), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n465), .B1(new_n972), .B2(new_n497), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n970), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n467), .A2(new_n470), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(G2105), .ZN(new_n978));
  INV_X1    g553(.A(G101), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n483), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(new_n484), .B2(G137), .ZN(new_n981));
  OAI211_X1 g556(.A(G40), .B(new_n978), .C1(new_n981), .C2(G2105), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n976), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G2067), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n817), .B(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1996), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n752), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n751), .A2(G1996), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n987), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n718), .A2(new_n720), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n818), .A2(new_n985), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n984), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n983), .B1(new_n987), .B2(new_n751), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n983), .A2(KEYINPUT46), .A3(new_n988), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT46), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n984), .B2(G1996), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n996), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  XOR2_X1   g575(.A(new_n1000), .B(KEYINPUT47), .Z(new_n1001));
  INV_X1    g576(.A(new_n992), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n991), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1003), .B1(new_n720), .B2(new_n718), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1004), .A2(new_n984), .ZN(new_n1005));
  NOR2_X1   g580(.A1(G290), .A2(G1986), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n983), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1007), .B(KEYINPUT48), .ZN(new_n1008));
  AOI211_X1 g583(.A(new_n995), .B(new_n1001), .C1(new_n1005), .C2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G8), .ZN(new_n1010));
  INV_X1    g585(.A(new_n974), .ZN(new_n1011));
  INV_X1    g586(.A(G40), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n464), .A2(new_n1012), .A3(new_n471), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1010), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1981), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n583), .A2(new_n587), .A3(new_n588), .A4(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT104), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT49), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(G305), .B2(G1981), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(G305), .A2(new_n1020), .A3(G1981), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1019), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AND3_X1   g599(.A1(G305), .A2(new_n1020), .A3(G1981), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n1025), .A2(new_n1021), .A3(new_n1018), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1014), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1976), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT52), .B1(G288), .B2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n575), .A2(new_n576), .A3(G1976), .A4(new_n577), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT103), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n1030), .A2(KEYINPUT103), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1029), .A2(new_n1014), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1013), .A2(new_n500), .A3(new_n970), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1034), .A2(G8), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT52), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1027), .A2(new_n1033), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT109), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1022), .A2(new_n1019), .A3(new_n1023), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1018), .B1(new_n1025), .B2(new_n1021), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1042), .A2(new_n1014), .B1(KEYINPUT52), .B2(new_n1035), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(KEYINPUT109), .A3(new_n1033), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(new_n500), .B2(new_n970), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1046), .A2(new_n982), .ZN(new_n1047));
  INV_X1    g622(.A(G2090), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1011), .A2(new_n1045), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT45), .B(new_n970), .C1(new_n971), .C2(new_n973), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n976), .A2(new_n1013), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n700), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1010), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT102), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G303), .A2(G8), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT101), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT55), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1057), .A2(KEYINPUT55), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1056), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1055), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1061), .B(KEYINPUT102), .C1(new_n1056), .C2(new_n1060), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1039), .A2(new_n1044), .B1(new_n1054), .B2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT110), .B(G2084), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1047), .A2(new_n1049), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1052), .A2(new_n769), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1071), .A2(new_n1010), .A3(G286), .ZN(new_n1072));
  AOI211_X1 g647(.A(KEYINPUT107), .B(new_n982), .C1(KEYINPUT50), .C2(new_n974), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT107), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n974), .A2(KEYINPUT50), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1074), .B1(new_n1075), .B2(new_n1013), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1049), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT108), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT108), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1079), .B(new_n1049), .C1(new_n1073), .C2(new_n1076), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1078), .A2(new_n1048), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1010), .B1(new_n1081), .B2(new_n1053), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1067), .B(new_n1072), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT63), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1037), .A2(KEYINPUT105), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT105), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1043), .A2(new_n1088), .A3(new_n1033), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n1054), .B2(new_n1066), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1054), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1083), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1085), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(new_n1072), .A3(new_n1094), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1042), .A2(G1976), .A3(G288), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1016), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1014), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1054), .A2(new_n1066), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1098), .B1(new_n1090), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT106), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT106), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1098), .B(new_n1102), .C1(new_n1090), .C2(new_n1099), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1086), .A2(new_n1095), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1069), .A2(G168), .A3(new_n1070), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1105), .B1(new_n1106), .B2(G8), .ZN(new_n1107));
  OAI21_X1  g682(.A(KEYINPUT51), .B1(new_n1071), .B2(G168), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1106), .A2(G8), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n1111));
  OR2_X1    g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n976), .A2(new_n789), .A3(new_n1013), .A4(new_n1051), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1113), .A2(KEYINPUT119), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1115), .B1(new_n1113), .B2(KEYINPUT119), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1119));
  INV_X1    g694(.A(G1961), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT120), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1113), .A2(new_n1124), .A3(new_n1115), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1121), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(G171), .B1(new_n1118), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1127), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1049), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT107), .B1(new_n1046), .B2(new_n982), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1075), .A2(new_n1074), .A3(new_n1013), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(G2090), .B1(new_n1133), .B2(new_n1079), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1134), .A2(new_n1078), .B1(new_n700), .B2(new_n1052), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1093), .B1(new_n1135), .B2(new_n1010), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1129), .B1(new_n1136), .B2(new_n1067), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1080), .A2(new_n1048), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1079), .B1(new_n1139), .B2(new_n1049), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1053), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1083), .B1(new_n1141), .B2(G8), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT109), .B1(new_n1043), .B2(new_n1033), .ZN(new_n1143));
  AND4_X1   g718(.A1(KEYINPUT109), .A2(new_n1027), .A3(new_n1033), .A4(new_n1036), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1099), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1142), .A2(new_n1145), .A3(KEYINPUT122), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1112), .B(new_n1128), .C1(new_n1137), .C2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1052), .ZN(new_n1148));
  XNOR2_X1  g723(.A(KEYINPUT56), .B(G2072), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1150), .B1(new_n1133), .B2(G1956), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT57), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n566), .B1(new_n564), .B2(G651), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT111), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1153), .A2(new_n1154), .A3(new_n573), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1154), .B1(new_n1153), .B2(new_n573), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1152), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(G299), .A2(KEYINPUT111), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1153), .A2(new_n1154), .A3(new_n573), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1158), .A2(KEYINPUT57), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1151), .A2(new_n1161), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1155), .A2(new_n1156), .A3(new_n1152), .ZN(new_n1163));
  AOI21_X1  g738(.A(KEYINPUT57), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1165), .B(new_n1150), .C1(G1956), .C2(new_n1133), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT118), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1162), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT61), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1151), .A2(KEYINPUT118), .A3(new_n1161), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1166), .A2(KEYINPUT61), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1034), .A2(G2067), .ZN(new_n1173));
  INV_X1    g748(.A(G1348), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1173), .B1(new_n1119), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1175), .A2(KEYINPUT60), .A3(new_n609), .ZN(new_n1176));
  XOR2_X1   g751(.A(KEYINPUT58), .B(G1341), .Z(new_n1177));
  NAND2_X1  g752(.A1(new_n1034), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT116), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1034), .A2(KEYINPUT116), .A3(new_n1177), .ZN(new_n1181));
  XNOR2_X1  g756(.A(KEYINPUT115), .B(G1996), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1180), .B(new_n1181), .C1(new_n1052), .C2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(new_n550), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT117), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1184), .A2(new_n1185), .A3(KEYINPUT59), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(KEYINPUT59), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1183), .A2(new_n550), .A3(new_n1187), .ZN(new_n1188));
  OR2_X1    g763(.A1(new_n1175), .A2(KEYINPUT60), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n609), .B1(new_n1175), .B2(KEYINPUT60), .ZN(new_n1190));
  AOI22_X1  g765(.A1(new_n1186), .A2(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1171), .A2(new_n1172), .A3(new_n1176), .A4(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1161), .B(KEYINPUT114), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT113), .ZN(new_n1194));
  OAI211_X1 g769(.A(new_n1194), .B(new_n1150), .C1(new_n1133), .C2(G1956), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1151), .A2(KEYINPUT113), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1193), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT112), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1198), .B1(new_n1175), .B2(new_n609), .ZN(new_n1199));
  OR3_X1    g774(.A1(new_n1175), .A2(new_n1198), .A3(new_n609), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1197), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1166), .ZN(new_n1202));
  AND2_X1   g777(.A1(new_n1192), .A2(new_n1202), .ZN(new_n1203));
  AND2_X1   g778(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1204));
  XNOR2_X1  g779(.A(KEYINPUT121), .B(G2078), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1148), .A2(KEYINPUT53), .A3(new_n1205), .ZN(new_n1206));
  NAND4_X1  g781(.A1(new_n1204), .A2(G301), .A3(new_n1121), .A4(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(KEYINPUT54), .B1(new_n1127), .B2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1208), .A2(new_n1110), .ZN(new_n1209));
  NAND4_X1  g784(.A1(new_n1204), .A2(KEYINPUT124), .A3(new_n1121), .A4(new_n1206), .ZN(new_n1210));
  NAND4_X1  g785(.A1(new_n1121), .A2(new_n1123), .A3(new_n1125), .A4(new_n1206), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT124), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1210), .A2(new_n1213), .A3(G171), .ZN(new_n1214));
  NAND4_X1  g789(.A1(new_n1204), .A2(G301), .A3(new_n1121), .A4(new_n1117), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1215), .A2(KEYINPUT123), .ZN(new_n1216));
  INV_X1    g791(.A(new_n1126), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT123), .ZN(new_n1218));
  NAND4_X1  g793(.A1(new_n1217), .A2(new_n1218), .A3(G301), .A4(new_n1117), .ZN(new_n1219));
  NAND4_X1  g794(.A1(new_n1214), .A2(new_n1216), .A3(KEYINPUT54), .A4(new_n1219), .ZN(new_n1220));
  OAI211_X1 g795(.A(new_n1209), .B(new_n1220), .C1(new_n1137), .C2(new_n1146), .ZN(new_n1221));
  OAI211_X1 g796(.A(new_n1104), .B(new_n1147), .C1(new_n1203), .C2(new_n1221), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT125), .ZN(new_n1223));
  INV_X1    g798(.A(G1986), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1004), .B1(new_n1224), .B2(new_n723), .ZN(new_n1225));
  OAI21_X1  g800(.A(new_n983), .B1(new_n1225), .B2(new_n1006), .ZN(new_n1226));
  AND3_X1   g801(.A1(new_n1222), .A2(new_n1223), .A3(new_n1226), .ZN(new_n1227));
  AOI21_X1  g802(.A(new_n1223), .B1(new_n1222), .B2(new_n1226), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1009), .B1(new_n1227), .B2(new_n1228), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g804(.A1(new_n652), .A2(G319), .A3(new_n668), .ZN(new_n1231));
  XNOR2_X1  g805(.A(new_n1231), .B(KEYINPUT126), .ZN(new_n1232));
  AOI21_X1  g806(.A(new_n1232), .B1(new_n898), .B2(new_n902), .ZN(new_n1233));
  AND3_X1   g807(.A1(new_n1233), .A2(new_n966), .A3(new_n687), .ZN(G308));
  NAND3_X1  g808(.A1(new_n1233), .A2(new_n966), .A3(new_n687), .ZN(G225));
endmodule


