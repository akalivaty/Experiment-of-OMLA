//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1167, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g0007(.A(KEYINPUT65), .B(G50), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR3_X1   g0009(.A1(new_n207), .A2(new_n209), .A3(G77), .ZN(G353));
  OAI21_X1  g0010(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G50), .A2(G226), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G97), .A2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n214), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n213), .B1(new_n218), .B2(KEYINPUT67), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n219), .B1(KEYINPUT67), .B2(new_n218), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G68), .A2(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G116), .ZN(new_n222));
  INV_X1    g0022(.A(G270), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n220), .B(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(KEYINPUT66), .B(G77), .Z(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n212), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT68), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n212), .A2(G13), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT0), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n231), .B(new_n234), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n235));
  NAND2_X1  g0035(.A1(G1), .A2(G13), .ZN(new_n236));
  INV_X1    g0036(.A(G20), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(G50), .ZN(new_n239));
  NOR2_X1   g0039(.A1(new_n206), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g0040(.A(new_n235), .B1(new_n238), .B2(new_n240), .ZN(G361));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  INV_X1    g0042(.A(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G238), .B(G244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G250), .B(G257), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G264), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n223), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G358));
  XNOR2_X1  g0050(.A(G68), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(new_n239), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(G58), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT69), .B(G107), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(G116), .ZN(new_n255));
  XNOR2_X1  g0055(.A(G87), .B(G97), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n253), .B(new_n257), .ZN(G351));
  AOI21_X1  g0058(.A(new_n236), .B1(G33), .B2(G41), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G226), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT3), .B(G33), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G222), .ZN(new_n267));
  INV_X1    g0067(.A(G223), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n265), .B(new_n267), .C1(new_n268), .C2(new_n266), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n269), .B(new_n259), .C1(new_n225), .C2(new_n265), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n262), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n264), .A2(new_n270), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G190), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(G20), .B1(new_n207), .B2(new_n209), .ZN(new_n277));
  XOR2_X1   g0077(.A(KEYINPUT8), .B(G58), .Z(new_n278));
  INV_X1    g0078(.A(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G20), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n278), .A2(new_n280), .B1(G150), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n236), .ZN(new_n285));
  INV_X1    g0085(.A(G13), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(G1), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n283), .A2(new_n285), .B1(new_n239), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n285), .B1(new_n261), .B2(G20), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n290), .B1(new_n239), .B2(new_n292), .ZN(new_n293));
  XOR2_X1   g0093(.A(new_n293), .B(KEYINPUT70), .Z(new_n294));
  AOI21_X1  g0094(.A(new_n276), .B1(new_n294), .B2(KEYINPUT9), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n293), .B(KEYINPUT70), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT9), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n274), .A2(G200), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n295), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT10), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n289), .A2(new_n278), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n302), .B1(new_n292), .B2(new_n278), .ZN(new_n303));
  INV_X1    g0103(.A(new_n285), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n279), .A2(KEYINPUT3), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT3), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT7), .B1(new_n308), .B2(new_n237), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT7), .ZN(new_n310));
  AOI211_X1 g0110(.A(new_n310), .B(G20), .C1(new_n305), .C2(new_n307), .ZN(new_n311));
  OAI21_X1  g0111(.A(G68), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G58), .A2(G68), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n204), .A2(new_n205), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT75), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n237), .A2(new_n279), .ZN(new_n316));
  INV_X1    g0116(.A(G159), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n281), .A2(KEYINPUT75), .A3(G159), .ZN(new_n319));
  AOI22_X1  g0119(.A1(G20), .A2(new_n314), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n312), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT16), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n304), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AND3_X1   g0123(.A1(new_n306), .A2(KEYINPUT74), .A3(G33), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT74), .B1(new_n306), .B2(G33), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n305), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(new_n310), .A3(new_n237), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n306), .A2(G33), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT74), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(new_n279), .B2(KEYINPUT3), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n306), .A2(KEYINPUT74), .A3(G33), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n328), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT7), .B1(new_n332), .B2(G20), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n327), .A2(new_n333), .A3(G68), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n320), .A2(KEYINPUT76), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n314), .A2(G20), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n318), .A2(new_n319), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT76), .ZN(new_n338));
  OAI211_X1 g0138(.A(KEYINPUT16), .B(new_n334), .C1(new_n335), .C2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n303), .B1(new_n323), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n330), .A2(new_n331), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n268), .A2(new_n266), .ZN(new_n342));
  OR2_X1    g0142(.A1(new_n266), .A2(G226), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n341), .A2(new_n305), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G33), .A2(G87), .ZN(new_n345));
  XOR2_X1   g0145(.A(new_n345), .B(KEYINPUT77), .Z(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n272), .B1(new_n347), .B2(new_n259), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n260), .A2(G232), .A3(new_n262), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n348), .A2(new_n275), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n260), .B1(new_n344), .B2(new_n346), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n352), .A2(new_n272), .A3(new_n349), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n351), .B1(new_n353), .B2(G200), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n340), .A2(KEYINPUT17), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT17), .B1(new_n340), .B2(new_n354), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n323), .A2(new_n339), .ZN(new_n358));
  INV_X1    g0158(.A(new_n303), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n353), .A2(G179), .ZN(new_n361));
  INV_X1    g0161(.A(G169), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n361), .B1(new_n353), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n360), .A2(KEYINPUT18), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT18), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n362), .B1(new_n348), .B2(new_n350), .ZN(new_n366));
  INV_X1    g0166(.A(G179), .ZN(new_n367));
  NOR4_X1   g0167(.A1(new_n352), .A2(new_n349), .A3(new_n367), .A4(new_n272), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n365), .B1(new_n340), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n364), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n301), .A2(new_n357), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G33), .A2(G97), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n373), .B(KEYINPUT71), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n243), .A2(G1698), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(G226), .B2(G1698), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n374), .B1(new_n308), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n272), .B1(new_n377), .B2(new_n259), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT13), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n263), .A2(G238), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n379), .B1(new_n378), .B2(new_n380), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OR3_X1    g0183(.A1(new_n383), .A2(KEYINPUT72), .A3(new_n275), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n289), .A2(new_n203), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT12), .B1(new_n385), .B2(KEYINPUT73), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(KEYINPUT73), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n386), .B(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n280), .ZN(new_n389));
  INV_X1    g0189(.A(G77), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n389), .A2(new_n390), .B1(new_n239), .B2(new_n316), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n237), .A2(G68), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n285), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT11), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n393), .A2(new_n394), .B1(G68), .B2(new_n291), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n388), .B(new_n395), .C1(new_n394), .C2(new_n393), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n383), .B2(G200), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT72), .B1(new_n383), .B2(new_n275), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n384), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(G169), .B1(new_n381), .B2(new_n382), .ZN(new_n400));
  OR2_X1    g0200(.A1(new_n400), .A2(KEYINPUT14), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(KEYINPUT14), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n401), .B(new_n402), .C1(new_n367), .C2(new_n383), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n396), .ZN(new_n404));
  AOI22_X1  g0204(.A1(G20), .A2(new_n225), .B1(new_n278), .B2(new_n281), .ZN(new_n405));
  XOR2_X1   g0205(.A(KEYINPUT15), .B(G87), .Z(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n405), .B1(new_n389), .B2(new_n407), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(new_n285), .B1(G77), .B2(new_n291), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n225), .B2(new_n288), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n263), .A2(G244), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G238), .A2(G1698), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n265), .B(new_n412), .C1(new_n243), .C2(G1698), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n413), .B(new_n259), .C1(G107), .C2(new_n265), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n411), .A2(new_n414), .A3(new_n273), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n415), .A2(G179), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n362), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n410), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n415), .A2(G200), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n275), .B2(new_n415), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n421), .A2(new_n410), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  OR2_X1    g0223(.A1(new_n274), .A2(G179), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n274), .A2(new_n362), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n293), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n399), .A2(new_n404), .A3(new_n423), .A4(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT6), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT78), .ZN(new_n429));
  INV_X1    g0229(.A(G107), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n429), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  XNOR2_X1  g0231(.A(G97), .B(G107), .ZN(new_n432));
  MUX2_X1   g0232(.A(new_n431), .B(new_n429), .S(new_n432), .Z(new_n433));
  OAI22_X1  g0233(.A1(new_n433), .A2(new_n237), .B1(new_n390), .B2(new_n316), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n309), .A2(new_n311), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(new_n430), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n285), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n304), .B(new_n288), .C1(G1), .C2(new_n279), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G97), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n437), .B(new_n440), .C1(G97), .C2(new_n288), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n266), .A2(G244), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT79), .B1(new_n326), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT4), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT79), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n332), .A2(new_n445), .A3(G244), .A4(new_n266), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n443), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  OAI22_X1  g0247(.A1(new_n442), .A2(new_n444), .B1(new_n217), .B2(new_n266), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n265), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G283), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G45), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(G1), .ZN(new_n453));
  AND2_X1   g0253(.A1(KEYINPUT5), .A2(G41), .ZN(new_n454));
  NOR2_X1   g0254(.A1(KEYINPUT5), .A2(G41), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n260), .A2(new_n456), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n451), .A2(new_n259), .B1(G257), .B2(new_n457), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n456), .A2(new_n271), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n441), .B1(new_n460), .B2(G200), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT80), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n462), .B1(new_n460), .B2(new_n275), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n458), .A2(KEYINPUT80), .A3(G190), .A4(new_n459), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n406), .A2(new_n288), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT19), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n237), .B1(new_n374), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT81), .ZN(new_n469));
  INV_X1    g0269(.A(G97), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n216), .A2(new_n470), .A3(new_n430), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT81), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n472), .B(new_n237), .C1(new_n374), .C2(new_n467), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n469), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n467), .B1(new_n389), .B2(new_n470), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n332), .A2(new_n237), .A3(G68), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n466), .B1(new_n477), .B2(new_n285), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n439), .A2(new_n406), .ZN(new_n479));
  NOR2_X1   g0279(.A1(G238), .A2(G1698), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n480), .B1(new_n227), .B2(G1698), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n332), .A2(new_n481), .B1(G33), .B2(G116), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(new_n260), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n453), .A2(G250), .ZN(new_n484));
  AOI211_X1 g0284(.A(new_n259), .B(new_n484), .C1(new_n271), .C2(new_n453), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n478), .A2(new_n479), .B1(new_n367), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n486), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n362), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n439), .A2(G87), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n478), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(G200), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(G190), .B2(new_n486), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n487), .A2(new_n489), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT22), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n237), .A2(G87), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n496), .B1(new_n308), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n332), .A2(KEYINPUT22), .A3(new_n237), .A4(G87), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n237), .A2(G33), .A3(G116), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT83), .ZN(new_n501));
  XNOR2_X1  g0301(.A(new_n500), .B(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n430), .A2(G20), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT23), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n503), .B(new_n504), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n502), .A2(KEYINPUT84), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT84), .B1(new_n502), .B2(new_n505), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n498), .B(new_n499), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT24), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n502), .A2(new_n505), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT84), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n502), .A2(KEYINPUT84), .A3(new_n505), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n515), .A2(KEYINPUT24), .A3(new_n498), .A4(new_n499), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n510), .A2(new_n516), .A3(new_n285), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n503), .A2(G1), .A3(new_n286), .ZN(new_n518));
  XNOR2_X1  g0318(.A(new_n518), .B(KEYINPUT25), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n457), .A2(G264), .ZN(new_n521));
  OR2_X1    g0321(.A1(new_n521), .A2(KEYINPUT85), .ZN(new_n522));
  INV_X1    g0322(.A(new_n459), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n217), .A2(new_n266), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n332), .B(new_n524), .C1(G257), .C2(new_n266), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G294), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n523), .B1(new_n527), .B2(new_n259), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n521), .A2(KEYINPUT85), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n522), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G200), .ZN(new_n531));
  INV_X1    g0331(.A(new_n530), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G190), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n439), .A2(G107), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n520), .A2(new_n531), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n460), .A2(new_n362), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n458), .A2(new_n367), .A3(new_n459), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(new_n441), .A3(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n465), .A2(new_n495), .A3(new_n535), .A4(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n332), .B1(G264), .B2(new_n266), .ZN(new_n540));
  NOR2_X1   g0340(.A1(G257), .A2(G1698), .ZN(new_n541));
  INV_X1    g0341(.A(G303), .ZN(new_n542));
  OAI22_X1  g0342(.A1(new_n540), .A2(new_n541), .B1(new_n542), .B2(new_n265), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n259), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n260), .A2(G270), .A3(new_n456), .ZN(new_n545));
  XNOR2_X1  g0345(.A(new_n545), .B(KEYINPUT82), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n459), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n289), .A2(new_n222), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n450), .B(new_n237), .C1(G33), .C2(new_n470), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n549), .B(new_n285), .C1(new_n237), .C2(G116), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT20), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n550), .A2(new_n551), .ZN(new_n553));
  OAI221_X1 g0353(.A(new_n548), .B1(new_n222), .B2(new_n438), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n547), .A2(G169), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT21), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AND4_X1   g0357(.A1(G179), .A2(new_n544), .A3(new_n459), .A4(new_n546), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n554), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n547), .A2(KEYINPUT21), .A3(G169), .A4(new_n554), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n517), .A2(new_n534), .A3(new_n519), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n530), .A2(new_n362), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n532), .A2(new_n367), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n547), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n554), .B1(new_n566), .B2(G190), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n492), .B2(new_n566), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n561), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  NOR4_X1   g0369(.A1(new_n372), .A2(new_n427), .A3(new_n539), .A4(new_n569), .ZN(G372));
  INV_X1    g0370(.A(new_n426), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT88), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n301), .B(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT87), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT18), .B1(new_n360), .B2(new_n363), .ZN(new_n575));
  NOR3_X1   g0375(.A1(new_n340), .A2(new_n369), .A3(new_n365), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n364), .A2(new_n370), .A3(KEYINPUT87), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n399), .A2(new_n419), .B1(new_n403), .B2(new_n396), .ZN(new_n580));
  INV_X1    g0380(.A(new_n357), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n571), .B1(new_n573), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n372), .A2(new_n427), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n487), .A2(new_n489), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n491), .A2(new_n494), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT26), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n587), .A2(new_n538), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n538), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT26), .B1(new_n495), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n585), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT86), .B1(new_n561), .B2(new_n565), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n561), .A2(new_n565), .A3(KEYINPUT86), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n539), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n584), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n583), .A2(new_n596), .ZN(G369));
  NAND2_X1  g0397(.A1(new_n287), .A2(new_n237), .ZN(new_n598));
  OR2_X1    g0398(.A1(new_n598), .A2(KEYINPUT27), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(KEYINPUT27), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(G213), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(G343), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n565), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n562), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n535), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n604), .B1(new_n606), .B2(new_n565), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n561), .A2(new_n603), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n609), .A2(new_n604), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n554), .A2(new_n603), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n561), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n561), .A2(new_n612), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n568), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(G330), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n607), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n610), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g0419(.A(new_n619), .B(KEYINPUT89), .Z(G399));
  INV_X1    g0420(.A(new_n232), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n621), .A2(G41), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n471), .A2(G116), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(G1), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n240), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n625), .B1(new_n626), .B2(new_n623), .ZN(new_n627));
  XNOR2_X1  g0427(.A(new_n627), .B(KEYINPUT28), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT92), .ZN(new_n629));
  OR3_X1    g0429(.A1(new_n539), .A2(new_n593), .A3(new_n594), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n588), .B1(new_n587), .B2(new_n538), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n495), .A2(new_n590), .A3(KEYINPUT26), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n631), .A2(new_n632), .B1(new_n489), .B2(new_n487), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n603), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n629), .B1(new_n634), .B2(KEYINPUT29), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n561), .A2(new_n565), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n539), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n603), .B1(new_n637), .B2(new_n633), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT29), .ZN(new_n639));
  INV_X1    g0439(.A(new_n603), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n595), .B2(new_n592), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT29), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(KEYINPUT92), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n635), .A2(new_n639), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n532), .B1(new_n458), .B2(new_n459), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT91), .ZN(new_n646));
  AOI21_X1  g0446(.A(G179), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n460), .A2(new_n530), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(KEYINPUT91), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n647), .A2(new_n488), .A3(new_n649), .A4(new_n547), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n532), .A2(new_n558), .A3(new_n486), .A4(new_n458), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT90), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT30), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n653), .B1(new_n651), .B2(new_n652), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT31), .B1(new_n657), .B2(new_n603), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n539), .A2(new_n569), .A3(new_n603), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n657), .A2(KEYINPUT31), .A3(new_n603), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n616), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n644), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n628), .B1(new_n665), .B2(G1), .ZN(G364));
  INV_X1    g0466(.A(new_n617), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n286), .A2(G20), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(G45), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n623), .A2(G1), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n615), .A2(new_n616), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT93), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n237), .A2(G179), .ZN(new_n674));
  NOR2_X1   g0474(.A1(G190), .A2(G200), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT32), .B1(new_n676), .B2(new_n317), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n237), .A2(new_n367), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT96), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT96), .B1(new_n237), .B2(new_n367), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(new_n675), .A3(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n275), .A2(G200), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n680), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  OAI221_X1 g0484(.A(new_n677), .B1(new_n682), .B2(new_n226), .C1(new_n202), .C2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n674), .A2(new_n275), .A3(G200), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n430), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n308), .ZN(new_n688));
  OR3_X1    g0488(.A1(new_n676), .A2(KEYINPUT32), .A3(new_n317), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n237), .B1(new_n683), .B2(new_n367), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G97), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n678), .A2(new_n275), .A3(G200), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G68), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n688), .A2(new_n689), .A3(new_n692), .A4(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n678), .A2(G200), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(new_n275), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n239), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n674), .A2(G190), .A3(G200), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n216), .ZN(new_n702));
  NOR4_X1   g0502(.A1(new_n685), .A2(new_n696), .A3(new_n700), .A4(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(G317), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n693), .B1(KEYINPUT33), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(KEYINPUT33), .B2(new_n704), .ZN(new_n706));
  INV_X1    g0506(.A(G322), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n698), .A2(G326), .B1(new_n691), .B2(G294), .ZN(new_n708));
  OAI221_X1 g0508(.A(new_n706), .B1(new_n707), .B2(new_n684), .C1(new_n708), .C2(KEYINPUT97), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n265), .B1(new_n708), .B2(KEYINPUT97), .ZN(new_n710));
  INV_X1    g0510(.A(new_n676), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G329), .ZN(new_n712));
  INV_X1    g0512(.A(G283), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n710), .B(new_n712), .C1(new_n713), .C2(new_n686), .ZN(new_n714));
  INV_X1    g0514(.A(new_n701), .ZN(new_n715));
  AOI211_X1 g0515(.A(new_n709), .B(new_n714), .C1(G303), .C2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n682), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G311), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n703), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT98), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n236), .B1(G20), .B2(new_n362), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(G13), .A2(G33), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G20), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n615), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n670), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n332), .A2(new_n621), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(new_n626), .B2(G45), .ZN(new_n729));
  XOR2_X1   g0529(.A(new_n729), .B(KEYINPUT94), .Z(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n452), .B2(new_n253), .ZN(new_n731));
  INV_X1    g0531(.A(G355), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n265), .A2(new_n232), .ZN(new_n733));
  OAI221_X1 g0533(.A(new_n731), .B1(G116), .B2(new_n232), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n725), .A2(new_n721), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT95), .Z(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n722), .A2(new_n726), .A3(new_n727), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n673), .A2(new_n738), .ZN(G396));
  NAND2_X1  g0539(.A1(new_n410), .A2(new_n603), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n423), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT102), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n423), .A2(KEYINPUT102), .A3(new_n740), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(new_n418), .B2(new_n640), .ZN(new_n746));
  OR3_X1    g0546(.A1(new_n634), .A2(KEYINPUT103), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(KEYINPUT103), .B1(new_n634), .B2(new_n746), .ZN(new_n748));
  INV_X1    g0548(.A(new_n745), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n640), .B(new_n749), .C1(new_n595), .C2(new_n592), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n747), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n751), .A2(new_n663), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n663), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n752), .A2(new_n670), .A3(new_n753), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n746), .A2(new_n724), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n721), .A2(new_n723), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT99), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n390), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n694), .A2(KEYINPUT100), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n694), .A2(KEYINPUT100), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n713), .ZN(new_n762));
  INV_X1    g0562(.A(G294), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n692), .B1(new_n684), .B2(new_n763), .C1(new_n699), .C2(new_n542), .ZN(new_n764));
  INV_X1    g0564(.A(G311), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n686), .A2(new_n216), .B1(new_n676), .B2(new_n765), .ZN(new_n766));
  NOR4_X1   g0566(.A1(new_n762), .A2(new_n764), .A3(new_n265), .A4(new_n766), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n767), .B1(new_n430), .B2(new_n701), .C1(new_n222), .C2(new_n682), .ZN(new_n768));
  INV_X1    g0568(.A(new_n684), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n769), .A2(G143), .B1(G150), .B2(new_n694), .ZN(new_n770));
  INV_X1    g0570(.A(G137), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n770), .B1(new_n771), .B2(new_n699), .C1(new_n317), .C2(new_n682), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT34), .Z(new_n773));
  INV_X1    g0573(.A(G132), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n332), .B1(new_n774), .B2(new_n676), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT101), .Z(new_n776));
  INV_X1    g0576(.A(new_n686), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G68), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n691), .A2(G58), .B1(new_n715), .B2(G50), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n768), .B1(new_n773), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n721), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n755), .A2(new_n727), .A3(new_n758), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n754), .A2(new_n783), .ZN(G384));
  NOR2_X1   g0584(.A1(new_n668), .A2(new_n261), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n403), .A2(new_n396), .A3(new_n640), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT107), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT38), .ZN(new_n789));
  INV_X1    g0589(.A(new_n601), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n360), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(new_n579), .B2(new_n357), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n340), .A2(new_n354), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n791), .A2(KEYINPUT87), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(KEYINPUT37), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n360), .A2(new_n363), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n796), .A2(new_n791), .A3(new_n793), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n791), .A2(new_n793), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n799), .A2(new_n574), .A3(KEYINPUT37), .A4(new_n796), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n789), .B1(new_n792), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT108), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n320), .B(KEYINPUT76), .ZN(new_n804));
  AOI21_X1  g0604(.A(KEYINPUT16), .B1(new_n804), .B2(new_n334), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n339), .A2(new_n285), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n359), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n369), .A2(new_n601), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n793), .ZN(new_n810));
  OAI21_X1  g0610(.A(KEYINPUT37), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(KEYINPUT37), .B2(new_n797), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT106), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n357), .A2(new_n371), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n807), .A2(new_n790), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n813), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  AOI211_X1 g0617(.A(KEYINPUT106), .B(new_n815), .C1(new_n357), .C2(new_n371), .ZN(new_n818));
  OAI211_X1 g0618(.A(KEYINPUT38), .B(new_n812), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n802), .A2(new_n803), .A3(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT39), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n802), .A2(KEYINPUT108), .A3(new_n819), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n812), .B1(new_n817), .B2(new_n818), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n789), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n826), .A2(KEYINPUT39), .A3(new_n819), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n822), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(KEYINPUT109), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n823), .A2(KEYINPUT39), .A3(new_n819), .A4(new_n826), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT109), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n830), .A2(new_n831), .A3(new_n822), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n788), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n579), .A2(new_n790), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n396), .A2(new_n603), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n403), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n404), .A2(new_n399), .A3(new_n835), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n838), .B1(new_n839), .B2(KEYINPUT105), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n838), .A2(KEYINPUT105), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n418), .A2(new_n603), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n843), .B1(new_n750), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n826), .A2(new_n819), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n834), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n833), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n635), .A2(new_n584), .A3(new_n639), .A4(new_n643), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n583), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n850), .B(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n746), .B1(new_n840), .B2(new_n842), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n660), .B2(new_n661), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n847), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT40), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n857), .B1(new_n802), .B2(new_n819), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n657), .A2(new_n603), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT31), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OR3_X1    g0664(.A1(new_n539), .A2(new_n569), .A3(new_n603), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n864), .A2(new_n865), .A3(new_n661), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n584), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n861), .B(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n868), .A2(new_n616), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n785), .B1(new_n853), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT110), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n853), .B2(new_n869), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n433), .B(KEYINPUT104), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT35), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n237), .B(new_n236), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n875), .B(G116), .C1(new_n874), .C2(new_n873), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT36), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n240), .A2(new_n225), .A3(new_n313), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n203), .B2(new_n209), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(G1), .A3(new_n286), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n872), .A2(new_n877), .A3(new_n880), .ZN(G367));
  INV_X1    g0681(.A(new_n728), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n735), .B1(new_n232), .B2(new_n407), .C1(new_n249), .C2(new_n882), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT112), .Z(new_n884));
  NOR2_X1   g0684(.A1(new_n701), .A2(new_n222), .ZN(new_n885));
  AOI22_X1  g0685(.A1(KEYINPUT46), .A2(new_n885), .B1(new_n698), .B2(G311), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n886), .B(new_n326), .C1(new_n542), .C2(new_n684), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(G107), .B2(new_n691), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n763), .B2(new_n761), .ZN(new_n889));
  OAI22_X1  g0689(.A1(new_n885), .A2(KEYINPUT46), .B1(new_n470), .B2(new_n686), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI221_X1 g0691(.A(new_n891), .B1(new_n713), .B2(new_n682), .C1(new_n704), .C2(new_n676), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n698), .A2(G143), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n203), .B2(new_n690), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n265), .B1(new_n701), .B2(new_n202), .ZN(new_n895));
  INV_X1    g0695(.A(G150), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n684), .A2(new_n896), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n226), .A2(new_n686), .B1(new_n771), .B2(new_n676), .ZN(new_n898));
  NOR4_X1   g0698(.A1(new_n894), .A2(new_n895), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  OAI221_X1 g0699(.A(new_n899), .B1(new_n317), .B2(new_n761), .C1(new_n208), .C2(new_n682), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n892), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT47), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n670), .B(new_n884), .C1(new_n902), .C2(new_n721), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n491), .A2(new_n640), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n495), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n585), .B2(new_n904), .ZN(new_n906));
  INV_X1    g0706(.A(new_n725), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n903), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n618), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n441), .A2(new_n603), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n465), .A2(new_n538), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n538), .B2(new_n640), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n609), .A2(new_n913), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT42), .Z(new_n916));
  OAI21_X1  g0716(.A(new_n538), .B1(new_n912), .B2(new_n565), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n640), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n906), .A2(KEYINPUT43), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n914), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n906), .A2(KEYINPUT43), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n919), .A2(new_n914), .A3(new_n920), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n923), .B1(new_n922), .B2(new_n924), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n669), .A2(G1), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n610), .A2(new_n913), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT45), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT45), .B1(new_n610), .B2(new_n913), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OR3_X1    g0734(.A1(new_n610), .A2(KEYINPUT44), .A3(new_n913), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT44), .B1(new_n610), .B2(new_n913), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n934), .A2(new_n937), .A3(new_n618), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n932), .A2(new_n933), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n935), .A2(new_n936), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n910), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n607), .B(new_n608), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT111), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n617), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT111), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n667), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n665), .B1(new_n942), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n622), .B(KEYINPUT41), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n929), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n909), .B1(new_n928), .B2(new_n952), .ZN(G387));
  AOI22_X1  g0753(.A1(G303), .A2(new_n717), .B1(new_n769), .B2(G317), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n954), .B1(new_n707), .B2(new_n699), .C1(new_n761), .C2(new_n765), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT48), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n956), .B1(new_n713), .B2(new_n690), .C1(new_n763), .C2(new_n701), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT49), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n711), .A2(G326), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n777), .A2(G116), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n959), .A2(new_n326), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(new_n958), .B2(new_n957), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n226), .A2(new_n701), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n278), .B2(new_n694), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n896), .B2(new_n676), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n699), .A2(new_n317), .B1(new_n407), .B2(new_n690), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n682), .A2(new_n203), .B1(new_n470), .B2(new_n686), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n332), .B1(new_n684), .B2(new_n239), .ZN(new_n969));
  NOR4_X1   g0769(.A1(new_n966), .A2(new_n967), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n721), .B1(new_n963), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n246), .A2(G45), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT113), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n278), .A2(new_n239), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT50), .Z(new_n975));
  AOI21_X1  g0775(.A(G45), .B1(G68), .B2(G77), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(new_n624), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n973), .A2(new_n728), .A3(new_n977), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(G107), .B2(new_n232), .C1(new_n624), .C2(new_n733), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n736), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n971), .A2(new_n727), .A3(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT114), .Z(new_n982));
  OR2_X1    g0782(.A1(new_n607), .A2(new_n907), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n982), .A2(new_n983), .B1(new_n929), .B2(new_n948), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n949), .A2(new_n664), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n665), .A2(new_n948), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n985), .A2(new_n622), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n984), .A2(new_n987), .ZN(G393));
  OR2_X1    g0788(.A1(new_n942), .A2(new_n986), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n623), .B1(new_n942), .B2(new_n986), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n938), .A2(new_n929), .A3(new_n941), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n769), .A2(G311), .B1(G317), .B2(new_n698), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n995));
  OAI22_X1  g0795(.A1(new_n994), .A2(new_n995), .B1(new_n222), .B2(new_n690), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n687), .B1(new_n994), .B2(new_n995), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n997), .B(new_n308), .C1(new_n542), .C2(new_n761), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n996), .B(new_n998), .C1(G322), .C2(new_n711), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n713), .B2(new_n701), .C1(new_n763), .C2(new_n682), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n690), .A2(new_n390), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n769), .A2(G159), .B1(G150), .B2(new_n698), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT51), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1003), .A2(new_n326), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n761), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n209), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n717), .A2(new_n278), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n203), .A2(new_n701), .B1(new_n686), .B2(new_n216), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(G143), .B2(new_n711), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1004), .A2(new_n1006), .A3(new_n1007), .A4(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1000), .B1(new_n1001), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n670), .B1(new_n1011), .B2(new_n721), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n735), .B1(new_n470), .B2(new_n232), .C1(new_n257), .C2(new_n882), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(new_n907), .C2(new_n913), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n992), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n991), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT116), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n991), .A2(KEYINPUT116), .A3(new_n1015), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(G390));
  NAND3_X1  g0820(.A1(new_n866), .A2(G330), .A3(new_n746), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n843), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n843), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n662), .A2(new_n746), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n750), .A2(new_n845), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n844), .B1(new_n638), .B2(new_n749), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1022), .A2(new_n1024), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n584), .A2(G330), .A3(new_n866), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n851), .A2(new_n583), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1026), .A2(new_n1023), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n788), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n829), .A2(new_n1036), .A3(new_n832), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n802), .A2(new_n819), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n1028), .B2(new_n843), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1039), .A2(new_n787), .ZN(new_n1040));
  AND3_X1   g0840(.A1(new_n1037), .A2(new_n1040), .A3(new_n1024), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1024), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1034), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1024), .ZN(new_n1044));
  AND3_X1   g0844(.A1(new_n830), .A2(new_n831), .A3(new_n822), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n831), .B1(new_n830), .B2(new_n822), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n787), .B1(new_n1026), .B2(new_n1023), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1039), .A2(new_n787), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1044), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1037), .A2(new_n1040), .A3(new_n1024), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1032), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1043), .A2(new_n1053), .A3(new_n622), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n829), .A2(new_n832), .A3(new_n723), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n1005), .A2(G137), .B1(G128), .B2(new_n698), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n774), .B2(new_n684), .C1(new_n317), .C2(new_n690), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n711), .A2(G125), .ZN(new_n1058));
  XOR2_X1   g0858(.A(KEYINPUT54), .B(G143), .Z(new_n1059));
  AND2_X1   g0859(.A1(new_n717), .A2(new_n1059), .ZN(new_n1060));
  NOR4_X1   g0860(.A1(new_n1057), .A2(new_n308), .A3(new_n1058), .A4(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n701), .A2(new_n896), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT53), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1061), .B(new_n1063), .C1(new_n208), .C2(new_n686), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT117), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n702), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n308), .B1(new_n676), .B2(new_n763), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n717), .A2(G97), .B1(G283), .B2(new_n698), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n761), .B2(new_n430), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT118), .Z(new_n1070));
  AOI211_X1 g0870(.A(new_n1067), .B(new_n1070), .C1(G116), .C2(new_n769), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1001), .ZN(new_n1072));
  AND4_X1   g0872(.A1(new_n1066), .A2(new_n1071), .A3(new_n778), .A4(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n721), .B1(new_n1065), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n278), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n670), .B1(new_n757), .B2(new_n1075), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n1055), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1077), .B1(new_n1078), .B2(new_n929), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1054), .A2(new_n1079), .ZN(G378));
  NAND2_X1  g0880(.A1(new_n1053), .A2(new_n1033), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n860), .ZN(new_n1082));
  AOI21_X1  g0882(.A(KEYINPUT40), .B1(new_n855), .B2(new_n847), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n1082), .A2(new_n1083), .A3(new_n616), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n833), .B2(new_n849), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n573), .A2(new_n426), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n296), .A2(new_n790), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1087), .B(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1086), .B(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n787), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n858), .A2(G330), .A3(new_n860), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1091), .A2(new_n1092), .A3(new_n848), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1085), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1085), .A2(new_n1093), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1090), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1081), .A2(KEYINPUT57), .A3(new_n1094), .A4(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n622), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1085), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1090), .B1(new_n1085), .B2(new_n1093), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT57), .B1(new_n1102), .B2(new_n1081), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1097), .A2(new_n929), .A3(new_n1094), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n670), .B1(new_n1096), .B2(new_n723), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n684), .A2(new_n430), .B1(new_n203), .B2(new_n690), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n964), .A2(G41), .A3(new_n332), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT119), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n686), .A2(new_n202), .B1(new_n676), .B2(new_n713), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT120), .Z(new_n1114));
  AOI211_X1 g0914(.A(new_n1107), .B(new_n1114), .C1(G116), .C2(new_n698), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1115), .B1(new_n470), .B2(new_n693), .C1(new_n407), .C2(new_n682), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT58), .Z(new_n1117));
  NAND2_X1  g0917(.A1(new_n715), .A2(new_n1059), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT121), .Z(new_n1119));
  NAND2_X1  g0919(.A1(new_n717), .A2(G137), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n769), .A2(G128), .B1(G132), .B2(new_n694), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n698), .A2(G125), .B1(new_n691), .B2(G150), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT59), .ZN(new_n1124));
  AOI211_X1 g0924(.A(G33), .B(G41), .C1(new_n711), .C2(G124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n317), .B2(new_n686), .ZN(new_n1126));
  AOI21_X1  g0926(.A(G41), .B1(new_n341), .B2(G33), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1124), .A2(new_n1126), .B1(G50), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n721), .B1(new_n1117), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n756), .A2(new_n208), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1106), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1105), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1104), .A2(new_n1132), .ZN(G375));
  OAI221_X1 g0933(.A(new_n308), .B1(new_n713), .B2(new_n684), .C1(new_n761), .C2(new_n222), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n698), .A2(G294), .B1(new_n691), .B2(new_n406), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1135), .B1(new_n390), .B2(new_n686), .C1(new_n542), .C2(new_n676), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n701), .A2(new_n470), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n682), .A2(new_n430), .ZN(new_n1138));
  NOR4_X1   g0938(.A1(new_n1134), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n682), .A2(new_n896), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n769), .A2(G137), .B1(G159), .B2(new_n715), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n698), .A2(G132), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n326), .B1(G128), .B2(new_n711), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n691), .A2(G50), .B1(new_n777), .B2(G58), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1140), .B(new_n1145), .C1(new_n1005), .C2(new_n1059), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n721), .B1(new_n1139), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n757), .A2(new_n203), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1147), .A2(new_n727), .A3(new_n1148), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT122), .Z(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n843), .B2(new_n723), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n1030), .B2(new_n929), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1027), .A2(new_n1032), .A3(new_n1029), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n951), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1152), .B1(new_n1154), .B2(new_n1052), .ZN(G381));
  INV_X1    g0955(.A(KEYINPUT123), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1054), .A2(new_n1079), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1156), .B1(new_n1054), .B2(new_n1079), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(G375), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n952), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n927), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1018), .A2(new_n1162), .A3(new_n909), .A4(new_n1019), .ZN(new_n1163));
  OR2_X1    g0963(.A1(G393), .A2(G396), .ZN(new_n1164));
  NOR4_X1   g0964(.A1(new_n1163), .A2(G384), .A3(G381), .A4(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1160), .A2(new_n1165), .ZN(G407));
  OAI21_X1  g0966(.A(new_n1160), .B1(new_n1165), .B2(new_n602), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(G213), .ZN(G409));
  OAI211_X1 g0968(.A(G378), .B(new_n1132), .C1(new_n1099), .C2(new_n1103), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1081), .A2(new_n951), .A3(new_n1094), .A4(new_n1097), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1170), .A2(new_n1105), .A3(new_n1131), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n1158), .B2(new_n1157), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(G213), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1174), .A2(G343), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT124), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1027), .A2(new_n1032), .A3(KEYINPUT60), .A4(new_n1029), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1034), .A2(new_n1179), .A3(new_n622), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT60), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1153), .A2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g0982(.A(G384), .B(new_n1152), .C1(new_n1180), .C2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1153), .A2(new_n1181), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1185), .A2(new_n622), .A3(new_n1034), .A4(new_n1179), .ZN(new_n1186));
  AOI21_X1  g0986(.A(G384), .B1(new_n1186), .B2(new_n1152), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1178), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1186), .A2(new_n1152), .ZN(new_n1189));
  INV_X1    g0989(.A(G384), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1191), .A2(KEYINPUT124), .A3(new_n1183), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1188), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1175), .A2(G2897), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1191), .A2(new_n1183), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1195), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1177), .A2(new_n1196), .A3(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1173), .A2(new_n1176), .A3(new_n1194), .ZN(new_n1201));
  AND2_X1   g1001(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT61), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1173), .A2(new_n1176), .A3(new_n1194), .A4(new_n1206), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1200), .A2(new_n1203), .A3(new_n1204), .A4(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(G390), .A2(G387), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(G393), .A2(G396), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1164), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(new_n1163), .A3(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1211), .B1(new_n1209), .B2(new_n1163), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1213), .A2(new_n1214), .A3(KEYINPUT127), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT127), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1209), .A2(new_n1163), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1211), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1216), .B1(new_n1219), .B2(new_n1212), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1215), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1208), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1201), .A2(KEYINPUT125), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(KEYINPUT63), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1173), .A2(new_n1176), .B1(new_n1198), .B2(new_n1197), .ZN(new_n1225));
  AOI21_X1  g1025(.A(KEYINPUT61), .B1(new_n1225), .B2(new_n1196), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1219), .A2(new_n1212), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT63), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1201), .A2(KEYINPUT125), .A3(new_n1229), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1224), .A2(new_n1226), .A3(new_n1228), .A4(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1222), .A2(new_n1231), .ZN(G405));
  AOI21_X1  g1032(.A(new_n1159), .B1(new_n1104), .B2(new_n1132), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1169), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n1197), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1194), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1236), .A2(new_n1227), .A3(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1227), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(G402));
endmodule


