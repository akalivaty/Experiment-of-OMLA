

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U549 ( .A(n709), .B(KEYINPUT29), .Z(n516) );
  XOR2_X1 U550 ( .A(n809), .B(KEYINPUT105), .Z(n517) );
  NOR2_X1 U551 ( .A1(n802), .A2(n750), .ZN(n518) );
  NOR2_X1 U552 ( .A1(G299), .A2(n685), .ZN(n686) );
  XNOR2_X1 U553 ( .A(KEYINPUT30), .B(KEYINPUT100), .ZN(n715) );
  XNOR2_X1 U554 ( .A(n716), .B(n715), .ZN(n717) );
  OR2_X1 U555 ( .A1(n733), .A2(n732), .ZN(n734) );
  INV_X1 U556 ( .A(KEYINPUT32), .ZN(n736) );
  NAND2_X1 U557 ( .A1(G8), .A2(n728), .ZN(n802) );
  AND2_X1 U558 ( .A1(n797), .A2(n800), .ZN(n798) );
  NAND2_X1 U559 ( .A1(n823), .A2(n925), .ZN(n810) );
  AND2_X2 U560 ( .A1(n532), .A2(G2104), .ZN(n886) );
  NOR2_X1 U561 ( .A1(G651), .A2(G543), .ZN(n638) );
  NAND2_X1 U562 ( .A1(G91), .A2(n638), .ZN(n520) );
  XOR2_X1 U563 ( .A(KEYINPUT0), .B(G543), .Z(n615) );
  INV_X1 U564 ( .A(G651), .ZN(n525) );
  NOR2_X1 U565 ( .A1(n615), .A2(n525), .ZN(n641) );
  NAND2_X1 U566 ( .A1(G78), .A2(n641), .ZN(n519) );
  NAND2_X1 U567 ( .A1(n520), .A2(n519), .ZN(n524) );
  NOR2_X1 U568 ( .A1(G651), .A2(n615), .ZN(n521) );
  XOR2_X2 U569 ( .A(KEYINPUT65), .B(n521), .Z(n642) );
  NAND2_X1 U570 ( .A1(G53), .A2(n642), .ZN(n522) );
  XNOR2_X1 U571 ( .A(KEYINPUT71), .B(n522), .ZN(n523) );
  NOR2_X1 U572 ( .A1(n524), .A2(n523), .ZN(n529) );
  NOR2_X1 U573 ( .A1(G543), .A2(n525), .ZN(n527) );
  XNOR2_X1 U574 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n526) );
  XNOR2_X1 U575 ( .A(n527), .B(n526), .ZN(n637) );
  NAND2_X1 U576 ( .A1(n637), .A2(G65), .ZN(n528) );
  NAND2_X1 U577 ( .A1(n529), .A2(n528), .ZN(G299) );
  INV_X1 U578 ( .A(G2105), .ZN(n530) );
  NOR2_X1 U579 ( .A1(n530), .A2(G2104), .ZN(n604) );
  NAND2_X1 U580 ( .A1(G125), .A2(n604), .ZN(n531) );
  XNOR2_X1 U581 ( .A(n531), .B(KEYINPUT66), .ZN(n535) );
  INV_X1 U582 ( .A(G2105), .ZN(n532) );
  NAND2_X1 U583 ( .A1(G101), .A2(n886), .ZN(n533) );
  XOR2_X1 U584 ( .A(KEYINPUT23), .B(n533), .Z(n534) );
  NAND2_X1 U585 ( .A1(n535), .A2(n534), .ZN(n540) );
  NOR2_X1 U586 ( .A1(G2104), .A2(G2105), .ZN(n536) );
  XOR2_X2 U587 ( .A(KEYINPUT17), .B(n536), .Z(n887) );
  NAND2_X1 U588 ( .A1(n887), .A2(G137), .ZN(n538) );
  AND2_X1 U589 ( .A1(G2104), .A2(G2105), .ZN(n882) );
  NAND2_X1 U590 ( .A1(G113), .A2(n882), .ZN(n537) );
  NAND2_X1 U591 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U592 ( .A1(n540), .A2(n539), .ZN(G160) );
  NAND2_X1 U593 ( .A1(G85), .A2(n638), .ZN(n542) );
  NAND2_X1 U594 ( .A1(G72), .A2(n641), .ZN(n541) );
  NAND2_X1 U595 ( .A1(n542), .A2(n541), .ZN(n546) );
  NAND2_X1 U596 ( .A1(G60), .A2(n637), .ZN(n544) );
  NAND2_X1 U597 ( .A1(G47), .A2(n642), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n544), .A2(n543), .ZN(n545) );
  OR2_X1 U599 ( .A1(n546), .A2(n545), .ZN(G290) );
  INV_X1 U600 ( .A(G132), .ZN(G219) );
  INV_X1 U601 ( .A(G82), .ZN(G220) );
  INV_X1 U602 ( .A(G57), .ZN(G237) );
  INV_X1 U603 ( .A(G120), .ZN(G236) );
  NAND2_X1 U604 ( .A1(G63), .A2(n637), .ZN(n548) );
  NAND2_X1 U605 ( .A1(G51), .A2(n642), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U607 ( .A(KEYINPUT6), .B(n549), .ZN(n556) );
  NAND2_X1 U608 ( .A1(n638), .A2(G89), .ZN(n550) );
  XNOR2_X1 U609 ( .A(n550), .B(KEYINPUT4), .ZN(n552) );
  NAND2_X1 U610 ( .A1(G76), .A2(n641), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U612 ( .A(KEYINPUT74), .B(n553), .Z(n554) );
  XNOR2_X1 U613 ( .A(KEYINPUT5), .B(n554), .ZN(n555) );
  NOR2_X1 U614 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U615 ( .A(KEYINPUT7), .B(n557), .Z(G168) );
  XOR2_X1 U616 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U617 ( .A1(G94), .A2(G452), .ZN(n558) );
  XOR2_X1 U618 ( .A(KEYINPUT70), .B(n558), .Z(G173) );
  NAND2_X1 U619 ( .A1(G7), .A2(G661), .ZN(n559) );
  XNOR2_X1 U620 ( .A(n559), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U621 ( .A(G223), .ZN(n828) );
  NAND2_X1 U622 ( .A1(n828), .A2(G567), .ZN(n560) );
  XOR2_X1 U623 ( .A(KEYINPUT11), .B(n560), .Z(G234) );
  XOR2_X1 U624 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n562) );
  NAND2_X1 U625 ( .A1(G56), .A2(n637), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n562), .B(n561), .ZN(n569) );
  XNOR2_X1 U627 ( .A(KEYINPUT13), .B(KEYINPUT73), .ZN(n567) );
  NAND2_X1 U628 ( .A1(n638), .A2(G81), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT12), .ZN(n565) );
  NAND2_X1 U630 ( .A1(G68), .A2(n641), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  NOR2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n642), .A2(G43), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n923) );
  INV_X1 U636 ( .A(G860), .ZN(n594) );
  OR2_X1 U637 ( .A1(n923), .A2(n594), .ZN(G153) );
  NAND2_X1 U638 ( .A1(G64), .A2(n637), .ZN(n573) );
  NAND2_X1 U639 ( .A1(G52), .A2(n642), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U641 ( .A(KEYINPUT68), .B(n574), .ZN(n580) );
  NAND2_X1 U642 ( .A1(G90), .A2(n638), .ZN(n576) );
  NAND2_X1 U643 ( .A1(G77), .A2(n641), .ZN(n575) );
  NAND2_X1 U644 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U645 ( .A(KEYINPUT69), .B(n577), .ZN(n578) );
  XNOR2_X1 U646 ( .A(KEYINPUT9), .B(n578), .ZN(n579) );
  NOR2_X1 U647 ( .A1(n580), .A2(n579), .ZN(G171) );
  INV_X1 U648 ( .A(G171), .ZN(G301) );
  NAND2_X1 U649 ( .A1(G868), .A2(G301), .ZN(n589) );
  NAND2_X1 U650 ( .A1(G79), .A2(n641), .ZN(n582) );
  NAND2_X1 U651 ( .A1(G54), .A2(n642), .ZN(n581) );
  NAND2_X1 U652 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U653 ( .A1(G66), .A2(n637), .ZN(n584) );
  NAND2_X1 U654 ( .A1(G92), .A2(n638), .ZN(n583) );
  NAND2_X1 U655 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U656 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U657 ( .A(n587), .B(KEYINPUT15), .ZN(n920) );
  INV_X1 U658 ( .A(G868), .ZN(n656) );
  NAND2_X1 U659 ( .A1(n920), .A2(n656), .ZN(n588) );
  NAND2_X1 U660 ( .A1(n589), .A2(n588), .ZN(G284) );
  NOR2_X1 U661 ( .A1(G868), .A2(G299), .ZN(n590) );
  XOR2_X1 U662 ( .A(KEYINPUT75), .B(n590), .Z(n592) );
  NOR2_X1 U663 ( .A1(G286), .A2(n656), .ZN(n591) );
  NOR2_X1 U664 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U665 ( .A(KEYINPUT76), .B(n593), .ZN(G297) );
  NAND2_X1 U666 ( .A1(n594), .A2(G559), .ZN(n595) );
  INV_X1 U667 ( .A(n920), .ZN(n635) );
  NAND2_X1 U668 ( .A1(n595), .A2(n635), .ZN(n596) );
  XNOR2_X1 U669 ( .A(n596), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U670 ( .A1(G559), .A2(n656), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n635), .A2(n597), .ZN(n598) );
  XNOR2_X1 U672 ( .A(n598), .B(KEYINPUT77), .ZN(n600) );
  NOR2_X1 U673 ( .A1(n923), .A2(G868), .ZN(n599) );
  NOR2_X1 U674 ( .A1(n600), .A2(n599), .ZN(G282) );
  NAND2_X1 U675 ( .A1(G99), .A2(n886), .ZN(n602) );
  NAND2_X1 U676 ( .A1(G111), .A2(n882), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U678 ( .A(KEYINPUT78), .B(n603), .ZN(n609) );
  BUF_X1 U679 ( .A(n604), .Z(n883) );
  NAND2_X1 U680 ( .A1(G123), .A2(n883), .ZN(n605) );
  XNOR2_X1 U681 ( .A(n605), .B(KEYINPUT18), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n887), .A2(G135), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n1004) );
  XNOR2_X1 U685 ( .A(G2096), .B(n1004), .ZN(n611) );
  INV_X1 U686 ( .A(G2100), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(G156) );
  NAND2_X1 U688 ( .A1(G49), .A2(n642), .ZN(n613) );
  NAND2_X1 U689 ( .A1(G74), .A2(G651), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U691 ( .A(KEYINPUT80), .B(n614), .Z(n619) );
  NAND2_X1 U692 ( .A1(G87), .A2(n615), .ZN(n616) );
  XNOR2_X1 U693 ( .A(KEYINPUT81), .B(n616), .ZN(n617) );
  NOR2_X1 U694 ( .A1(n637), .A2(n617), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(G288) );
  NAND2_X1 U696 ( .A1(G62), .A2(n637), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G75), .A2(n641), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U699 ( .A1(G88), .A2(n638), .ZN(n622) );
  XNOR2_X1 U700 ( .A(KEYINPUT83), .B(n622), .ZN(n623) );
  NOR2_X1 U701 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n642), .A2(G50), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n626), .A2(n625), .ZN(G303) );
  XOR2_X1 U704 ( .A(KEYINPUT2), .B(KEYINPUT82), .Z(n628) );
  NAND2_X1 U705 ( .A1(G73), .A2(n641), .ZN(n627) );
  XNOR2_X1 U706 ( .A(n628), .B(n627), .ZN(n632) );
  NAND2_X1 U707 ( .A1(G61), .A2(n637), .ZN(n630) );
  NAND2_X1 U708 ( .A1(G86), .A2(n638), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U710 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U711 ( .A1(n642), .A2(G48), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n634), .A2(n633), .ZN(G305) );
  NAND2_X1 U713 ( .A1(G559), .A2(n635), .ZN(n636) );
  XNOR2_X1 U714 ( .A(n636), .B(n923), .ZN(n834) );
  NAND2_X1 U715 ( .A1(G67), .A2(n637), .ZN(n640) );
  NAND2_X1 U716 ( .A1(G93), .A2(n638), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n640), .A2(n639), .ZN(n646) );
  NAND2_X1 U718 ( .A1(G80), .A2(n641), .ZN(n644) );
  NAND2_X1 U719 ( .A1(G55), .A2(n642), .ZN(n643) );
  NAND2_X1 U720 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U721 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U722 ( .A(KEYINPUT79), .B(n647), .ZN(n835) );
  XOR2_X1 U723 ( .A(n835), .B(G299), .Z(n648) );
  XNOR2_X1 U724 ( .A(n648), .B(G288), .ZN(n649) );
  XNOR2_X1 U725 ( .A(KEYINPUT19), .B(n649), .ZN(n651) );
  XNOR2_X1 U726 ( .A(G290), .B(KEYINPUT84), .ZN(n650) );
  XNOR2_X1 U727 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U728 ( .A(n652), .B(G303), .ZN(n653) );
  XNOR2_X1 U729 ( .A(n653), .B(G305), .ZN(n899) );
  XOR2_X1 U730 ( .A(n899), .B(KEYINPUT85), .Z(n654) );
  XNOR2_X1 U731 ( .A(n834), .B(n654), .ZN(n655) );
  NAND2_X1 U732 ( .A1(n655), .A2(G868), .ZN(n658) );
  NAND2_X1 U733 ( .A1(n656), .A2(n835), .ZN(n657) );
  NAND2_X1 U734 ( .A1(n658), .A2(n657), .ZN(G295) );
  NAND2_X1 U735 ( .A1(G2078), .A2(G2084), .ZN(n659) );
  XOR2_X1 U736 ( .A(KEYINPUT20), .B(n659), .Z(n660) );
  NAND2_X1 U737 ( .A1(G2090), .A2(n660), .ZN(n661) );
  XNOR2_X1 U738 ( .A(KEYINPUT21), .B(n661), .ZN(n662) );
  NAND2_X1 U739 ( .A1(n662), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U740 ( .A(KEYINPUT86), .B(G44), .ZN(n663) );
  XNOR2_X1 U741 ( .A(n663), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U742 ( .A1(G236), .A2(G237), .ZN(n664) );
  NAND2_X1 U743 ( .A1(G69), .A2(n664), .ZN(n665) );
  XNOR2_X1 U744 ( .A(KEYINPUT87), .B(n665), .ZN(n666) );
  NAND2_X1 U745 ( .A1(n666), .A2(G108), .ZN(n832) );
  NAND2_X1 U746 ( .A1(n832), .A2(G567), .ZN(n671) );
  NOR2_X1 U747 ( .A1(G220), .A2(G219), .ZN(n667) );
  XOR2_X1 U748 ( .A(KEYINPUT22), .B(n667), .Z(n668) );
  NOR2_X1 U749 ( .A1(G218), .A2(n668), .ZN(n669) );
  NAND2_X1 U750 ( .A1(G96), .A2(n669), .ZN(n833) );
  NAND2_X1 U751 ( .A1(n833), .A2(G2106), .ZN(n670) );
  NAND2_X1 U752 ( .A1(n671), .A2(n670), .ZN(n837) );
  NAND2_X1 U753 ( .A1(G661), .A2(G483), .ZN(n672) );
  NOR2_X1 U754 ( .A1(n837), .A2(n672), .ZN(n831) );
  NAND2_X1 U755 ( .A1(n831), .A2(G36), .ZN(G176) );
  NAND2_X1 U756 ( .A1(G102), .A2(n886), .ZN(n674) );
  NAND2_X1 U757 ( .A1(G138), .A2(n887), .ZN(n673) );
  NAND2_X1 U758 ( .A1(n674), .A2(n673), .ZN(n678) );
  NAND2_X1 U759 ( .A1(G114), .A2(n882), .ZN(n676) );
  NAND2_X1 U760 ( .A1(G126), .A2(n883), .ZN(n675) );
  NAND2_X1 U761 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U762 ( .A1(n678), .A2(n677), .ZN(G164) );
  INV_X1 U763 ( .A(G303), .ZN(G166) );
  NAND2_X1 U764 ( .A1(G160), .A2(G40), .ZN(n752) );
  XOR2_X1 U765 ( .A(KEYINPUT96), .B(n752), .Z(n679) );
  NOR2_X1 U766 ( .A1(G164), .A2(G1384), .ZN(n753) );
  NAND2_X2 U767 ( .A1(n679), .A2(n753), .ZN(n728) );
  INV_X2 U768 ( .A(n728), .ZN(n710) );
  NAND2_X1 U769 ( .A1(n710), .A2(G2072), .ZN(n680) );
  XOR2_X1 U770 ( .A(n680), .B(KEYINPUT27), .Z(n682) );
  NAND2_X1 U771 ( .A1(G1956), .A2(n728), .ZN(n681) );
  NAND2_X1 U772 ( .A1(n682), .A2(n681), .ZN(n685) );
  NAND2_X1 U773 ( .A1(n685), .A2(G299), .ZN(n683) );
  XNOR2_X1 U774 ( .A(n683), .B(KEYINPUT97), .ZN(n684) );
  XNOR2_X1 U775 ( .A(n684), .B(KEYINPUT28), .ZN(n708) );
  XNOR2_X1 U776 ( .A(n686), .B(KEYINPUT99), .ZN(n701) );
  XNOR2_X1 U777 ( .A(G1996), .B(KEYINPUT98), .ZN(n977) );
  NAND2_X1 U778 ( .A1(n977), .A2(n710), .ZN(n688) );
  XNOR2_X1 U779 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n694) );
  INV_X1 U780 ( .A(n694), .ZN(n687) );
  NAND2_X1 U781 ( .A1(n688), .A2(n687), .ZN(n692) );
  INV_X1 U782 ( .A(G1341), .ZN(n922) );
  NAND2_X1 U783 ( .A1(G1348), .A2(n920), .ZN(n689) );
  NAND2_X1 U784 ( .A1(n922), .A2(n689), .ZN(n690) );
  NAND2_X1 U785 ( .A1(n728), .A2(n690), .ZN(n691) );
  NAND2_X1 U786 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U787 ( .A1(n923), .A2(n693), .ZN(n699) );
  NAND2_X1 U788 ( .A1(n920), .A2(G2067), .ZN(n696) );
  NAND2_X1 U789 ( .A1(n694), .A2(n977), .ZN(n695) );
  NAND2_X1 U790 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U791 ( .A1(n697), .A2(n710), .ZN(n698) );
  NAND2_X1 U792 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U793 ( .A1(n701), .A2(n700), .ZN(n706) );
  NAND2_X1 U794 ( .A1(G1348), .A2(n728), .ZN(n703) );
  NAND2_X1 U795 ( .A1(G2067), .A2(n710), .ZN(n702) );
  NAND2_X1 U796 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U797 ( .A1(n920), .A2(n704), .ZN(n705) );
  NOR2_X1 U798 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U799 ( .A(G2078), .B(KEYINPUT25), .Z(n983) );
  NOR2_X1 U800 ( .A1(n983), .A2(n728), .ZN(n712) );
  NOR2_X1 U801 ( .A1(n710), .A2(G1961), .ZN(n711) );
  NOR2_X1 U802 ( .A1(n712), .A2(n711), .ZN(n719) );
  NOR2_X1 U803 ( .A1(n719), .A2(G301), .ZN(n713) );
  NOR2_X1 U804 ( .A1(n516), .A2(n713), .ZN(n724) );
  NOR2_X1 U805 ( .A1(G1966), .A2(n802), .ZN(n739) );
  NOR2_X1 U806 ( .A1(G2084), .A2(n728), .ZN(n738) );
  NOR2_X1 U807 ( .A1(n739), .A2(n738), .ZN(n714) );
  NAND2_X1 U808 ( .A1(G8), .A2(n714), .ZN(n716) );
  NOR2_X1 U809 ( .A1(G168), .A2(n717), .ZN(n718) );
  XNOR2_X1 U810 ( .A(n718), .B(KEYINPUT101), .ZN(n721) );
  NAND2_X1 U811 ( .A1(n719), .A2(G301), .ZN(n720) );
  NAND2_X1 U812 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U813 ( .A(KEYINPUT31), .B(n722), .Z(n723) );
  NOR2_X1 U814 ( .A1(n724), .A2(n723), .ZN(n726) );
  INV_X1 U815 ( .A(KEYINPUT102), .ZN(n725) );
  XNOR2_X1 U816 ( .A(n726), .B(n725), .ZN(n740) );
  NAND2_X1 U817 ( .A1(n740), .A2(G286), .ZN(n735) );
  INV_X1 U818 ( .A(G8), .ZN(n733) );
  NOR2_X1 U819 ( .A1(G1971), .A2(n802), .ZN(n727) );
  XNOR2_X1 U820 ( .A(KEYINPUT103), .B(n727), .ZN(n731) );
  NOR2_X1 U821 ( .A1(G2090), .A2(n728), .ZN(n729) );
  NOR2_X1 U822 ( .A1(G166), .A2(n729), .ZN(n730) );
  NAND2_X1 U823 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U824 ( .A1(n735), .A2(n734), .ZN(n737) );
  XNOR2_X1 U825 ( .A(n737), .B(n736), .ZN(n745) );
  NAND2_X1 U826 ( .A1(G8), .A2(n738), .ZN(n743) );
  INV_X1 U827 ( .A(n740), .ZN(n741) );
  NOR2_X1 U828 ( .A1(n739), .A2(n741), .ZN(n742) );
  NAND2_X1 U829 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U830 ( .A1(n745), .A2(n744), .ZN(n799) );
  NOR2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n932) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n746) );
  NOR2_X1 U833 ( .A1(n932), .A2(n746), .ZN(n748) );
  INV_X1 U834 ( .A(KEYINPUT33), .ZN(n747) );
  AND2_X1 U835 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U836 ( .A1(n799), .A2(n749), .ZN(n791) );
  NAND2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n929) );
  INV_X1 U838 ( .A(n929), .ZN(n750) );
  NOR2_X1 U839 ( .A1(KEYINPUT33), .A2(n518), .ZN(n789) );
  NAND2_X1 U840 ( .A1(n932), .A2(KEYINPUT33), .ZN(n751) );
  OR2_X1 U841 ( .A1(n751), .A2(n802), .ZN(n787) );
  XOR2_X1 U842 ( .A(G1981), .B(G305), .Z(n942) );
  NOR2_X1 U843 ( .A1(n753), .A2(n752), .ZN(n823) );
  NAND2_X1 U844 ( .A1(G104), .A2(n886), .ZN(n755) );
  NAND2_X1 U845 ( .A1(G140), .A2(n887), .ZN(n754) );
  NAND2_X1 U846 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U847 ( .A(KEYINPUT34), .B(n756), .ZN(n762) );
  NAND2_X1 U848 ( .A1(G116), .A2(n882), .ZN(n758) );
  NAND2_X1 U849 ( .A1(G128), .A2(n883), .ZN(n757) );
  NAND2_X1 U850 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U851 ( .A(KEYINPUT88), .B(n759), .Z(n760) );
  XNOR2_X1 U852 ( .A(KEYINPUT35), .B(n760), .ZN(n761) );
  NOR2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U854 ( .A(KEYINPUT36), .B(n763), .ZN(n876) );
  XNOR2_X1 U855 ( .A(KEYINPUT37), .B(G2067), .ZN(n820) );
  OR2_X1 U856 ( .A1(n876), .A2(n820), .ZN(n764) );
  XNOR2_X1 U857 ( .A(n764), .B(KEYINPUT89), .ZN(n1017) );
  NAND2_X1 U858 ( .A1(n823), .A2(n1017), .ZN(n818) );
  NAND2_X1 U859 ( .A1(G95), .A2(n886), .ZN(n766) );
  NAND2_X1 U860 ( .A1(G131), .A2(n887), .ZN(n765) );
  NAND2_X1 U861 ( .A1(n766), .A2(n765), .ZN(n767) );
  XOR2_X1 U862 ( .A(KEYINPUT90), .B(n767), .Z(n771) );
  NAND2_X1 U863 ( .A1(G107), .A2(n882), .ZN(n769) );
  NAND2_X1 U864 ( .A1(G119), .A2(n883), .ZN(n768) );
  AND2_X1 U865 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U866 ( .A1(n771), .A2(n770), .ZN(n879) );
  NAND2_X1 U867 ( .A1(G1991), .A2(n879), .ZN(n772) );
  XNOR2_X1 U868 ( .A(KEYINPUT91), .B(n772), .ZN(n784) );
  NAND2_X1 U869 ( .A1(G117), .A2(n882), .ZN(n774) );
  NAND2_X1 U870 ( .A1(G129), .A2(n883), .ZN(n773) );
  NAND2_X1 U871 ( .A1(n774), .A2(n773), .ZN(n777) );
  NAND2_X1 U872 ( .A1(n886), .A2(G105), .ZN(n775) );
  XOR2_X1 U873 ( .A(KEYINPUT38), .B(n775), .Z(n776) );
  NOR2_X1 U874 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U875 ( .A(KEYINPUT92), .B(n778), .ZN(n781) );
  NAND2_X1 U876 ( .A1(n887), .A2(G141), .ZN(n779) );
  XOR2_X1 U877 ( .A(KEYINPUT93), .B(n779), .Z(n780) );
  NAND2_X1 U878 ( .A1(n781), .A2(n780), .ZN(n875) );
  NAND2_X1 U879 ( .A1(G1996), .A2(n875), .ZN(n782) );
  XOR2_X1 U880 ( .A(KEYINPUT94), .B(n782), .Z(n783) );
  NOR2_X1 U881 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U882 ( .A(KEYINPUT95), .B(n785), .ZN(n1016) );
  NAND2_X1 U883 ( .A1(n823), .A2(n1016), .ZN(n812) );
  AND2_X1 U884 ( .A1(n818), .A2(n812), .ZN(n801) );
  AND2_X1 U885 ( .A1(n942), .A2(n801), .ZN(n786) );
  NAND2_X1 U886 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U887 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U888 ( .A1(n791), .A2(n790), .ZN(n808) );
  NOR2_X1 U889 ( .A1(G2090), .A2(G303), .ZN(n792) );
  XNOR2_X1 U890 ( .A(n792), .B(KEYINPUT104), .ZN(n793) );
  NAND2_X1 U891 ( .A1(n793), .A2(G8), .ZN(n797) );
  NOR2_X1 U892 ( .A1(G1981), .A2(G305), .ZN(n794) );
  XOR2_X1 U893 ( .A(n794), .B(KEYINPUT24), .Z(n795) );
  NOR2_X1 U894 ( .A1(n802), .A2(n795), .ZN(n796) );
  NAND2_X1 U895 ( .A1(n801), .A2(n796), .ZN(n800) );
  NAND2_X1 U896 ( .A1(n799), .A2(n798), .ZN(n806) );
  INV_X1 U897 ( .A(n800), .ZN(n804) );
  AND2_X1 U898 ( .A1(n802), .A2(n801), .ZN(n803) );
  OR2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U901 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U902 ( .A(G1986), .B(G290), .ZN(n925) );
  NAND2_X1 U903 ( .A1(n517), .A2(n810), .ZN(n811) );
  XNOR2_X1 U904 ( .A(n811), .B(KEYINPUT106), .ZN(n825) );
  NOR2_X1 U905 ( .A1(G1996), .A2(n875), .ZN(n1012) );
  INV_X1 U906 ( .A(n812), .ZN(n815) );
  NOR2_X1 U907 ( .A1(G1991), .A2(n879), .ZN(n1008) );
  NOR2_X1 U908 ( .A1(G1986), .A2(G290), .ZN(n813) );
  NOR2_X1 U909 ( .A1(n1008), .A2(n813), .ZN(n814) );
  NOR2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U911 ( .A1(n1012), .A2(n816), .ZN(n817) );
  XNOR2_X1 U912 ( .A(n817), .B(KEYINPUT39), .ZN(n819) );
  NAND2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n820), .A2(n876), .ZN(n1009) );
  NAND2_X1 U915 ( .A1(n821), .A2(n1009), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n825), .A2(n824), .ZN(n827) );
  XOR2_X1 U918 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n826) );
  XNOR2_X1 U919 ( .A(n827), .B(n826), .ZN(G329) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n828), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U922 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n831), .A2(n830), .ZN(G188) );
  INV_X1 U926 ( .A(G108), .ZN(G238) );
  INV_X1 U927 ( .A(G96), .ZN(G221) );
  NOR2_X1 U928 ( .A1(n833), .A2(n832), .ZN(G325) );
  INV_X1 U929 ( .A(G325), .ZN(G261) );
  NOR2_X1 U930 ( .A1(n834), .A2(G860), .ZN(n836) );
  XOR2_X1 U931 ( .A(n836), .B(n835), .Z(G145) );
  INV_X1 U932 ( .A(n837), .ZN(G319) );
  XOR2_X1 U933 ( .A(G2096), .B(KEYINPUT43), .Z(n839) );
  XNOR2_X1 U934 ( .A(G2072), .B(KEYINPUT108), .ZN(n838) );
  XNOR2_X1 U935 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U936 ( .A(n840), .B(G2678), .Z(n842) );
  XNOR2_X1 U937 ( .A(G2067), .B(G2090), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U939 ( .A(KEYINPUT42), .B(G2100), .Z(n844) );
  XNOR2_X1 U940 ( .A(G2078), .B(G2084), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U942 ( .A(n846), .B(n845), .ZN(G227) );
  XOR2_X1 U943 ( .A(G1976), .B(G1981), .Z(n848) );
  XNOR2_X1 U944 ( .A(G1986), .B(G1971), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U946 ( .A(G1961), .B(G1966), .Z(n850) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1991), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U949 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U950 ( .A(KEYINPUT109), .B(G2474), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n854), .B(n853), .ZN(n856) );
  XOR2_X1 U952 ( .A(G1956), .B(KEYINPUT41), .Z(n855) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(G229) );
  NAND2_X1 U954 ( .A1(n887), .A2(G136), .ZN(n863) );
  NAND2_X1 U955 ( .A1(G100), .A2(n886), .ZN(n858) );
  NAND2_X1 U956 ( .A1(G112), .A2(n882), .ZN(n857) );
  NAND2_X1 U957 ( .A1(n858), .A2(n857), .ZN(n861) );
  NAND2_X1 U958 ( .A1(n883), .A2(G124), .ZN(n859) );
  XOR2_X1 U959 ( .A(KEYINPUT44), .B(n859), .Z(n860) );
  NOR2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n862) );
  NAND2_X1 U961 ( .A1(n863), .A2(n862), .ZN(n864) );
  XOR2_X1 U962 ( .A(KEYINPUT110), .B(n864), .Z(G162) );
  XOR2_X1 U963 ( .A(KEYINPUT48), .B(KEYINPUT111), .Z(n873) );
  NAND2_X1 U964 ( .A1(G103), .A2(n886), .ZN(n866) );
  NAND2_X1 U965 ( .A1(G139), .A2(n887), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n871) );
  NAND2_X1 U967 ( .A1(G115), .A2(n882), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G127), .A2(n883), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U970 ( .A(KEYINPUT47), .B(n869), .Z(n870) );
  NOR2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n999) );
  XNOR2_X1 U972 ( .A(n999), .B(KEYINPUT46), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U974 ( .A(n875), .B(n874), .ZN(n878) );
  XOR2_X1 U975 ( .A(G164), .B(n876), .Z(n877) );
  XNOR2_X1 U976 ( .A(n878), .B(n877), .ZN(n880) );
  XNOR2_X1 U977 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U978 ( .A(n881), .B(G162), .ZN(n894) );
  NAND2_X1 U979 ( .A1(G118), .A2(n882), .ZN(n885) );
  NAND2_X1 U980 ( .A1(G130), .A2(n883), .ZN(n884) );
  NAND2_X1 U981 ( .A1(n885), .A2(n884), .ZN(n892) );
  NAND2_X1 U982 ( .A1(G106), .A2(n886), .ZN(n889) );
  NAND2_X1 U983 ( .A1(G142), .A2(n887), .ZN(n888) );
  NAND2_X1 U984 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U985 ( .A(KEYINPUT45), .B(n890), .Z(n891) );
  NOR2_X1 U986 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U987 ( .A(n894), .B(n893), .Z(n896) );
  XNOR2_X1 U988 ( .A(G160), .B(n1004), .ZN(n895) );
  XNOR2_X1 U989 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U990 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U991 ( .A(G171), .B(n920), .ZN(n898) );
  XNOR2_X1 U992 ( .A(KEYINPUT112), .B(n898), .ZN(n901) );
  XNOR2_X1 U993 ( .A(n923), .B(n899), .ZN(n900) );
  XNOR2_X1 U994 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U995 ( .A(n902), .B(G286), .ZN(n903) );
  NOR2_X1 U996 ( .A1(G37), .A2(n903), .ZN(G397) );
  XOR2_X1 U997 ( .A(G2451), .B(G2430), .Z(n905) );
  XNOR2_X1 U998 ( .A(G2438), .B(G2443), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n905), .B(n904), .ZN(n911) );
  XOR2_X1 U1000 ( .A(G2435), .B(G2454), .Z(n907) );
  XNOR2_X1 U1001 ( .A(G1341), .B(G1348), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n909) );
  XOR2_X1 U1003 ( .A(G2446), .B(G2427), .Z(n908) );
  XNOR2_X1 U1004 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1005 ( .A(n911), .B(n910), .Z(n912) );
  NAND2_X1 U1006 ( .A1(G14), .A2(n912), .ZN(n919) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n919), .ZN(n916) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n913) );
  XOR2_X1 U1009 ( .A(KEYINPUT49), .B(n913), .Z(n914) );
  XNOR2_X1 U1010 ( .A(n914), .B(KEYINPUT113), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1013 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G69), .ZN(G235) );
  INV_X1 U1016 ( .A(n919), .ZN(G401) );
  XNOR2_X1 U1017 ( .A(G16), .B(KEYINPUT56), .ZN(n950) );
  XNOR2_X1 U1018 ( .A(n920), .B(G1348), .ZN(n921) );
  XNOR2_X1 U1019 ( .A(n921), .B(KEYINPUT119), .ZN(n940) );
  XNOR2_X1 U1020 ( .A(n923), .B(n922), .ZN(n927) );
  XNOR2_X1 U1021 ( .A(G1961), .B(G301), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n938) );
  XNOR2_X1 U1024 ( .A(G299), .B(G1956), .ZN(n935) );
  XNOR2_X1 U1025 ( .A(G166), .B(G1971), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(n928), .B(KEYINPUT120), .ZN(n930) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1029 ( .A(KEYINPUT121), .B(n933), .ZN(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1031 ( .A(KEYINPUT122), .B(n936), .Z(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n947) );
  XNOR2_X1 U1034 ( .A(KEYINPUT118), .B(KEYINPUT57), .ZN(n945) );
  XOR2_X1 U1035 ( .A(G1966), .B(G168), .Z(n941) );
  XNOR2_X1 U1036 ( .A(KEYINPUT117), .B(n941), .ZN(n943) );
  NAND2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1038 ( .A(n945), .B(n944), .Z(n946) );
  NOR2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(KEYINPUT123), .B(n948), .ZN(n949) );
  NAND2_X1 U1041 ( .A1(n950), .A2(n949), .ZN(n1027) );
  XOR2_X1 U1042 ( .A(G16), .B(KEYINPUT124), .Z(n975) );
  XNOR2_X1 U1043 ( .A(G1966), .B(G21), .ZN(n952) );
  XNOR2_X1 U1044 ( .A(G5), .B(G1961), .ZN(n951) );
  NOR2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n965) );
  XNOR2_X1 U1046 ( .A(KEYINPUT127), .B(KEYINPUT60), .ZN(n963) );
  XNOR2_X1 U1047 ( .A(KEYINPUT59), .B(KEYINPUT126), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(n953), .B(G4), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(G1348), .B(n954), .ZN(n961) );
  XNOR2_X1 U1050 ( .A(G1956), .B(G20), .ZN(n959) );
  XNOR2_X1 U1051 ( .A(G1341), .B(G19), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(G1981), .B(G6), .ZN(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(KEYINPUT125), .B(n957), .ZN(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(n963), .B(n962), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n972) );
  XNOR2_X1 U1059 ( .A(G1971), .B(G22), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(G23), .B(G1976), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n969) );
  XOR2_X1 U1062 ( .A(G1986), .B(G24), .Z(n968) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(KEYINPUT58), .B(n970), .ZN(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(n973), .B(KEYINPUT61), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1068 ( .A1(G11), .A2(n976), .ZN(n1025) );
  XNOR2_X1 U1069 ( .A(G1991), .B(G25), .ZN(n988) );
  XNOR2_X1 U1070 ( .A(n977), .B(G32), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(G26), .B(G2067), .ZN(n978) );
  NOR2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n982) );
  XOR2_X1 U1073 ( .A(G2072), .B(KEYINPUT114), .Z(n980) );
  XNOR2_X1 U1074 ( .A(G33), .B(n980), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n985) );
  XNOR2_X1 U1076 ( .A(G27), .B(n983), .ZN(n984) );
  NOR2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(KEYINPUT115), .B(n986), .ZN(n987) );
  NOR2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1080 ( .A1(G28), .A2(n989), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(KEYINPUT53), .B(n990), .ZN(n994) );
  XOR2_X1 U1082 ( .A(G34), .B(KEYINPUT116), .Z(n992) );
  XNOR2_X1 U1083 ( .A(G2084), .B(KEYINPUT54), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(n992), .B(n991), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(G35), .B(G2090), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(G29), .A2(n997), .ZN(n998) );
  XNOR2_X1 U1089 ( .A(n998), .B(KEYINPUT55), .ZN(n1023) );
  XOR2_X1 U1090 ( .A(G2072), .B(n999), .Z(n1001) );
  XOR2_X1 U1091 ( .A(G164), .B(G2078), .Z(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(KEYINPUT50), .B(n1002), .ZN(n1006) );
  XOR2_X1 U1094 ( .A(G160), .B(G2084), .Z(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1015) );
  XOR2_X1 U1099 ( .A(G2090), .B(G162), .Z(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(n1013), .B(KEYINPUT51), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1019) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(KEYINPUT52), .B(n1020), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(G29), .A2(n1021), .ZN(n1022) );
  NAND2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1109 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1028), .Z(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

