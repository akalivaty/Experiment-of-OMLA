//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1292, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1360, new_n1361, new_n1362, new_n1363;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  XOR2_X1   g0008(.A(KEYINPUT66), .B(G244), .Z(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G77), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT65), .B(G68), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n210), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(KEYINPUT67), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n214), .A2(KEYINPUT67), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n208), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n208), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT0), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n206), .A2(KEYINPUT64), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT64), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G20), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  AND2_X1   g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n202), .A2(G50), .ZN(new_n232));
  OAI22_X1  g0032(.A1(new_n224), .A2(new_n225), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(new_n225), .B2(new_n224), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n221), .A2(new_n222), .A3(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT68), .Z(G361));
  XOR2_X1   g0036(.A(G238), .B(G244), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT69), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G13), .ZN(new_n253));
  NOR3_X1   g0053(.A1(new_n253), .A2(new_n206), .A3(G1), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G50), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G1), .A2(G13), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(G1), .B2(new_n206), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n256), .B1(new_n262), .B2(G50), .ZN(new_n263));
  OAI21_X1  g0063(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G150), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT64), .B(G20), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G33), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT8), .B(G58), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n264), .B(new_n266), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n259), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT9), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT9), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT10), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(G222), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G77), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n283), .A2(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(G223), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n285), .B1(new_n286), .B2(new_n283), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT71), .ZN(new_n290));
  AND2_X1   g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n290), .B1(new_n291), .B2(new_n258), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n230), .A2(KEYINPUT71), .A3(new_n293), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n230), .A2(new_n293), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G226), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT70), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n205), .B(KEYINPUT70), .C1(G41), .C2(G45), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n302), .A2(new_n297), .A3(G274), .A4(new_n303), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n296), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G190), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT74), .B(G200), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n277), .A2(new_n278), .A3(new_n309), .A4(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n274), .A2(new_n312), .A3(new_n276), .ZN(new_n314));
  OAI21_X1  g0114(.A(KEYINPUT10), .B1(new_n314), .B2(new_n308), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n306), .ZN(new_n317));
  INV_X1    g0117(.A(G179), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(KEYINPUT72), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n319), .A2(KEYINPUT72), .ZN(new_n321));
  OAI221_X1 g0121(.A(new_n272), .B1(G169), .B2(new_n317), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n299), .A2(new_n209), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n304), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n283), .A2(G232), .A3(new_n284), .ZN(new_n325));
  INV_X1    g0125(.A(G107), .ZN(new_n326));
  OAI221_X1 g0126(.A(new_n325), .B1(new_n326), .B2(new_n283), .C1(new_n287), .C2(new_n212), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n324), .B1(new_n327), .B2(new_n295), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n318), .ZN(new_n329));
  INV_X1    g0129(.A(new_n269), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n330), .A2(new_n265), .B1(new_n229), .B2(G77), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT15), .B(G87), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(G33), .A3(new_n267), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n260), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT73), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n255), .B2(G77), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n254), .A2(KEYINPUT73), .A3(new_n286), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n337), .B(new_n338), .C1(new_n261), .C2(new_n286), .ZN(new_n339));
  OAI221_X1 g0139(.A(new_n329), .B1(G169), .B2(new_n328), .C1(new_n335), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n328), .A2(G190), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n339), .A2(new_n335), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n341), .B(new_n342), .C1(new_n310), .C2(new_n328), .ZN(new_n343));
  AND4_X1   g0143(.A1(new_n316), .A2(new_n322), .A3(new_n340), .A4(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G68), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(new_n261), .B2(KEYINPUT12), .ZN(new_n346));
  AND3_X1   g0146(.A1(new_n213), .A2(new_n254), .A3(KEYINPUT12), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n254), .A2(KEYINPUT12), .ZN(new_n348));
  OR3_X1    g0148(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n213), .A2(G20), .B1(G50), .B2(new_n265), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n286), .B2(new_n268), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT75), .B(KEYINPUT11), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n259), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n259), .ZN(new_n354));
  INV_X1    g0154(.A(new_n352), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n349), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  AND2_X1   g0157(.A1(KEYINPUT3), .A2(G33), .ZN(new_n358));
  NOR2_X1   g0158(.A1(KEYINPUT3), .A2(G33), .ZN(new_n359));
  OAI211_X1 g0159(.A(G232), .B(G1698), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  OAI211_X1 g0160(.A(G226), .B(new_n284), .C1(new_n358), .C2(new_n359), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G33), .A2(G97), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n363), .A2(new_n295), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n297), .A2(G238), .A3(new_n298), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n304), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(KEYINPUT13), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n366), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n363), .A2(new_n295), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT13), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G200), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n367), .A2(G190), .A3(new_n371), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n357), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n364), .A2(KEYINPUT13), .A3(new_n366), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n370), .B1(new_n368), .B2(new_n369), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n378), .A2(KEYINPUT77), .A3(G179), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n367), .A2(G179), .A3(new_n371), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT77), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G169), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(KEYINPUT76), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT14), .B1(new_n372), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT14), .ZN(new_n386));
  INV_X1    g0186(.A(new_n384), .ZN(new_n387));
  AOI211_X1 g0187(.A(new_n386), .B(new_n387), .C1(new_n367), .C2(new_n371), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n379), .B(new_n382), .C1(new_n385), .C2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n357), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n375), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n261), .A2(new_n330), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n255), .A2(new_n269), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n358), .A2(new_n359), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT7), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(new_n267), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n281), .A2(new_n206), .A3(new_n282), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT7), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n399), .A3(G68), .ZN(new_n400));
  INV_X1    g0200(.A(G58), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n202), .B1(new_n213), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G20), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n265), .A2(G159), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n400), .A2(new_n403), .A3(KEYINPUT16), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n259), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT7), .B1(new_n229), .B2(new_n283), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n345), .A2(KEYINPUT65), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT65), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(G68), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n407), .B(new_n411), .C1(KEYINPUT7), .C2(new_n398), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n402), .A2(G20), .B1(G159), .B2(new_n265), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT16), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n394), .B1(new_n406), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(G200), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n292), .A2(new_n294), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G87), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n288), .A2(new_n284), .ZN(new_n420));
  INV_X1    g0220(.A(G226), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G1698), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n420), .B(new_n422), .C1(new_n358), .C2(new_n359), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n418), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n297), .A2(G232), .A3(new_n298), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n304), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n417), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n423), .A2(new_n419), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n295), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n429), .A2(new_n307), .A3(new_n304), .A4(new_n425), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n427), .A2(new_n430), .A3(KEYINPUT78), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n424), .A2(new_n426), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT78), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(new_n307), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n416), .A2(new_n435), .A3(KEYINPUT17), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n420), .A2(new_n422), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n437), .A2(new_n283), .B1(G33), .B2(G87), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n304), .B(new_n425), .C1(new_n438), .C2(new_n418), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G169), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n318), .B2(new_n439), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n415), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT18), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT16), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n396), .B1(new_n395), .B2(new_n267), .ZN(new_n445));
  NOR4_X1   g0245(.A1(new_n358), .A2(new_n359), .A3(KEYINPUT7), .A4(G20), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n445), .A2(new_n446), .A3(new_n213), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n201), .B1(new_n411), .B2(G58), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n404), .B1(new_n448), .B2(new_n206), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n444), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(new_n259), .A3(new_n405), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n451), .A2(new_n431), .A3(new_n394), .A4(new_n434), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT17), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT18), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n415), .A2(new_n455), .A3(new_n441), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n436), .A2(new_n443), .A3(new_n454), .A4(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n344), .A2(new_n391), .A3(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n333), .A2(new_n255), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n226), .A2(new_n228), .A3(G33), .A4(G97), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT19), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT82), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n461), .A2(KEYINPUT82), .A3(new_n462), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n283), .A2(new_n267), .A3(G68), .ZN(new_n467));
  INV_X1    g0267(.A(G87), .ZN(new_n468));
  INV_X1    g0268(.A(G97), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(new_n469), .A3(new_n326), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n362), .A2(new_n462), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n470), .B1(new_n229), .B2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n465), .A2(new_n466), .A3(new_n467), .A4(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n460), .B1(new_n473), .B2(new_n259), .ZN(new_n474));
  OAI211_X1 g0274(.A(G238), .B(new_n284), .C1(new_n358), .C2(new_n359), .ZN(new_n475));
  OAI211_X1 g0275(.A(G244), .B(G1698), .C1(new_n358), .C2(new_n359), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G116), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n295), .ZN(new_n479));
  INV_X1    g0279(.A(G45), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(G1), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G274), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT81), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(KEYINPUT81), .A3(G274), .ZN(new_n485));
  INV_X1    g0285(.A(G250), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n484), .A2(new_n485), .B1(new_n297), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n479), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n311), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n205), .A2(G33), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n255), .A2(new_n260), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G87), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n474), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT83), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n489), .B2(new_n307), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n479), .A2(new_n488), .A3(KEYINPUT83), .A4(G190), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n492), .A2(new_n332), .ZN(new_n500));
  AOI211_X1 g0300(.A(new_n460), .B(new_n500), .C1(new_n473), .C2(new_n259), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n479), .A2(new_n318), .A3(new_n488), .ZN(new_n502));
  INV_X1    g0302(.A(new_n489), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(G169), .ZN(new_n504));
  OAI22_X1  g0304(.A1(new_n495), .A2(new_n499), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT84), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n500), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n474), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(G169), .B1(new_n479), .B2(new_n488), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n510), .B1(new_n318), .B2(new_n503), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n512), .B(KEYINPUT84), .C1(new_n495), .C2(new_n499), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(KEYINPUT23), .A2(G107), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n227), .A2(G20), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n206), .A2(KEYINPUT64), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g0319(.A1(KEYINPUT23), .A2(G107), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT23), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n477), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n520), .B1(new_n522), .B2(new_n206), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n226), .B(new_n228), .C1(new_n358), .C2(new_n359), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT22), .B1(new_n525), .B2(new_n468), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT22), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n283), .A2(new_n267), .A3(new_n527), .A4(G87), .ZN(new_n528));
  AOI211_X1 g0328(.A(KEYINPUT24), .B(new_n524), .C1(new_n526), .C2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT24), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n526), .A2(new_n528), .ZN(new_n531));
  INV_X1    g0331(.A(new_n524), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n259), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT85), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT85), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n536), .B(new_n259), .C1(new_n529), .C2(new_n533), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(G250), .B(new_n284), .C1(new_n358), .C2(new_n359), .ZN(new_n539));
  OAI211_X1 g0339(.A(G257), .B(G1698), .C1(new_n358), .C2(new_n359), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G294), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n295), .ZN(new_n543));
  XNOR2_X1  g0343(.A(KEYINPUT5), .B(G41), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n544), .A2(new_n481), .B1(new_n230), .B2(new_n293), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G264), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n544), .A2(new_n297), .A3(G274), .A4(new_n481), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n543), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(KEYINPUT86), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT86), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n542), .A2(new_n295), .B1(new_n545), .B2(G264), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n550), .B1(new_n551), .B2(new_n547), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n307), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT87), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n548), .A2(new_n554), .A3(new_n417), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n548), .A2(new_n417), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT87), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n553), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT25), .B1(new_n254), .B2(new_n326), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n254), .A2(KEYINPUT25), .A3(new_n326), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n493), .A2(G107), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n538), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n562), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n535), .B2(new_n537), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n548), .A2(new_n318), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n549), .A2(new_n552), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(G169), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n283), .A2(G264), .A3(G1698), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n283), .A2(G257), .A3(new_n284), .ZN(new_n572));
  INV_X1    g0372(.A(G303), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n571), .B(new_n572), .C1(new_n573), .C2(new_n283), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n295), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n297), .A2(G274), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n544), .A2(new_n481), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n576), .A2(new_n578), .B1(new_n545), .B2(G270), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n383), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n493), .A2(G116), .ZN(new_n581));
  INV_X1    g0381(.A(G116), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n254), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n257), .A2(new_n258), .B1(G20), .B2(new_n582), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G33), .A2(G283), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n469), .B2(G33), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n584), .B1(new_n229), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT20), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n587), .A2(new_n588), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n581), .B(new_n583), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n580), .A2(new_n591), .A3(KEYINPUT21), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT21), .B1(new_n580), .B2(new_n591), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n589), .A2(new_n590), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n583), .B1(new_n492), .B2(new_n582), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n575), .A2(new_n579), .A3(G179), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR3_X1   g0398(.A1(new_n592), .A2(new_n593), .A3(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(G244), .B(new_n284), .C1(new_n358), .C2(new_n359), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT4), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n283), .A2(KEYINPUT4), .A3(G244), .A4(new_n284), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n283), .A2(G250), .A3(G1698), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .A4(new_n585), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n295), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n577), .A2(G257), .A3(new_n297), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n547), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n383), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n608), .B1(new_n295), .B2(new_n605), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n318), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n445), .A2(new_n446), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n614), .A2(G107), .B1(G77), .B2(new_n265), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT80), .ZN(new_n616));
  AND2_X1   g0416(.A1(KEYINPUT79), .A2(KEYINPUT6), .ZN(new_n617));
  NOR2_X1   g0417(.A1(KEYINPUT79), .A2(KEYINPUT6), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n469), .A2(G107), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n616), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OR2_X1    g0421(.A1(KEYINPUT79), .A2(KEYINPUT6), .ZN(new_n622));
  NAND2_X1  g0422(.A1(KEYINPUT79), .A2(KEYINPUT6), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n616), .A2(new_n622), .A3(new_n620), .A4(new_n623), .ZN(new_n624));
  OAI22_X1  g0424(.A1(new_n621), .A2(new_n624), .B1(new_n469), .B2(G107), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n622), .A2(new_n620), .A3(new_n623), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT80), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n619), .A2(new_n616), .A3(new_n620), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n469), .A2(G107), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n625), .A2(new_n229), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n260), .B1(new_n615), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n254), .A2(new_n469), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n492), .B2(new_n469), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n611), .B(new_n613), .C1(new_n632), .C2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n615), .A2(new_n631), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n634), .B1(new_n636), .B2(new_n259), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n606), .A2(new_n307), .A3(new_n609), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(G200), .B2(new_n612), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n575), .A2(new_n579), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n591), .B1(G200), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(new_n307), .B2(new_n641), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n599), .A2(new_n635), .A3(new_n640), .A4(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  AND4_X1   g0445(.A1(new_n459), .A2(new_n515), .A3(new_n570), .A4(new_n645), .ZN(G372));
  NAND2_X1  g0446(.A1(new_n443), .A2(new_n456), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n389), .A2(new_n390), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n375), .B2(new_n340), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n436), .A2(new_n454), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n647), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT88), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n316), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n313), .A2(KEYINPUT88), .A3(new_n315), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n322), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT89), .ZN(new_n657));
  INV_X1    g0457(.A(new_n635), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n507), .A2(new_n513), .A3(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(KEYINPUT26), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n503), .A2(G190), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n661), .A2(new_n474), .A3(new_n490), .A4(new_n494), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n512), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(new_n658), .A3(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n640), .A2(new_n635), .A3(new_n662), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n538), .A2(new_n558), .A3(new_n562), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n580), .A2(new_n591), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT21), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n580), .A2(new_n591), .A3(KEYINPUT21), .ZN(new_n672));
  INV_X1    g0472(.A(new_n597), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n591), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n671), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n531), .A2(new_n532), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT24), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n531), .A2(new_n530), .A3(new_n532), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n536), .B1(new_n679), .B2(new_n259), .ZN(new_n680));
  INV_X1    g0480(.A(new_n537), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n562), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n549), .A2(new_n552), .ZN(new_n683));
  OAI22_X1  g0483(.A1(new_n683), .A2(new_n383), .B1(new_n318), .B2(new_n548), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n675), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n512), .B(new_n665), .C1(new_n668), .C2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n459), .B1(new_n660), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n657), .A2(new_n687), .ZN(G369));
  INV_X1    g0488(.A(KEYINPUT90), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n682), .A2(new_n684), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n667), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n229), .A2(new_n253), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n205), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT27), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n692), .A2(new_n695), .A3(new_n205), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n694), .A2(G213), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n682), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n689), .B1(new_n691), .B2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n690), .A2(new_n700), .A3(KEYINPUT90), .A4(new_n667), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n699), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n690), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(KEYINPUT91), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT91), .ZN(new_n710));
  AOI211_X1 g0510(.A(new_n710), .B(new_n706), .C1(new_n702), .C2(new_n703), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n705), .A2(new_n596), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n675), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n599), .A2(new_n643), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n715), .B1(new_n716), .B2(new_n714), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G330), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n713), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT92), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n675), .A2(new_n705), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT93), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(new_n708), .B2(new_n711), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n690), .A2(new_n699), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n721), .A2(new_n728), .ZN(G399));
  INV_X1    g0529(.A(new_n223), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G41), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n470), .A2(G116), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n732), .A2(G1), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(new_n232), .B2(new_n732), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT28), .ZN(new_n736));
  INV_X1    g0536(.A(G330), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT94), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT30), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n551), .A2(new_n479), .A3(new_n488), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n612), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n739), .B1(new_n741), .B2(new_n597), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n673), .A2(KEYINPUT30), .A3(new_n612), .A4(new_n740), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n503), .A2(G179), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n744), .A2(new_n548), .A3(new_n610), .A4(new_n641), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT31), .B1(new_n746), .B2(new_n699), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n738), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n746), .A2(new_n699), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT31), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n752), .A2(KEYINPUT94), .A3(new_n753), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n570), .A2(new_n645), .A3(new_n515), .A4(new_n705), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n737), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n705), .B1(new_n686), .B2(new_n660), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT29), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n666), .A2(new_n667), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n690), .A2(new_n599), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n761), .A2(new_n762), .B1(new_n509), .B2(new_n511), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n659), .A2(KEYINPUT95), .A3(new_n664), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n663), .A2(KEYINPUT26), .A3(new_n658), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(KEYINPUT95), .B1(new_n659), .B2(new_n664), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n763), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n768), .A2(KEYINPUT29), .A3(new_n705), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n757), .B1(new_n760), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n736), .B1(new_n770), .B2(G1), .ZN(G364));
  AOI21_X1  g0571(.A(new_n258), .B1(G20), .B2(new_n383), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n310), .A2(G179), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n267), .A2(G190), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT96), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G107), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n206), .A2(new_n307), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n774), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n778), .B(new_n283), .C1(new_n468), .C2(new_n780), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT97), .Z(new_n782));
  NOR2_X1   g0582(.A1(G179), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n775), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G159), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT32), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n267), .A2(new_n318), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n307), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G200), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G50), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n789), .A2(G190), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n417), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n788), .B1(new_n792), .B2(new_n286), .C1(new_n793), .C2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n267), .B1(G190), .B2(new_n783), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n798), .A2(KEYINPUT98), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(KEYINPUT98), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G97), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n794), .A2(G200), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n790), .A2(new_n417), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G58), .A2(new_n804), .B1(new_n805), .B2(G68), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n803), .B(new_n806), .C1(new_n787), .C2(new_n786), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n782), .A2(new_n797), .A3(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(KEYINPUT100), .B(KEYINPUT33), .ZN(new_n809));
  INV_X1    g0609(.A(G317), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n809), .B(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n805), .ZN(new_n812));
  INV_X1    g0612(.A(new_n804), .ZN(new_n813));
  INV_X1    g0613(.A(G322), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n811), .A2(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT101), .Z(new_n816));
  INV_X1    g0616(.A(new_n784), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n283), .B1(new_n817), .B2(G329), .ZN(new_n818));
  INV_X1    g0618(.A(G326), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n796), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G294), .ZN(new_n821));
  INV_X1    g0621(.A(G311), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n801), .A2(new_n821), .B1(new_n792), .B2(new_n822), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n780), .B(KEYINPUT99), .Z(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n777), .ZN(new_n826));
  INV_X1    g0626(.A(G283), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n825), .A2(new_n573), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR4_X1   g0628(.A1(new_n816), .A2(new_n820), .A3(new_n823), .A4(new_n828), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n808), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n773), .B1(new_n830), .B2(KEYINPUT102), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(KEYINPUT102), .B2(new_n830), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n205), .B1(new_n692), .B2(G45), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(new_n731), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n248), .A2(G45), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n730), .A2(new_n283), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n837), .B(new_n838), .C1(G45), .C2(new_n232), .ZN(new_n839));
  INV_X1    g0639(.A(G355), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n223), .A2(new_n283), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n839), .B1(G116), .B2(new_n223), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(G13), .A2(G33), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n844), .A2(G20), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n845), .A2(new_n772), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n836), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n845), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n832), .B(new_n847), .C1(new_n717), .C2(new_n848), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT103), .Z(new_n850));
  NOR2_X1   g0650(.A1(new_n717), .A2(G330), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n719), .A2(new_n851), .A3(new_n835), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(G396));
  OAI21_X1  g0654(.A(new_n343), .B1(new_n342), .B2(new_n705), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n340), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n340), .A2(new_n699), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n758), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n858), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n705), .B(new_n860), .C1(new_n686), .C2(new_n660), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n757), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n732), .B2(new_n833), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n757), .A2(new_n859), .A3(new_n861), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n772), .A2(new_n843), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n836), .B1(new_n286), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n283), .B1(new_n817), .B2(G311), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n803), .B(new_n868), .C1(new_n825), .C2(new_n326), .ZN(new_n869));
  AOI22_X1  g0669(.A1(G116), .A2(new_n791), .B1(new_n795), .B2(G303), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n870), .B1(new_n827), .B2(new_n812), .C1(new_n821), .C2(new_n813), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n826), .A2(new_n468), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n869), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI22_X1  g0673(.A1(G137), .A2(new_n795), .B1(new_n805), .B2(G150), .ZN(new_n874));
  INV_X1    g0674(.A(G143), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n874), .B1(new_n875), .B2(new_n813), .C1(new_n785), .C2(new_n792), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT34), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n825), .A2(new_n793), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n826), .A2(new_n345), .ZN(new_n880));
  INV_X1    g0680(.A(G132), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n283), .B1(new_n881), .B2(new_n784), .C1(new_n801), .C2(new_n401), .ZN(new_n882));
  NOR4_X1   g0682(.A1(new_n878), .A2(new_n879), .A3(new_n880), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n876), .A2(new_n877), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n873), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI221_X1 g0685(.A(new_n867), .B1(new_n860), .B2(new_n844), .C1(new_n885), .C2(new_n773), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n865), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(G384));
  NOR2_X1   g0688(.A1(new_n692), .A2(new_n205), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n747), .A2(new_n748), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n756), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT40), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n390), .A2(new_n699), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n386), .B1(new_n378), .B2(new_n387), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n372), .A2(KEYINPUT14), .A3(new_n384), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n380), .B(KEYINPUT77), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n893), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n391), .B2(new_n893), .ZN(new_n899));
  AOI211_X1 g0699(.A(new_n858), .B(new_n899), .C1(new_n756), .C2(new_n890), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT38), .ZN(new_n901));
  INV_X1    g0701(.A(new_n697), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n457), .A2(new_n415), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT37), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n440), .B(new_n697), .C1(new_n318), .C2(new_n439), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n415), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n905), .B1(new_n907), .B2(new_n452), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n907), .A2(new_n452), .A3(new_n905), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n909), .A2(KEYINPUT105), .A3(new_n910), .ZN(new_n911));
  AOI211_X1 g0711(.A(KEYINPUT105), .B(new_n905), .C1(new_n907), .C2(new_n452), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n901), .B1(new_n904), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT16), .B1(new_n413), .B2(new_n400), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n394), .B1(new_n406), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n457), .A2(new_n902), .A3(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n416), .A2(new_n435), .B1(new_n917), .B2(new_n906), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n910), .B1(new_n919), .B2(new_n905), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n918), .A2(KEYINPUT38), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n915), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n892), .B1(new_n900), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n899), .ZN(new_n924));
  NOR4_X1   g0724(.A1(new_n691), .A2(new_n644), .A3(new_n514), .A4(new_n699), .ZN(new_n925));
  INV_X1    g0725(.A(new_n890), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n860), .B(new_n924), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n921), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT38), .B1(new_n918), .B2(new_n920), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n892), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n459), .B(new_n891), .C1(new_n923), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n910), .A2(KEYINPUT105), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n933), .A2(new_n908), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n934), .A2(new_n912), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT38), .B1(new_n935), .B2(new_n903), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n936), .A2(new_n928), .ZN(new_n937));
  OAI21_X1  g0737(.A(KEYINPUT40), .B1(new_n937), .B2(new_n927), .ZN(new_n938));
  INV_X1    g0738(.A(new_n929), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n921), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n900), .A2(new_n892), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n459), .A2(new_n891), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n938), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n932), .A2(G330), .A3(new_n943), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT106), .Z(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n769), .A2(new_n459), .A3(new_n760), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n657), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT39), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n936), .B2(new_n928), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n648), .A2(new_n699), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n939), .A2(KEYINPUT39), .A3(new_n921), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n861), .A2(new_n857), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(new_n924), .A3(new_n940), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n647), .A2(new_n697), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n948), .B(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n889), .B1(new_n946), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n946), .B2(new_n958), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n231), .A2(new_n582), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n625), .A2(new_n630), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT35), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n963), .B2(new_n962), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT36), .Z(new_n966));
  AOI211_X1 g0766(.A(new_n286), .B(new_n232), .C1(new_n411), .C2(G58), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT104), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n967), .A2(new_n968), .B1(new_n793), .B2(G68), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n968), .B2(new_n967), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n970), .A2(G1), .A3(new_n253), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n960), .A2(new_n966), .A3(new_n971), .ZN(G367));
  OAI22_X1  g0772(.A1(new_n793), .A2(new_n792), .B1(new_n796), .B2(new_n875), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(G159), .B2(new_n805), .ZN(new_n974));
  XOR2_X1   g0774(.A(KEYINPUT111), .B(G137), .Z(new_n975));
  OAI22_X1  g0775(.A1(new_n776), .A2(new_n286), .B1(new_n784), .B2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n780), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n395), .B(new_n976), .C1(G58), .C2(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n801), .A2(new_n345), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(G150), .B2(new_n804), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n974), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT46), .B1(new_n977), .B2(G116), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT46), .ZN(new_n983));
  NOR3_X1   g0783(.A1(new_n825), .A2(new_n983), .A3(new_n582), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n982), .B(new_n984), .C1(G294), .C2(new_n805), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(KEYINPUT110), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n573), .A2(new_n813), .B1(new_n796), .B2(new_n822), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n801), .A2(new_n326), .B1(new_n792), .B2(new_n827), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n395), .B1(new_n784), .B2(new_n810), .C1(new_n469), .C2(new_n776), .ZN(new_n989));
  NOR3_X1   g0789(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n986), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n985), .A2(KEYINPUT110), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n981), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT47), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n772), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n474), .A2(new_n494), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n699), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n663), .A2(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n997), .A2(new_n512), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n998), .A2(new_n845), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n838), .A2(new_n243), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n846), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n730), .B2(new_n333), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n836), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n995), .A2(new_n1000), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n713), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n723), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n719), .A2(KEYINPUT109), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1007), .A2(new_n725), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n713), .A2(new_n724), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n723), .B1(new_n709), .B2(new_n712), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n718), .B(KEYINPUT109), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1009), .B(new_n770), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n640), .B(new_n635), .C1(new_n637), .C2(new_n705), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n658), .A2(new_n699), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n725), .A2(new_n727), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT45), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n725), .A2(KEYINPUT45), .A3(new_n727), .A4(new_n1017), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n725), .A2(new_n727), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1017), .ZN(new_n1024));
  AOI21_X1  g0824(.A(KEYINPUT44), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT44), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1026), .B(new_n1017), .C1(new_n725), .C2(new_n727), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1022), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n721), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1014), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n721), .B(new_n1022), .C1(new_n1025), .C2(new_n1027), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n770), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n731), .B(KEYINPUT41), .Z(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n834), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n721), .A2(new_n1024), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n998), .A2(new_n999), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT107), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1039), .A2(KEYINPUT43), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(KEYINPUT43), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1038), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(KEYINPUT43), .B2(new_n1038), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n635), .B1(new_n690), .B2(new_n1015), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n705), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1011), .A2(new_n1017), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1046), .B1(new_n1047), .B2(KEYINPUT42), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT108), .ZN(new_n1049));
  OR3_X1    g0849(.A1(new_n725), .A2(KEYINPUT42), .A3(new_n1024), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1049), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1043), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1053), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1055), .A2(new_n1051), .A3(new_n1042), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1037), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1054), .A2(new_n1056), .A3(new_n1037), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1005), .B1(new_n1036), .B2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT112), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(G387));
  INV_X1    g0863(.A(new_n770), .ZN(new_n1064));
  AND3_X1   g0864(.A1(new_n1007), .A2(new_n725), .A3(new_n1008), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1013), .B1(new_n1007), .B2(new_n725), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1064), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1067), .A2(new_n731), .A3(new_n1014), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n395), .B1(new_n784), .B2(new_n819), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G303), .A2(new_n791), .B1(new_n804), .B2(G317), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n822), .B2(new_n812), .C1(new_n814), .C2(new_n796), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT48), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n802), .A2(G283), .B1(G294), .B2(new_n977), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1076), .B(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n776), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1069), .B(new_n1078), .C1(G116), .C2(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G68), .A2(new_n791), .B1(new_n795), .B2(G159), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n793), .B2(new_n813), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n780), .A2(new_n286), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n395), .B(new_n1083), .C1(G150), .C2(new_n817), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n802), .A2(new_n333), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(new_n269), .C2(new_n812), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1082), .B(new_n1086), .C1(G97), .C2(new_n777), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n772), .B1(new_n1080), .B2(new_n1087), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n841), .A2(new_n733), .B1(G107), .B2(new_n223), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n240), .A2(new_n480), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n733), .ZN(new_n1091));
  AOI211_X1 g0891(.A(G45), .B(new_n1091), .C1(G68), .C2(G77), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n269), .A2(G50), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT50), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n730), .B(new_n283), .C1(new_n1092), .C2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1089), .B1(new_n1090), .B2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1088), .B(new_n835), .C1(new_n1002), .C2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n1006), .B2(new_n845), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1098), .B1(new_n1099), .B2(new_n834), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1068), .A2(new_n1100), .ZN(G393));
  NAND2_X1  g0901(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT114), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n1031), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1028), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1105), .A2(KEYINPUT114), .A3(new_n721), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT115), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1104), .A2(KEYINPUT115), .A3(new_n1106), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n834), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1104), .A2(new_n1014), .A3(new_n1106), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n732), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1024), .A2(new_n845), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n846), .B1(new_n469), .B2(new_n223), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n838), .B2(new_n251), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n283), .B1(new_n780), .B2(new_n213), .C1(new_n875), .C2(new_n784), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n872), .A2(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n802), .A2(G77), .B1(G50), .B2(new_n805), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1118), .B(new_n1119), .C1(new_n269), .C2(new_n792), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(G150), .A2(new_n795), .B1(new_n804), .B2(G159), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT51), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G311), .A2(new_n804), .B1(new_n795), .B2(G317), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT52), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n802), .A2(G116), .B1(G303), .B2(new_n805), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n791), .A2(G294), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n395), .B1(new_n780), .B2(new_n827), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(G322), .B2(new_n817), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1125), .A2(new_n778), .A3(new_n1126), .A4(new_n1128), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n1120), .A2(new_n1122), .B1(new_n1124), .B2(new_n1129), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n836), .B(new_n1116), .C1(new_n1130), .C2(new_n772), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1112), .A2(new_n1113), .B1(new_n1114), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1111), .A2(new_n1132), .ZN(G390));
  AOI21_X1  g0933(.A(new_n899), .B1(new_n861), .B2(new_n857), .ZN(new_n1134));
  AOI21_X1  g0934(.A(KEYINPUT39), .B1(new_n915), .B2(new_n921), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n928), .A2(new_n929), .A3(new_n949), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n1134), .A2(new_n951), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n768), .A2(new_n705), .A3(new_n856), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n899), .B1(new_n1138), .B2(new_n857), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n951), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n922), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1137), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT116), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n891), .A2(G330), .A3(new_n860), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1144), .A2(new_n899), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1142), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n757), .A2(new_n860), .A3(new_n924), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1137), .B(new_n1147), .C1(new_n1139), .C2(new_n1141), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1143), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1146), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n924), .B1(new_n757), .B2(new_n860), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n954), .B1(new_n1151), .B2(new_n1145), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1144), .A2(new_n899), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1147), .A2(new_n857), .A3(new_n1138), .A4(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n459), .A2(G330), .A3(new_n891), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n657), .A2(new_n947), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n732), .B1(new_n1150), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n1150), .B2(new_n1159), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n866), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n395), .B1(new_n821), .B2(new_n784), .C1(new_n801), .C2(new_n286), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1163), .B(new_n880), .C1(G87), .C2(new_n824), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n582), .A2(new_n813), .B1(new_n796), .B2(new_n827), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n469), .A2(new_n792), .B1(new_n812), .B2(new_n326), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n395), .B1(new_n817), .B2(G125), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n793), .B2(new_n776), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT117), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT53), .ZN(new_n1171));
  INV_X1    g0971(.A(G150), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n780), .A2(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1171), .A2(new_n1173), .B1(new_n795), .B2(G128), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n881), .B2(new_n813), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT54), .B(G143), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n801), .A2(new_n785), .B1(new_n792), .B2(new_n1176), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n812), .A2(new_n975), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1175), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1164), .A2(new_n1167), .B1(new_n1170), .B2(new_n1179), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n835), .B1(new_n330), .B2(new_n1162), .C1(new_n1180), .C2(new_n773), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT118), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1182), .B1(new_n1184), .B2(new_n843), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1138), .A2(new_n857), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1141), .B1(new_n1186), .B2(new_n924), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n954), .A2(new_n924), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1188), .A2(new_n1140), .B1(new_n950), .B2(new_n952), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1145), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1190), .A2(KEYINPUT116), .A3(new_n1148), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1142), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1185), .B1(new_n1193), .B2(new_n834), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1161), .A2(new_n1194), .ZN(G378));
  AND3_X1   g0995(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n1196));
  OAI21_X1  g0996(.A(G330), .B1(new_n923), .B2(new_n931), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n938), .A2(new_n941), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n957), .A2(new_n1199), .A3(G330), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n653), .A2(new_n322), .A3(new_n654), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(KEYINPUT120), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT120), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n653), .A2(new_n1203), .A3(new_n322), .A4(new_n654), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  XOR2_X1   g1005(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n273), .A2(new_n697), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1206), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1202), .A2(new_n1204), .A3(new_n1209), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1207), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1208), .B1(new_n1207), .B2(new_n1210), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1198), .A2(new_n1200), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1213), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n834), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n836), .B1(new_n793), .B2(new_n866), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n802), .A2(G150), .B1(G132), .B2(new_n805), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1176), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n804), .A2(G128), .B1(new_n977), .B2(new_n1220), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G125), .A2(new_n795), .B1(new_n791), .B2(G137), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1219), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1079), .A2(G159), .ZN(new_n1226));
  AOI211_X1 g1026(.A(G33), .B(G41), .C1(new_n817), .C2(G124), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1079), .A2(G58), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n827), .B2(new_n784), .ZN(new_n1230));
  OR3_X1    g1030(.A1(new_n1083), .A2(G41), .A3(new_n283), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1230), .B(new_n979), .C1(KEYINPUT119), .C2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(KEYINPUT119), .B2(new_n1231), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n795), .A2(G116), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n805), .A2(G97), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n326), .B2(new_n813), .C1(new_n332), .C2(new_n792), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1233), .A2(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1238), .A2(KEYINPUT58), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(KEYINPUT58), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n793), .B1(new_n358), .B2(G41), .ZN(new_n1241));
  AND4_X1   g1041(.A1(new_n1228), .A2(new_n1239), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1218), .B1(new_n773), .B2(new_n1242), .C1(new_n1213), .C2(new_n844), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1217), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1158), .B1(new_n1150), .B2(new_n1159), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT57), .B1(new_n1246), .B2(new_n1216), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n731), .B1(new_n1247), .B2(KEYINPUT122), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT121), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1246), .A2(new_n1249), .A3(KEYINPUT57), .A4(new_n1216), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1159), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1216), .B(KEYINPUT57), .C1(new_n1251), .C2(new_n1157), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT121), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT57), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1159), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1157), .B1(new_n1193), .B2(new_n1255), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1257));
  OAI211_X1 g1057(.A(KEYINPUT122), .B(new_n1254), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1250), .A2(new_n1253), .A3(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1245), .B1(new_n1248), .B2(new_n1259), .ZN(G375));
  OAI22_X1  g1060(.A1(new_n825), .A2(new_n469), .B1(new_n826), .B2(new_n286), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1085), .B(new_n395), .C1(new_n573), .C2(new_n784), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n1261), .B(new_n1262), .C1(G283), .C2(new_n804), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(G116), .A2(new_n805), .B1(new_n795), .B2(G294), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n326), .B2(new_n792), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(KEYINPUT124), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1229), .A2(new_n283), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(KEYINPUT125), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n805), .A2(new_n1220), .B1(new_n817), .B2(G128), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n825), .B2(new_n785), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n881), .A2(new_n796), .B1(new_n813), .B2(new_n975), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n801), .A2(new_n793), .B1(new_n792), .B2(new_n1172), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1263), .A2(new_n1266), .B1(new_n1268), .B2(new_n1273), .ZN(new_n1274));
  OAI221_X1 g1074(.A(new_n835), .B1(G68), .B2(new_n1162), .C1(new_n1274), .C2(new_n773), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(new_n843), .B2(new_n899), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n833), .B(KEYINPUT123), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1276), .B1(new_n1155), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1159), .A2(new_n1035), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1278), .B1(new_n1279), .B2(new_n1280), .ZN(G381));
  INV_X1    g1081(.A(G378), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1250), .A2(new_n1253), .A3(new_n1258), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1254), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT122), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n732), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1244), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1068), .A2(new_n1100), .A3(new_n853), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n887), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(G390), .A2(G381), .A3(new_n1289), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1062), .A2(new_n1282), .A3(new_n1287), .A4(new_n1290), .ZN(G407));
  NAND2_X1  g1091(.A1(new_n1287), .A2(new_n1282), .ZN(new_n1292));
  OAI211_X1 g1092(.A(G407), .B(G213), .C1(G343), .C2(new_n1292), .ZN(G409));
  INV_X1    g1093(.A(new_n1005), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n833), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1059), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1297), .A2(new_n1057), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1294), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT112), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n853), .B1(new_n1068), .B2(new_n1100), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1300), .B1(new_n1288), .B2(new_n1301), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1111), .A2(new_n1132), .A3(new_n1302), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1288), .A2(new_n1301), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1304), .B1(new_n1111), .B2(new_n1132), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1299), .B1(new_n1303), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1304), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(G390), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1111), .A2(new_n1132), .A3(new_n1302), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1308), .A2(new_n1061), .A3(new_n1309), .ZN(new_n1310));
  AND2_X1   g1110(.A1(new_n1306), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(G375), .A2(G378), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1216), .A2(new_n1277), .ZN(new_n1314));
  AND2_X1   g1114(.A1(new_n1314), .A2(new_n1243), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1246), .A2(new_n1035), .A3(new_n1216), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1161), .A2(new_n1315), .A3(new_n1316), .A4(new_n1194), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n698), .A2(G213), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT60), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT126), .ZN(new_n1323));
  OR3_X1    g1123(.A1(new_n1322), .A2(new_n1280), .A3(new_n1323), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1323), .B1(new_n1322), .B2(new_n1280), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n732), .B1(new_n1280), .B2(KEYINPUT60), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1324), .A2(new_n1325), .A3(new_n1326), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1327), .A2(G384), .A3(new_n1278), .ZN(new_n1328));
  AOI21_X1  g1128(.A(G384), .B1(new_n1327), .B2(new_n1278), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1313), .A2(new_n1320), .A3(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(KEYINPUT62), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1319), .B1(G375), .B2(G378), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT62), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1333), .A2(new_n1334), .A3(new_n1330), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1332), .A2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n698), .A2(G213), .A3(G2897), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1338), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1327), .A2(new_n1278), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(new_n887), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1327), .A2(G384), .A3(new_n1278), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1341), .A2(new_n1342), .A3(new_n1337), .ZN(new_n1343));
  AND2_X1   g1143(.A1(new_n1339), .A2(new_n1343), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1286), .A2(new_n1258), .A3(new_n1253), .A4(new_n1250), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1282), .B1(new_n1345), .B2(new_n1245), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1344), .B1(new_n1346), .B2(new_n1319), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT61), .ZN(new_n1348));
  AOI21_X1  g1148(.A(KEYINPUT127), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1312), .B1(new_n1336), .B2(new_n1349), .ZN(new_n1350));
  AND4_X1   g1150(.A1(KEYINPUT63), .A2(new_n1313), .A3(new_n1320), .A4(new_n1330), .ZN(new_n1351));
  AOI21_X1  g1151(.A(KEYINPUT63), .B1(new_n1333), .B2(new_n1330), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1311), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1353));
  AOI21_X1  g1153(.A(KEYINPUT127), .B1(new_n1306), .B2(new_n1310), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1339), .A2(new_n1343), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1348), .B1(new_n1333), .B2(new_n1355), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1354), .A2(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1353), .A2(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1350), .A2(new_n1358), .ZN(G405));
  NAND2_X1  g1159(.A1(new_n1292), .A2(new_n1313), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1360), .A2(new_n1330), .ZN(new_n1361));
  OAI211_X1 g1161(.A(new_n1292), .B(new_n1313), .C1(new_n1329), .C2(new_n1328), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  XNOR2_X1  g1163(.A(new_n1363), .B(new_n1311), .ZN(G402));
endmodule


