//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1248, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G77), .ZN(new_n211));
  INV_X1    g0011(.A(G244), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT65), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n213), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n218), .B1(new_n214), .B2(new_n217), .ZN(new_n219));
  INV_X1    g0019(.A(G1), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT66), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT64), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n221), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n223), .A2(G13), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT0), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n231), .B(new_n234), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n226), .A2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  OR2_X1    g0051(.A1(KEYINPUT67), .A2(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  NAND2_X1  g0053(.A1(KEYINPUT67), .A2(G41), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n220), .A2(G274), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n229), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n253), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n220), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G226), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n258), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n272), .A2(G223), .B1(G77), .B2(new_n270), .ZN(new_n273));
  INV_X1    g0073(.A(G222), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n260), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n271), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n273), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT68), .ZN(new_n282));
  XNOR2_X1  g0082(.A(new_n281), .B(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n267), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(G179), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT69), .ZN(new_n288));
  INV_X1    g0088(.A(G58), .ZN(new_n289));
  OR3_X1    g0089(.A1(new_n289), .A2(KEYINPUT69), .A3(KEYINPUT8), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n288), .A2(new_n221), .A3(G33), .A4(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n292), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n259), .B1(new_n222), .B2(G33), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G13), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n297), .A2(new_n221), .A3(G1), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G50), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n295), .B1(G1), .B2(new_n221), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(new_n202), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n296), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n284), .A2(G169), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n286), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT9), .B1(new_n296), .B2(new_n303), .ZN(new_n307));
  INV_X1    g0107(.A(new_n303), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n308), .B(new_n309), .C1(new_n295), .C2(new_n294), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n285), .A2(G200), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT71), .B1(new_n284), .B2(G190), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT10), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT10), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n311), .A2(new_n312), .A3(new_n316), .A4(new_n313), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n306), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n272), .A2(G238), .B1(G107), .B2(new_n270), .ZN(new_n319));
  INV_X1    g0119(.A(G232), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(new_n279), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n283), .ZN(new_n322));
  INV_X1    g0122(.A(new_n265), .ZN(new_n323));
  AOI22_X1  g0123(.A1(G244), .A2(new_n323), .B1(new_n255), .B2(new_n257), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G179), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n302), .A2(new_n211), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT70), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n328), .B(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n298), .A2(new_n211), .ZN(new_n331));
  INV_X1    g0131(.A(new_n287), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n332), .A2(new_n292), .B1(G20), .B2(G77), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n221), .A2(G33), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT15), .B(G87), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n295), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n330), .A2(new_n331), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n322), .A2(new_n324), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n327), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n339), .B1(G200), .B2(new_n340), .ZN(new_n344));
  INV_X1    g0144(.A(G190), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n344), .B1(new_n345), .B2(new_n340), .ZN(new_n346));
  AND3_X1   g0146(.A1(new_n318), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n289), .A2(new_n209), .ZN(new_n348));
  OAI21_X1  g0148(.A(G20), .B1(new_n348), .B2(new_n201), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n292), .A2(G159), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AND2_X1   g0151(.A1(KEYINPUT75), .A2(G33), .ZN(new_n352));
  NOR2_X1   g0152(.A1(KEYINPUT75), .A2(G33), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT3), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n354), .A2(new_n221), .A3(new_n276), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n355), .A2(KEYINPUT7), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT7), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n354), .A2(new_n357), .A3(new_n221), .A4(new_n276), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G68), .ZN(new_n359));
  OAI211_X1 g0159(.A(KEYINPUT16), .B(new_n351), .C1(new_n356), .C2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT76), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n355), .A2(KEYINPUT7), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n363), .A2(G68), .A3(new_n358), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n364), .A2(KEYINPUT76), .A3(KEYINPUT16), .A4(new_n351), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT75), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n260), .ZN(new_n368));
  NAND2_X1  g0168(.A1(KEYINPUT75), .A2(G33), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(new_n275), .A3(new_n369), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n277), .A2(KEYINPUT7), .A3(new_n221), .ZN(new_n371));
  AOI21_X1  g0171(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n276), .A2(new_n372), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n370), .A2(new_n371), .B1(new_n373), .B2(new_n357), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n351), .B1(new_n374), .B2(new_n209), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT16), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n366), .A2(new_n337), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n258), .B1(new_n265), .B2(new_n320), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n275), .B1(new_n368), .B2(new_n369), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n380), .A2(new_n269), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n266), .A2(G1698), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(G223), .B2(G1698), .ZN(new_n383));
  INV_X1    g0183(.A(G87), .ZN(new_n384));
  OAI22_X1  g0184(.A1(new_n381), .A2(new_n383), .B1(new_n260), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n379), .B1(new_n385), .B2(new_n283), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G190), .ZN(new_n387));
  INV_X1    g0187(.A(G200), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n387), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n288), .A2(new_n290), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n302), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n299), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n378), .A2(new_n390), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT17), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n377), .A2(new_n337), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n362), .B2(new_n365), .ZN(new_n400));
  INV_X1    g0200(.A(new_n395), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n400), .A2(new_n389), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT17), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n386), .A2(new_n341), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n386), .A2(G179), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n400), .B2(new_n401), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT18), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n406), .B(new_n409), .C1(new_n400), .C2(new_n401), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n398), .A2(new_n403), .A3(new_n408), .A4(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n292), .A2(G50), .B1(G20), .B2(new_n209), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n211), .B2(new_n334), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n337), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT11), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n299), .A2(KEYINPUT12), .A3(G68), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT12), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n298), .B2(new_n209), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n419), .A2(new_n421), .B1(new_n302), .B2(new_n209), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n415), .A2(new_n416), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n418), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT14), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n278), .A2(G226), .A3(new_n271), .ZN(new_n427));
  INV_X1    g0227(.A(G97), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT72), .B1(new_n260), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT72), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(G33), .A3(G97), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n278), .A2(G1698), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n427), .B(new_n432), .C1(new_n433), .C2(new_n320), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n283), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n258), .B1(new_n265), .B2(new_n210), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT13), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n435), .A2(KEYINPUT73), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n436), .B1(new_n283), .B2(new_n434), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n439), .B1(new_n440), .B2(new_n438), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT73), .B1(new_n440), .B2(new_n438), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n426), .B(G169), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n438), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT74), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OR2_X1    g0246(.A1(new_n440), .A2(new_n438), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n440), .A2(KEYINPUT74), .A3(new_n438), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n446), .A2(new_n447), .A3(G179), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n443), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT73), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n452), .A2(new_n447), .A3(new_n439), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n426), .B1(new_n453), .B2(G169), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n425), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(G200), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n446), .A2(new_n447), .A3(G190), .A4(new_n448), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n456), .A2(new_n424), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n347), .A2(new_n412), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT78), .ZN(new_n462));
  INV_X1    g0262(.A(G107), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n374), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n277), .A2(new_n221), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n357), .B1(new_n465), .B2(new_n269), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n372), .A2(KEYINPUT7), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n469), .A2(KEYINPUT78), .A3(G107), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT77), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT6), .ZN(new_n472));
  AND2_X1   g0272(.A1(G97), .A2(G107), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(new_n205), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n463), .A2(KEYINPUT6), .A3(G97), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n221), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n292), .A2(G77), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n471), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n463), .A2(KEYINPUT6), .A3(G97), .ZN(new_n480));
  XNOR2_X1  g0280(.A(G97), .B(G107), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n480), .B1(new_n481), .B2(new_n472), .ZN(new_n482));
  OAI211_X1 g0282(.A(KEYINPUT77), .B(new_n477), .C1(new_n482), .C2(new_n221), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n464), .A2(new_n470), .A3(new_n479), .A4(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n337), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n299), .A2(G97), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n220), .A2(G33), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n295), .A2(new_n299), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n486), .B1(new_n489), .B2(G97), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT80), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(new_n261), .A3(KEYINPUT5), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(new_n220), .A3(G45), .ZN(new_n493));
  NAND2_X1  g0293(.A1(KEYINPUT67), .A2(KEYINPUT80), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n252), .A2(new_n254), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT5), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G274), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n495), .A2(new_n496), .ZN(new_n499));
  OAI211_X1 g0299(.A(G257), .B(new_n262), .C1(new_n499), .C2(new_n493), .ZN(new_n500));
  AND2_X1   g0300(.A1(KEYINPUT4), .A2(G244), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n271), .B(new_n501), .C1(new_n268), .C2(new_n269), .ZN(new_n502));
  OAI211_X1 g0302(.A(G250), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G283), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(G244), .B(new_n271), .C1(new_n380), .C2(new_n269), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT4), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n283), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n498), .B(new_n500), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n485), .A2(new_n490), .B1(new_n510), .B2(new_n341), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT79), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n508), .B2(new_n509), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n212), .B1(new_n354), .B2(new_n276), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT4), .B1(new_n514), .B2(new_n271), .ZN(new_n515));
  OAI211_X1 g0315(.A(KEYINPUT79), .B(new_n283), .C1(new_n515), .C2(new_n505), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n500), .A2(new_n498), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n326), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n511), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n388), .B1(new_n517), .B2(new_n518), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT81), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n485), .A2(new_n490), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n518), .B(G190), .C1(new_n509), .C2(new_n508), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n523), .A2(new_n524), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n485), .A3(new_n490), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT81), .B1(new_n528), .B2(new_n522), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n521), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(G116), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n368), .B2(new_n369), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n221), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n463), .A2(G20), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT23), .ZN(new_n535));
  XNOR2_X1  g0335(.A(new_n534), .B(new_n535), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n354), .A2(new_n276), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n538), .A2(KEYINPUT22), .A3(new_n221), .A4(G87), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT22), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n221), .A2(G87), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n540), .B1(new_n270), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n537), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n543), .A2(KEYINPUT24), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n543), .A2(KEYINPUT24), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n337), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(G1698), .B1(new_n354), .B2(new_n276), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G250), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n538), .A2(G257), .A3(G1698), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n368), .A2(new_n369), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G294), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n283), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n497), .A2(new_n281), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G264), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n498), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G200), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n298), .A2(KEYINPUT25), .A3(new_n463), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT25), .B1(new_n298), .B2(new_n463), .ZN(new_n559));
  OAI22_X1  g0359(.A1(new_n488), .A2(new_n463), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n553), .A2(G190), .A3(new_n498), .A4(new_n555), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n546), .A2(new_n557), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n335), .A2(new_n298), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT19), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n429), .B2(new_n431), .ZN(new_n566));
  OAI22_X1  g0366(.A1(new_n566), .A2(G20), .B1(G87), .B2(new_n206), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n538), .A2(new_n221), .A3(G68), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n565), .B1(new_n334), .B2(new_n428), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n564), .B1(new_n570), .B2(new_n337), .ZN(new_n571));
  XNOR2_X1  g0371(.A(new_n335), .B(KEYINPUT83), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n571), .B1(new_n488), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(G244), .B(G1698), .C1(new_n380), .C2(new_n269), .ZN(new_n574));
  OAI211_X1 g0374(.A(G238), .B(new_n271), .C1(new_n380), .C2(new_n269), .ZN(new_n575));
  INV_X1    g0375(.A(new_n532), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n283), .ZN(new_n578));
  OAI21_X1  g0378(.A(G250), .B1(new_n253), .B2(G1), .ZN(new_n579));
  OAI22_X1  g0379(.A1(new_n281), .A2(new_n579), .B1(new_n253), .B2(new_n256), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT82), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI221_X1 g0382(.A(KEYINPUT82), .B1(new_n253), .B2(new_n256), .C1(new_n281), .C2(new_n579), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n341), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n577), .A2(new_n283), .B1(new_n582), .B2(new_n583), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n326), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n573), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n578), .A2(G190), .A3(new_n584), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT84), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT84), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n587), .A2(new_n592), .A3(G190), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n532), .B1(new_n547), .B2(G238), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n509), .B1(new_n594), .B2(new_n574), .ZN(new_n595));
  INV_X1    g0395(.A(new_n584), .ZN(new_n596));
  OAI21_X1  g0396(.A(G200), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n488), .A2(new_n384), .ZN(new_n598));
  AOI211_X1 g0398(.A(new_n564), .B(new_n598), .C1(new_n570), .C2(new_n337), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n591), .A2(new_n593), .A3(new_n597), .A4(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n563), .A2(new_n589), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n530), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(G264), .A2(G1698), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT85), .B1(new_n381), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT85), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n538), .A2(new_n605), .A3(G264), .A4(G1698), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n538), .A2(G257), .A3(new_n271), .ZN(new_n608));
  XOR2_X1   g0408(.A(KEYINPUT86), .B(G303), .Z(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n270), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n509), .B1(new_n607), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n554), .A2(G270), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n498), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G190), .ZN(new_n616));
  OAI21_X1  g0416(.A(G200), .B1(new_n612), .B2(new_n614), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n504), .B(new_n221), .C1(G33), .C2(new_n428), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT20), .ZN(new_n619));
  AOI22_X1  g0419(.A1(KEYINPUT87), .A2(new_n619), .B1(new_n531), .B2(G20), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n337), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n619), .A2(KEYINPUT87), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n299), .A2(new_n531), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(new_n489), .B2(new_n531), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n621), .A2(new_n622), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n616), .A2(new_n617), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  XNOR2_X1  g0430(.A(KEYINPUT89), .B(KEYINPUT21), .ZN(new_n631));
  OAI21_X1  g0431(.A(G169), .B1(new_n612), .B2(new_n614), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n631), .B1(new_n632), .B2(new_n628), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n546), .A2(new_n561), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n556), .A2(new_n341), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n634), .B(new_n635), .C1(G179), .C2(new_n556), .ZN(new_n636));
  OAI211_X1 g0436(.A(KEYINPUT21), .B(G169), .C1(new_n612), .C2(new_n614), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n554), .A2(G270), .B1(G274), .B2(new_n497), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n608), .A2(new_n610), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n639), .B1(new_n606), .B2(new_n604), .ZN(new_n640));
  OAI211_X1 g0440(.A(G179), .B(new_n638), .C1(new_n640), .C2(new_n509), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT88), .B1(new_n642), .B2(new_n627), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT88), .ZN(new_n644));
  AOI211_X1 g0444(.A(new_n644), .B(new_n628), .C1(new_n637), .C2(new_n641), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n633), .B(new_n636), .C1(new_n643), .C2(new_n645), .ZN(new_n646));
  NOR4_X1   g0446(.A1(new_n461), .A2(new_n602), .A3(new_n630), .A4(new_n646), .ZN(G372));
  AND2_X1   g0447(.A1(new_n408), .A2(new_n410), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n455), .A2(new_n343), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n398), .A2(new_n403), .A3(new_n458), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n315), .A2(new_n317), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n306), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n600), .A2(new_n589), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n654), .A2(KEYINPUT92), .A3(KEYINPUT26), .A4(new_n521), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT92), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n600), .A2(new_n519), .A3(new_n589), .A4(new_n511), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n511), .A2(new_n519), .A3(KEYINPUT90), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n600), .A2(new_n589), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT90), .B1(new_n511), .B2(new_n519), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(KEYINPUT91), .B1(new_n665), .B2(KEYINPUT26), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT90), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n520), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n654), .A2(new_n661), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT91), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(new_n670), .A3(new_n658), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n660), .A2(new_n666), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT93), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n672), .A2(new_n673), .A3(new_n589), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n673), .B1(new_n672), .B2(new_n589), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n642), .A2(new_n627), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n676), .A2(new_n633), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n602), .B1(new_n677), .B2(new_n636), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n674), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n653), .B1(new_n679), .B2(new_n461), .ZN(G369));
  OR2_X1    g0480(.A1(new_n643), .A2(new_n645), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n633), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n220), .A2(new_n221), .A3(G13), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(KEYINPUT27), .ZN(new_n684));
  XOR2_X1   g0484(.A(new_n684), .B(KEYINPUT94), .Z(new_n685));
  INV_X1    g0485(.A(G213), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n683), .B2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G343), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n627), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n629), .A2(new_n691), .ZN(new_n692));
  OAI22_X1  g0492(.A1(new_n682), .A2(new_n692), .B1(new_n677), .B2(new_n691), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n636), .A2(new_n690), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n634), .A2(new_n690), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n563), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n696), .B1(new_n636), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n696), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n690), .B1(new_n681), .B2(new_n633), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n699), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n700), .A2(new_n701), .A3(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n232), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n252), .A2(new_n254), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n228), .ZN(new_n708));
  INV_X1    g0508(.A(new_n707), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n708), .B1(new_n711), .B2(KEYINPUT95), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(KEYINPUT95), .B2(new_n711), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n713), .B(KEYINPUT28), .Z(new_n714));
  AND2_X1   g0514(.A1(new_n530), .A2(new_n601), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n646), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n589), .B1(new_n657), .B2(KEYINPUT26), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n717), .B1(KEYINPUT26), .B2(new_n669), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n690), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT29), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n672), .A2(new_n589), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n678), .B1(new_n721), .B2(KEYINPUT93), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n672), .A2(new_n673), .A3(new_n589), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n690), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n720), .B1(new_n724), .B2(KEYINPUT29), .ZN(new_n725));
  INV_X1    g0525(.A(G330), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT96), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n641), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n553), .A2(new_n555), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n729), .A2(new_n585), .A3(new_n510), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n607), .A2(new_n611), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(new_n283), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(KEYINPUT96), .A3(G179), .A4(new_n638), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n728), .A2(new_n730), .A3(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n728), .A2(new_n730), .A3(new_n733), .A4(KEYINPUT30), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n615), .A2(G179), .A3(new_n587), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n517), .A2(new_n518), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n738), .A2(new_n739), .A3(new_n556), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n736), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n690), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(KEYINPUT31), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT31), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n741), .A2(new_n744), .A3(new_n690), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n646), .A2(new_n630), .ZN(new_n747));
  INV_X1    g0547(.A(new_n690), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n747), .A2(new_n715), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n726), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n725), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n714), .B1(new_n752), .B2(G1), .ZN(G364));
  NOR2_X1   g0553(.A1(new_n297), .A2(G20), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n220), .B1(new_n754), .B2(G45), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n707), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n693), .A2(G330), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n695), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT97), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n232), .A2(new_n278), .ZN(new_n761));
  INV_X1    g0561(.A(G355), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n761), .A2(new_n762), .B1(G116), .B2(new_n232), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n705), .A2(new_n538), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(new_n253), .B2(new_n228), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n247), .A2(new_n253), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n763), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G13), .A2(G33), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n229), .B1(G20), .B2(new_n341), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n757), .B1(new_n768), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n771), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n693), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n221), .A2(G179), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n778), .A2(new_n345), .A3(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n463), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n778), .A2(G190), .A3(G200), .ZN(new_n781));
  NOR4_X1   g0581(.A1(new_n221), .A2(new_n326), .A3(new_n345), .A4(G200), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n278), .B1(new_n384), .B2(new_n781), .C1(new_n783), .C2(new_n289), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G179), .A2(G200), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n221), .B1(new_n785), .B2(G190), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n780), .B(new_n784), .C1(G97), .C2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G190), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(new_n345), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n790), .A2(G68), .B1(new_n791), .B2(G50), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n785), .A2(G20), .A3(new_n345), .ZN(new_n793));
  INV_X1    g0593(.A(G159), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT99), .B(KEYINPUT32), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR4_X1   g0597(.A1(new_n221), .A2(new_n326), .A3(G190), .A4(G200), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n798), .A2(KEYINPUT98), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(KEYINPUT98), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G77), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n788), .A2(new_n792), .A3(new_n797), .A4(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n793), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n805), .A2(KEYINPUT100), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(KEYINPUT100), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n779), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n809), .A2(G329), .B1(G283), .B2(new_n810), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT101), .Z(new_n812));
  INV_X1    g0612(.A(G322), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n270), .B1(new_n783), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G294), .B2(new_n787), .ZN(new_n815));
  INV_X1    g0615(.A(new_n791), .ZN(new_n816));
  INV_X1    g0616(.A(G326), .ZN(new_n817));
  INV_X1    g0617(.A(G303), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n816), .A2(new_n817), .B1(new_n781), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(KEYINPUT33), .B(G317), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(new_n790), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G311), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n815), .B(new_n821), .C1(new_n822), .C2(new_n801), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n804), .B1(new_n812), .B2(new_n823), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n775), .B(new_n777), .C1(new_n772), .C2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n760), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G396));
  NAND2_X1  g0627(.A1(new_n339), .A2(new_n690), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n346), .A2(new_n343), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(KEYINPUT103), .B1(new_n343), .B2(new_n748), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n339), .A2(new_n342), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT103), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n831), .A2(new_n832), .A3(new_n327), .A4(new_n690), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n748), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n724), .A2(new_n835), .B1(new_n679), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n757), .B1(new_n837), .B2(new_n751), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n751), .B2(new_n837), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n779), .A2(new_n209), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(G58), .B2(new_n787), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n841), .B(new_n538), .C1(new_n202), .C2(new_n781), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n782), .A2(G143), .B1(G137), .B2(new_n791), .ZN(new_n843));
  INV_X1    g0643(.A(G150), .ZN(new_n844));
  INV_X1    g0644(.A(new_n790), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n843), .B1(new_n844), .B2(new_n845), .C1(new_n801), .C2(new_n794), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT34), .Z(new_n847));
  AOI211_X1 g0647(.A(new_n842), .B(new_n847), .C1(G132), .C2(new_n809), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n278), .B1(new_n782), .B2(G294), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n849), .B1(new_n428), .B2(new_n786), .C1(new_n808), .C2(new_n822), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n801), .A2(new_n531), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n384), .A2(new_n779), .B1(new_n781), .B2(new_n463), .ZN(new_n852));
  XOR2_X1   g0652(.A(KEYINPUT102), .B(G283), .Z(new_n853));
  OAI22_X1  g0653(.A1(new_n845), .A2(new_n853), .B1(new_n816), .B2(new_n818), .ZN(new_n854));
  NOR4_X1   g0654(.A1(new_n850), .A2(new_n851), .A3(new_n852), .A4(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n772), .B1(new_n848), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n757), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n772), .A2(new_n769), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n857), .B1(new_n211), .B2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n856), .B(new_n859), .C1(new_n835), .C2(new_n770), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n839), .A2(new_n860), .ZN(G384));
  NOR2_X1   g0661(.A1(new_n754), .A2(new_n220), .ZN(new_n862));
  INV_X1    g0662(.A(new_n461), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n863), .B(new_n720), .C1(new_n724), .C2(KEYINPUT29), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n864), .A2(new_n653), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT105), .ZN(new_n866));
  INV_X1    g0666(.A(new_n688), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n648), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n867), .B1(new_n400), .B2(new_n401), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n396), .A2(new_n407), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT37), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n396), .A2(new_n407), .A3(new_n869), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n412), .B2(new_n869), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n364), .A2(new_n351), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n295), .B1(new_n878), .B2(new_n376), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n366), .A2(new_n879), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n880), .A2(new_n395), .B1(new_n404), .B2(new_n405), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n688), .B1(new_n880), .B2(new_n395), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n881), .A2(new_n882), .A3(new_n402), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n873), .B1(new_n883), .B2(new_n872), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n411), .A2(new_n882), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n877), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT39), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT38), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT38), .B1(new_n884), .B2(new_n885), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT39), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n455), .A2(new_n690), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n868), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n884), .A2(new_n885), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n876), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n886), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n748), .A2(new_n424), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n455), .A2(new_n458), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n903), .B1(new_n455), .B2(new_n458), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n836), .B1(new_n722), .B2(new_n723), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n343), .A2(new_n690), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n901), .B(new_n907), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n898), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n866), .B(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n835), .B1(new_n904), .B2(new_n905), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n746), .B2(new_n749), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n901), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT40), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n877), .B2(new_n886), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n916), .A2(new_n917), .B1(new_n918), .B2(new_n915), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n461), .B1(new_n746), .B2(new_n749), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT106), .ZN(new_n922));
  OR2_X1    g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n920), .A2(new_n922), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(G330), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n862), .B1(new_n913), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n913), .B2(new_n925), .ZN(new_n927));
  INV_X1    g0727(.A(new_n482), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n928), .A2(KEYINPUT35), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(KEYINPUT35), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n929), .A2(new_n930), .A3(G116), .A4(new_n230), .ZN(new_n931));
  XOR2_X1   g0731(.A(KEYINPUT104), .B(KEYINPUT36), .Z(new_n932));
  XNOR2_X1  g0732(.A(new_n931), .B(new_n932), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n228), .B(G77), .C1(new_n289), .C2(new_n209), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(G50), .B2(new_n209), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(G1), .A3(new_n297), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n927), .A2(new_n933), .A3(new_n936), .ZN(G367));
  OAI21_X1  g0737(.A(new_n530), .B1(new_n525), .B2(new_n748), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n521), .A2(new_n690), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n940), .A2(new_n703), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n942), .A2(KEYINPUT42), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n938), .A2(new_n636), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n690), .B1(new_n944), .B2(new_n520), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n942), .B2(KEYINPUT42), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n748), .A2(new_n599), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n663), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n589), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n948), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT43), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n947), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n943), .A2(new_n946), .A3(new_n954), .A4(new_n953), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n700), .A2(new_n940), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n707), .B(KEYINPUT41), .Z(new_n962));
  NAND2_X1  g0762(.A1(new_n703), .A2(new_n701), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n940), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT44), .Z(new_n965));
  NOR2_X1   g0765(.A1(new_n963), .A2(new_n940), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT45), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n968), .A2(new_n695), .A3(new_n699), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n702), .B(new_n699), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n695), .B(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n965), .A2(new_n700), .A3(new_n967), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n969), .A2(new_n752), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n962), .B1(new_n973), .B2(new_n752), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n961), .B1(new_n974), .B2(new_n756), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n773), .B1(new_n232), .B2(new_n335), .C1(new_n765), .C2(new_n243), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n976), .A2(new_n757), .ZN(new_n977));
  INV_X1    g0777(.A(new_n609), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n783), .A2(new_n978), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n538), .B(new_n979), .C1(G317), .C2(new_n805), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n779), .A2(new_n428), .ZN(new_n981));
  INV_X1    g0781(.A(G294), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n845), .A2(new_n982), .B1(new_n786), .B2(new_n463), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n981), .B(new_n983), .C1(G311), .C2(new_n791), .ZN(new_n984));
  INV_X1    g0784(.A(new_n853), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n802), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n781), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(G116), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT46), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n980), .A2(new_n984), .A3(new_n986), .A4(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n779), .A2(new_n211), .ZN(new_n991));
  INV_X1    g0791(.A(G137), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n278), .B1(new_n793), .B2(new_n992), .C1(new_n783), .C2(new_n844), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n991), .B(new_n993), .C1(G159), .C2(new_n790), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n202), .B2(new_n801), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n786), .A2(new_n209), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n791), .B2(G143), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n289), .B2(new_n781), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n990), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT47), .Z(new_n1000));
  INV_X1    g0800(.A(new_n772), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n977), .B1(new_n952), .B2(new_n776), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n975), .A2(new_n1002), .ZN(G387));
  AOI21_X1  g0803(.A(new_n709), .B1(new_n752), .B2(new_n971), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n752), .B2(new_n971), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n240), .A2(new_n253), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT108), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n287), .A2(G50), .ZN(new_n1008));
  XOR2_X1   g0808(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n1009));
  XNOR2_X1  g0809(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n710), .B(new_n253), .C1(new_n209), .C2(new_n211), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n764), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1006), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(G107), .B2(new_n232), .C1(new_n710), .C2(new_n761), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n857), .B1(new_n1015), .B2(new_n773), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n801), .A2(new_n209), .B1(new_n391), .B2(new_n845), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT109), .Z(new_n1018));
  NOR2_X1   g0818(.A1(new_n781), .A2(new_n211), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n981), .B(new_n1019), .C1(G159), .C2(new_n791), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n572), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n787), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n783), .A2(new_n202), .B1(new_n844), .B2(new_n793), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1023), .A2(new_n381), .ZN(new_n1024));
  AND4_X1   g0824(.A1(new_n1018), .A2(new_n1020), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n782), .A2(G317), .B1(G311), .B2(new_n790), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n813), .B2(new_n816), .C1(new_n801), .C2(new_n978), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT48), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n787), .A2(new_n985), .B1(new_n987), .B2(G294), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT49), .Z(new_n1033));
  OR2_X1    g0833(.A1(new_n1033), .A2(KEYINPUT110), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n381), .B1(new_n531), .B2(new_n779), .C1(new_n817), .C2(new_n793), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT111), .Z(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n1033), .B2(KEYINPUT110), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1025), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1016), .B1(new_n1038), .B2(new_n1001), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n699), .A2(new_n776), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n971), .B2(new_n756), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1005), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT112), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1005), .A2(KEYINPUT112), .A3(new_n1042), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(G393));
  NAND2_X1  g0847(.A1(new_n969), .A2(new_n972), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1048), .A2(new_n755), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n940), .A2(new_n771), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n773), .B1(new_n428), .B2(new_n232), .C1(new_n765), .C2(new_n250), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n757), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n782), .A2(G311), .B1(G317), .B2(new_n791), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT52), .Z(new_n1054));
  OAI22_X1  g0854(.A1(new_n978), .A2(new_n845), .B1(new_n531), .B2(new_n786), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n987), .B2(new_n985), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n802), .A2(G294), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n278), .B(new_n780), .C1(G322), .C2(new_n805), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1054), .A2(new_n1056), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n786), .A2(new_n211), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n845), .A2(new_n202), .B1(new_n781), .B2(new_n209), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(G87), .C2(new_n810), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n381), .B1(G143), .B2(new_n805), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(new_n287), .C2(new_n801), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n782), .A2(G159), .B1(G150), .B2(new_n791), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT51), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1059), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1052), .B1(new_n1067), .B2(new_n772), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1049), .B1(new_n1050), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n752), .A2(new_n971), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1048), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1071), .A2(new_n707), .A3(new_n973), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1069), .A2(new_n1072), .ZN(G390));
  NAND2_X1  g0873(.A1(new_n750), .A2(new_n863), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n864), .A2(new_n653), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n745), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n744), .B1(new_n741), .B2(new_n690), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NOR4_X1   g0879(.A1(new_n602), .A2(new_n646), .A3(new_n630), .A4(new_n690), .ZN(new_n1080));
  OAI211_X1 g0880(.A(G330), .B(new_n835), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n906), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n750), .A2(new_n835), .A3(new_n907), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n909), .B1(new_n719), .B2(new_n835), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n909), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n679), .B2(new_n836), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1085), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1076), .A2(new_n1090), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n665), .A2(KEYINPUT91), .A3(KEYINPUT26), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n670), .B1(new_n669), .B2(new_n658), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n655), .A2(new_n659), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(KEYINPUT93), .B1(new_n1095), .B2(new_n950), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n678), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1096), .A2(new_n723), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n836), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n909), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n896), .B1(new_n1100), .B2(new_n906), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n894), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1084), .A2(new_n906), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n887), .A2(new_n896), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1083), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1083), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1108), .B(new_n1105), .C1(new_n1101), .C2(new_n894), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1091), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n895), .B1(new_n1111), .B2(new_n896), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1108), .B1(new_n1112), .B2(new_n1105), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n897), .B1(new_n1087), .B2(new_n907), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1083), .B(new_n1106), .C1(new_n1114), .C2(new_n895), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1075), .A2(new_n1089), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1113), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1110), .A2(new_n707), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1113), .A2(new_n1115), .A3(new_n756), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n801), .A2(new_n428), .B1(new_n463), .B2(new_n845), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1120), .A2(KEYINPUT113), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(KEYINPUT113), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1060), .B(new_n840), .C1(G283), .C2(new_n791), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n270), .B1(new_n384), .B2(new_n781), .C1(new_n783), .C2(new_n531), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n809), .B2(G294), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(G132), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n278), .B1(new_n786), .B2(new_n794), .C1(new_n783), .C2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n809), .B2(G125), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n791), .A2(G128), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1130), .B1(new_n779), .B2(new_n202), .C1(new_n992), .C2(new_n845), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT53), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n781), .B2(new_n844), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n987), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1131), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT54), .B(G143), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1129), .B(new_n1135), .C1(new_n801), .C2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1126), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1001), .B1(new_n1138), .B2(KEYINPUT114), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(KEYINPUT114), .B2(new_n1138), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n858), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1140), .B(new_n757), .C1(new_n392), .C2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n894), .B2(new_n769), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT115), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1119), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1118), .A2(new_n1145), .ZN(G378));
  NAND2_X1  g0946(.A1(new_n1117), .A2(new_n1076), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n304), .A2(new_n688), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n318), .A2(new_n1149), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1148), .B(new_n306), .C1(new_n315), .C2(new_n317), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n1150), .A2(new_n1151), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1153), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n919), .B2(G330), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n905), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n455), .A2(new_n458), .A3(new_n903), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1159), .A2(new_n1160), .B1(new_n829), .B2(new_n834), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n917), .B1(new_n1162), .B2(new_n892), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n918), .A2(new_n915), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT118), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1156), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n1154), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1155), .A2(KEYINPUT118), .A3(new_n1156), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AND4_X1   g0969(.A1(G330), .A2(new_n1163), .A3(new_n1164), .A4(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1158), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n911), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n898), .B(new_n910), .C1(new_n1158), .C2(new_n1170), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1172), .A2(KEYINPUT57), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1147), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1117), .B2(new_n1076), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1175), .B(new_n707), .C1(KEYINPUT57), .C2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n857), .B1(new_n202), .B2(new_n858), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1021), .A2(new_n802), .B1(new_n809), .B2(G283), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n816), .A2(new_n531), .B1(new_n779), .B2(new_n289), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1019), .B(new_n1181), .C1(G97), .C2(new_n790), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n783), .A2(new_n463), .ZN(new_n1183));
  NOR4_X1   g0983(.A1(new_n1183), .A2(new_n538), .A3(new_n706), .A4(new_n996), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1180), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT58), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n202), .B1(G33), .B2(G41), .C1(new_n538), .C2(new_n706), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n791), .A2(G125), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n845), .B2(new_n1127), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G150), .B2(new_n787), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1136), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n987), .A2(new_n1191), .B1(new_n782), .B2(G128), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1190), .B(new_n1192), .C1(new_n992), .C2(new_n801), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT116), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(KEYINPUT59), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n810), .A2(G159), .ZN(new_n1197));
  AOI211_X1 g0997(.A(G33), .B(G41), .C1(new_n805), .C2(G124), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1195), .A2(KEYINPUT59), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1186), .B(new_n1187), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT117), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n772), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1179), .B1(new_n1204), .B2(new_n1205), .C1(new_n1169), .C2(new_n770), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n1176), .B2(new_n755), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT119), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  OAI211_X1 g1009(.A(KEYINPUT119), .B(new_n1206), .C1(new_n1176), .C2(new_n755), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1178), .A2(new_n1211), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT120), .Z(G375));
  INV_X1    g1013(.A(new_n962), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1075), .A2(new_n1089), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1091), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n906), .A2(new_n769), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n757), .B1(G68), .B2(new_n1141), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G107), .A2(new_n802), .B1(new_n809), .B2(G303), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n278), .B(new_n991), .C1(G283), .C2(new_n782), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1219), .A2(new_n1022), .A3(new_n1220), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n987), .A2(G97), .B1(G116), .B2(new_n790), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n982), .B2(new_n816), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n802), .A2(G150), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n809), .A2(G128), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n381), .B1(G137), .B2(new_n782), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n810), .A2(G58), .B1(new_n787), .B2(G50), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n987), .A2(G159), .B1(new_n1191), .B2(new_n790), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1127), .B2(new_n816), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n1221), .A2(new_n1223), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1218), .B1(new_n1231), .B2(new_n772), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1090), .A2(new_n756), .B1(new_n1217), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1216), .A2(new_n1233), .ZN(G381));
  INV_X1    g1034(.A(G390), .ZN(new_n1235));
  INV_X1    g1035(.A(G384), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1045), .A2(new_n826), .A3(new_n1046), .ZN(new_n1238));
  NOR4_X1   g1038(.A1(new_n1237), .A2(new_n1238), .A3(G387), .A4(G381), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT121), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1119), .A2(new_n1144), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n709), .B1(new_n1242), .B2(new_n1091), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1241), .B1(new_n1243), .B2(new_n1117), .ZN(new_n1244));
  INV_X1    g1044(.A(G375), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1240), .A2(new_n1244), .A3(new_n1245), .ZN(G407));
  NOR2_X1   g1046(.A1(new_n686), .A2(G343), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1245), .A2(new_n1244), .A3(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(G407), .A2(G213), .A3(new_n1248), .ZN(G409));
  INV_X1    g1049(.A(new_n1238), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n826), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n1250), .A2(new_n1235), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G393), .A2(G396), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G390), .B1(new_n1253), .B2(new_n1238), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT126), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(new_n975), .B2(new_n1002), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n975), .A2(new_n1255), .A3(new_n1002), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n1252), .A2(new_n1254), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1235), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1258), .A2(new_n1256), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1253), .A2(G390), .A3(new_n1238), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1259), .A2(new_n1263), .ZN(new_n1264));
  XOR2_X1   g1064(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1265));
  OAI21_X1  g1065(.A(KEYINPUT60), .B1(new_n1075), .B2(new_n1089), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n709), .B1(new_n1266), .B2(new_n1215), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1075), .A2(new_n1089), .A3(KEYINPUT60), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1267), .A2(KEYINPUT124), .A3(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT124), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1233), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1236), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G384), .B(new_n1233), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1247), .A2(G2897), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1272), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1274), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT123), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1207), .B1(new_n1177), .B2(new_n1214), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1278), .B1(new_n1279), .B2(G378), .ZN(new_n1280));
  AOI211_X1 g1080(.A(new_n962), .B(new_n1176), .C1(new_n1117), .C2(new_n1076), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1244), .B(KEYINPUT123), .C1(new_n1207), .C2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1280), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1175), .A2(new_n707), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1177), .A2(KEYINPUT57), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G378), .B(new_n1211), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(KEYINPUT122), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT122), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1178), .A2(new_n1288), .A3(G378), .A4(new_n1211), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1283), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1277), .B1(new_n1290), .B2(new_n1247), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1290), .A2(new_n1247), .A3(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT62), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1265), .B(new_n1291), .C1(new_n1293), .C2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1283), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1247), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1292), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1301), .A2(KEYINPUT62), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1264), .B1(new_n1295), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT61), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1259), .A2(new_n1304), .A3(new_n1263), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1305), .B1(new_n1293), .B2(KEYINPUT63), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT125), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1277), .B(new_n1307), .C1(new_n1247), .C2(new_n1290), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1301), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1291), .A2(KEYINPUT125), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1306), .A2(new_n1308), .A3(new_n1310), .A4(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1303), .A2(new_n1312), .ZN(G405));
  NAND2_X1  g1113(.A1(G375), .A2(new_n1244), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1314), .A2(new_n1296), .A3(new_n1292), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1292), .B1(new_n1314), .B2(new_n1296), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1264), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1314), .A2(new_n1296), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1300), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1264), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1314), .A2(new_n1296), .A3(new_n1292), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1319), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1317), .A2(new_n1322), .ZN(G402));
endmodule


