

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U557 ( .A1(n840), .A2(n839), .ZN(n843) );
  OR2_X2 U558 ( .A1(n769), .A2(n784), .ZN(n526) );
  AND2_X1 U559 ( .A1(n759), .A2(n758), .ZN(n762) );
  OR2_X1 U560 ( .A1(n988), .A2(n716), .ZN(n717) );
  NAND2_X1 U561 ( .A1(n747), .A2(n525), .ZN(n752) );
  NOR2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n529) );
  AND2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n908) );
  OR2_X1 U564 ( .A1(G301), .A2(n742), .ZN(n524) );
  XNOR2_X1 U565 ( .A(n746), .B(n745), .ZN(n525) );
  INV_X1 U566 ( .A(G2105), .ZN(n533) );
  XOR2_X1 U567 ( .A(n730), .B(KEYINPUT29), .Z(n527) );
  INV_X2 U568 ( .A(n753), .ZN(n731) );
  NAND2_X2 U569 ( .A1(n705), .A2(n804), .ZN(n753) );
  XOR2_X1 U570 ( .A(KEYINPUT23), .B(n539), .Z(n528) );
  INV_X1 U571 ( .A(KEYINPUT26), .ZN(n712) );
  INV_X1 U572 ( .A(KEYINPUT98), .ZN(n707) );
  INV_X1 U573 ( .A(KEYINPUT99), .ZN(n738) );
  XNOR2_X1 U574 ( .A(n738), .B(KEYINPUT30), .ZN(n739) );
  XNOR2_X1 U575 ( .A(n740), .B(n739), .ZN(n741) );
  NAND2_X1 U576 ( .A1(n527), .A2(n524), .ZN(n747) );
  INV_X1 U577 ( .A(KEYINPUT103), .ZN(n765) );
  XNOR2_X1 U578 ( .A(n760), .B(KEYINPUT101), .ZN(n761) );
  NOR2_X1 U579 ( .A1(G164), .A2(G1384), .ZN(n804) );
  INV_X1 U580 ( .A(n973), .ZN(n773) );
  NOR2_X1 U581 ( .A1(G651), .A2(n648), .ZN(n672) );
  NOR2_X1 U582 ( .A1(n546), .A2(n545), .ZN(n703) );
  BUF_X1 U583 ( .A(n703), .Z(G160) );
  XOR2_X1 U584 ( .A(KEYINPUT17), .B(n529), .Z(n541) );
  INV_X1 U585 ( .A(n541), .ZN(n530) );
  INV_X1 U586 ( .A(n530), .ZN(n904) );
  NAND2_X1 U587 ( .A1(G138), .A2(n904), .ZN(n532) );
  AND2_X1 U588 ( .A1(n533), .A2(G2104), .ZN(n905) );
  NAND2_X1 U589 ( .A1(G102), .A2(n905), .ZN(n531) );
  NAND2_X1 U590 ( .A1(n532), .A2(n531), .ZN(n538) );
  NAND2_X1 U591 ( .A1(G114), .A2(n908), .ZN(n536) );
  NOR2_X1 U592 ( .A1(n533), .A2(G2104), .ZN(n534) );
  XNOR2_X2 U593 ( .A(n534), .B(KEYINPUT64), .ZN(n909) );
  NAND2_X1 U594 ( .A1(G126), .A2(n909), .ZN(n535) );
  NAND2_X1 U595 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U596 ( .A1(n538), .A2(n537), .ZN(G164) );
  NAND2_X1 U597 ( .A1(G125), .A2(n909), .ZN(n540) );
  NAND2_X1 U598 ( .A1(G101), .A2(n905), .ZN(n539) );
  NAND2_X1 U599 ( .A1(n540), .A2(n528), .ZN(n546) );
  NAND2_X1 U600 ( .A1(n908), .A2(G113), .ZN(n543) );
  NAND2_X1 U601 ( .A1(n541), .A2(G137), .ZN(n542) );
  NAND2_X1 U602 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U603 ( .A(n544), .B(KEYINPUT65), .Z(n545) );
  XOR2_X1 U604 ( .A(G2443), .B(G2446), .Z(n548) );
  XNOR2_X1 U605 ( .A(G2427), .B(G2451), .ZN(n547) );
  XNOR2_X1 U606 ( .A(n548), .B(n547), .ZN(n554) );
  XOR2_X1 U607 ( .A(G2430), .B(G2454), .Z(n550) );
  XNOR2_X1 U608 ( .A(G1348), .B(G1341), .ZN(n549) );
  XNOR2_X1 U609 ( .A(n550), .B(n549), .ZN(n552) );
  XOR2_X1 U610 ( .A(G2435), .B(G2438), .Z(n551) );
  XNOR2_X1 U611 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U612 ( .A(n554), .B(n553), .Z(n555) );
  AND2_X1 U613 ( .A1(G14), .A2(n555), .ZN(G401) );
  AND2_X1 U614 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U615 ( .A(G57), .ZN(G237) );
  INV_X1 U616 ( .A(G132), .ZN(G219) );
  INV_X1 U617 ( .A(G82), .ZN(G220) );
  INV_X1 U618 ( .A(G651), .ZN(n561) );
  NOR2_X1 U619 ( .A1(G543), .A2(n561), .ZN(n556) );
  XOR2_X1 U620 ( .A(KEYINPUT1), .B(n556), .Z(n667) );
  NAND2_X1 U621 ( .A1(G63), .A2(n667), .ZN(n558) );
  XOR2_X1 U622 ( .A(G543), .B(KEYINPUT0), .Z(n648) );
  NAND2_X1 U623 ( .A1(G51), .A2(n672), .ZN(n557) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(KEYINPUT6), .B(n559), .ZN(n567) );
  NOR2_X1 U626 ( .A1(G651), .A2(G543), .ZN(n666) );
  NAND2_X1 U627 ( .A1(n666), .A2(G89), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n560), .B(KEYINPUT4), .ZN(n563) );
  NOR2_X1 U629 ( .A1(n648), .A2(n561), .ZN(n663) );
  NAND2_X1 U630 ( .A1(G76), .A2(n663), .ZN(n562) );
  NAND2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U632 ( .A(KEYINPUT75), .B(n564), .ZN(n565) );
  XNOR2_X1 U633 ( .A(KEYINPUT5), .B(n565), .ZN(n566) );
  NOR2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U635 ( .A(KEYINPUT7), .B(n568), .Z(G168) );
  XOR2_X1 U636 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U637 ( .A1(G7), .A2(G661), .ZN(n569) );
  XNOR2_X1 U638 ( .A(n569), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U639 ( .A(G223), .ZN(n844) );
  NAND2_X1 U640 ( .A1(n844), .A2(G567), .ZN(n570) );
  XOR2_X1 U641 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  NAND2_X1 U642 ( .A1(G56), .A2(n667), .ZN(n571) );
  XOR2_X1 U643 ( .A(KEYINPUT14), .B(n571), .Z(n577) );
  NAND2_X1 U644 ( .A1(n666), .A2(G81), .ZN(n572) );
  XNOR2_X1 U645 ( .A(n572), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U646 ( .A1(G68), .A2(n663), .ZN(n573) );
  NAND2_X1 U647 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U648 ( .A(KEYINPUT13), .B(n575), .Z(n576) );
  NOR2_X1 U649 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U650 ( .A1(n672), .A2(G43), .ZN(n578) );
  NAND2_X1 U651 ( .A1(n579), .A2(n578), .ZN(n988) );
  INV_X1 U652 ( .A(G860), .ZN(n638) );
  OR2_X1 U653 ( .A1(n988), .A2(n638), .ZN(G153) );
  NAND2_X1 U654 ( .A1(n663), .A2(G77), .ZN(n580) );
  XNOR2_X1 U655 ( .A(n580), .B(KEYINPUT68), .ZN(n582) );
  NAND2_X1 U656 ( .A1(G90), .A2(n666), .ZN(n581) );
  NAND2_X1 U657 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U658 ( .A(KEYINPUT9), .B(n583), .ZN(n587) );
  NAND2_X1 U659 ( .A1(G64), .A2(n667), .ZN(n585) );
  NAND2_X1 U660 ( .A1(G52), .A2(n672), .ZN(n584) );
  AND2_X1 U661 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U662 ( .A1(n587), .A2(n586), .ZN(G301) );
  NAND2_X1 U663 ( .A1(G79), .A2(n663), .ZN(n588) );
  XNOR2_X1 U664 ( .A(n588), .B(KEYINPUT72), .ZN(n595) );
  NAND2_X1 U665 ( .A1(G66), .A2(n667), .ZN(n590) );
  NAND2_X1 U666 ( .A1(G54), .A2(n672), .ZN(n589) );
  NAND2_X1 U667 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U668 ( .A1(G92), .A2(n666), .ZN(n591) );
  XNOR2_X1 U669 ( .A(KEYINPUT71), .B(n591), .ZN(n592) );
  NOR2_X1 U670 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U671 ( .A1(n595), .A2(n594), .ZN(n597) );
  XOR2_X1 U672 ( .A(KEYINPUT73), .B(KEYINPUT15), .Z(n596) );
  XNOR2_X1 U673 ( .A(n597), .B(n596), .ZN(n871) );
  INV_X1 U674 ( .A(n871), .ZN(n977) );
  NOR2_X1 U675 ( .A1(G868), .A2(n977), .ZN(n599) );
  INV_X1 U676 ( .A(G868), .ZN(n685) );
  NOR2_X1 U677 ( .A1(n685), .A2(G301), .ZN(n598) );
  NOR2_X1 U678 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U679 ( .A(KEYINPUT74), .B(n600), .ZN(G284) );
  NAND2_X1 U680 ( .A1(n667), .A2(G65), .ZN(n603) );
  NAND2_X1 U681 ( .A1(G53), .A2(n672), .ZN(n601) );
  XOR2_X1 U682 ( .A(KEYINPUT69), .B(n601), .Z(n602) );
  NAND2_X1 U683 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U684 ( .A1(G91), .A2(n666), .ZN(n605) );
  NAND2_X1 U685 ( .A1(G78), .A2(n663), .ZN(n604) );
  NAND2_X1 U686 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U687 ( .A1(n607), .A2(n606), .ZN(n976) );
  XOR2_X1 U688 ( .A(n976), .B(KEYINPUT70), .Z(G299) );
  NOR2_X1 U689 ( .A1(G299), .A2(G868), .ZN(n609) );
  NOR2_X1 U690 ( .A1(G286), .A2(n685), .ZN(n608) );
  NOR2_X1 U691 ( .A1(n609), .A2(n608), .ZN(G297) );
  NAND2_X1 U692 ( .A1(n638), .A2(G559), .ZN(n610) );
  NAND2_X1 U693 ( .A1(n610), .A2(n871), .ZN(n611) );
  XNOR2_X1 U694 ( .A(n611), .B(KEYINPUT16), .ZN(n613) );
  XOR2_X1 U695 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n612) );
  XNOR2_X1 U696 ( .A(n613), .B(n612), .ZN(G148) );
  NOR2_X1 U697 ( .A1(G868), .A2(n988), .ZN(n614) );
  XNOR2_X1 U698 ( .A(KEYINPUT78), .B(n614), .ZN(n617) );
  NAND2_X1 U699 ( .A1(G868), .A2(n871), .ZN(n615) );
  NOR2_X1 U700 ( .A1(G559), .A2(n615), .ZN(n616) );
  NOR2_X1 U701 ( .A1(n617), .A2(n616), .ZN(G282) );
  XNOR2_X1 U702 ( .A(G2096), .B(KEYINPUT82), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n905), .A2(G99), .ZN(n618) );
  XNOR2_X1 U704 ( .A(n618), .B(KEYINPUT80), .ZN(n620) );
  NAND2_X1 U705 ( .A1(G111), .A2(n908), .ZN(n619) );
  NAND2_X1 U706 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U707 ( .A(KEYINPUT81), .B(n621), .ZN(n627) );
  NAND2_X1 U708 ( .A1(G123), .A2(n909), .ZN(n622) );
  XNOR2_X1 U709 ( .A(n622), .B(KEYINPUT18), .ZN(n624) );
  NAND2_X1 U710 ( .A1(G135), .A2(n904), .ZN(n623) );
  NAND2_X1 U711 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U712 ( .A(KEYINPUT79), .B(n625), .ZN(n626) );
  NAND2_X1 U713 ( .A1(n627), .A2(n626), .ZN(n954) );
  XNOR2_X1 U714 ( .A(n628), .B(n954), .ZN(n629) );
  NOR2_X1 U715 ( .A1(G2100), .A2(n629), .ZN(n630) );
  XNOR2_X1 U716 ( .A(KEYINPUT83), .B(n630), .ZN(G156) );
  NAND2_X1 U717 ( .A1(G93), .A2(n666), .ZN(n632) );
  NAND2_X1 U718 ( .A1(G67), .A2(n667), .ZN(n631) );
  NAND2_X1 U719 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U720 ( .A1(G80), .A2(n663), .ZN(n634) );
  NAND2_X1 U721 ( .A1(G55), .A2(n672), .ZN(n633) );
  NAND2_X1 U722 ( .A1(n634), .A2(n633), .ZN(n635) );
  OR2_X1 U723 ( .A1(n636), .A2(n635), .ZN(n684) );
  XNOR2_X1 U724 ( .A(n684), .B(KEYINPUT84), .ZN(n640) );
  NAND2_X1 U725 ( .A1(G559), .A2(n871), .ZN(n637) );
  XOR2_X1 U726 ( .A(n988), .B(n637), .Z(n682) );
  NAND2_X1 U727 ( .A1(n682), .A2(n638), .ZN(n639) );
  XNOR2_X1 U728 ( .A(n640), .B(n639), .ZN(G145) );
  NAND2_X1 U729 ( .A1(G75), .A2(n663), .ZN(n642) );
  NAND2_X1 U730 ( .A1(G62), .A2(n667), .ZN(n641) );
  NAND2_X1 U731 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U732 ( .A1(G88), .A2(n666), .ZN(n643) );
  XNOR2_X1 U733 ( .A(KEYINPUT87), .B(n643), .ZN(n644) );
  NOR2_X1 U734 ( .A1(n645), .A2(n644), .ZN(n647) );
  NAND2_X1 U735 ( .A1(n672), .A2(G50), .ZN(n646) );
  NAND2_X1 U736 ( .A1(n647), .A2(n646), .ZN(G303) );
  INV_X1 U737 ( .A(G303), .ZN(G166) );
  NAND2_X1 U738 ( .A1(G49), .A2(n672), .ZN(n650) );
  NAND2_X1 U739 ( .A1(G87), .A2(n648), .ZN(n649) );
  NAND2_X1 U740 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U741 ( .A1(n667), .A2(n651), .ZN(n654) );
  NAND2_X1 U742 ( .A1(G74), .A2(G651), .ZN(n652) );
  XOR2_X1 U743 ( .A(KEYINPUT85), .B(n652), .Z(n653) );
  NAND2_X1 U744 ( .A1(n654), .A2(n653), .ZN(G288) );
  NAND2_X1 U745 ( .A1(G85), .A2(n666), .ZN(n655) );
  XNOR2_X1 U746 ( .A(n655), .B(KEYINPUT66), .ZN(n657) );
  NAND2_X1 U747 ( .A1(n667), .A2(G60), .ZN(n656) );
  NAND2_X1 U748 ( .A1(n657), .A2(n656), .ZN(n660) );
  NAND2_X1 U749 ( .A1(G72), .A2(n663), .ZN(n658) );
  XNOR2_X1 U750 ( .A(KEYINPUT67), .B(n658), .ZN(n659) );
  NOR2_X1 U751 ( .A1(n660), .A2(n659), .ZN(n662) );
  NAND2_X1 U752 ( .A1(n672), .A2(G47), .ZN(n661) );
  NAND2_X1 U753 ( .A1(n662), .A2(n661), .ZN(G290) );
  XOR2_X1 U754 ( .A(KEYINPUT86), .B(KEYINPUT2), .Z(n665) );
  NAND2_X1 U755 ( .A1(G73), .A2(n663), .ZN(n664) );
  XNOR2_X1 U756 ( .A(n665), .B(n664), .ZN(n671) );
  NAND2_X1 U757 ( .A1(G86), .A2(n666), .ZN(n669) );
  NAND2_X1 U758 ( .A1(G61), .A2(n667), .ZN(n668) );
  NAND2_X1 U759 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U760 ( .A1(n671), .A2(n670), .ZN(n674) );
  NAND2_X1 U761 ( .A1(n672), .A2(G48), .ZN(n673) );
  NAND2_X1 U762 ( .A1(n674), .A2(n673), .ZN(G305) );
  XOR2_X1 U763 ( .A(KEYINPUT89), .B(KEYINPUT19), .Z(n676) );
  XNOR2_X1 U764 ( .A(G166), .B(KEYINPUT88), .ZN(n675) );
  XNOR2_X1 U765 ( .A(n676), .B(n675), .ZN(n677) );
  XOR2_X1 U766 ( .A(n684), .B(n677), .Z(n679) );
  XNOR2_X1 U767 ( .A(G288), .B(G299), .ZN(n678) );
  XNOR2_X1 U768 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U769 ( .A(n680), .B(G290), .ZN(n681) );
  XNOR2_X1 U770 ( .A(n681), .B(G305), .ZN(n870) );
  XNOR2_X1 U771 ( .A(n682), .B(n870), .ZN(n683) );
  NAND2_X1 U772 ( .A1(n683), .A2(G868), .ZN(n687) );
  NAND2_X1 U773 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U774 ( .A1(n687), .A2(n686), .ZN(G295) );
  XOR2_X1 U775 ( .A(KEYINPUT90), .B(KEYINPUT20), .Z(n689) );
  NAND2_X1 U776 ( .A1(G2078), .A2(G2084), .ZN(n688) );
  XNOR2_X1 U777 ( .A(n689), .B(n688), .ZN(n690) );
  NAND2_X1 U778 ( .A1(n690), .A2(G2090), .ZN(n691) );
  XOR2_X1 U779 ( .A(KEYINPUT21), .B(n691), .Z(n692) );
  XNOR2_X1 U780 ( .A(KEYINPUT91), .B(n692), .ZN(n693) );
  NAND2_X1 U781 ( .A1(n693), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U782 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U783 ( .A1(G220), .A2(G219), .ZN(n694) );
  XOR2_X1 U784 ( .A(KEYINPUT22), .B(n694), .Z(n695) );
  NOR2_X1 U785 ( .A1(G218), .A2(n695), .ZN(n696) );
  NAND2_X1 U786 ( .A1(G96), .A2(n696), .ZN(n848) );
  NAND2_X1 U787 ( .A1(n848), .A2(G2106), .ZN(n700) );
  NAND2_X1 U788 ( .A1(G69), .A2(G120), .ZN(n697) );
  NOR2_X1 U789 ( .A1(G237), .A2(n697), .ZN(n698) );
  NAND2_X1 U790 ( .A1(G108), .A2(n698), .ZN(n849) );
  NAND2_X1 U791 ( .A1(n849), .A2(G567), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n850) );
  NAND2_X1 U793 ( .A1(G661), .A2(G483), .ZN(n701) );
  NOR2_X1 U794 ( .A1(n850), .A2(n701), .ZN(n847) );
  NAND2_X1 U795 ( .A1(n847), .A2(G36), .ZN(G176) );
  NOR2_X1 U796 ( .A1(G1976), .A2(G288), .ZN(n771) );
  NOR2_X1 U797 ( .A1(G1971), .A2(G303), .ZN(n702) );
  NOR2_X1 U798 ( .A1(n771), .A2(n702), .ZN(n991) );
  NAND2_X1 U799 ( .A1(G40), .A2(n703), .ZN(n704) );
  XNOR2_X1 U800 ( .A(n704), .B(KEYINPUT92), .ZN(n805) );
  INV_X1 U801 ( .A(n805), .ZN(n705) );
  NOR2_X1 U802 ( .A1(G2084), .A2(n753), .ZN(n735) );
  NAND2_X1 U803 ( .A1(n735), .A2(G8), .ZN(n751) );
  NAND2_X1 U804 ( .A1(G8), .A2(n753), .ZN(n784) );
  NOR2_X1 U805 ( .A1(G1966), .A2(n784), .ZN(n749) );
  NAND2_X1 U806 ( .A1(G1348), .A2(n753), .ZN(n706) );
  XNOR2_X1 U807 ( .A(KEYINPUT97), .B(n706), .ZN(n710) );
  NAND2_X1 U808 ( .A1(n731), .A2(G2067), .ZN(n708) );
  XNOR2_X1 U809 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U810 ( .A1(n710), .A2(n709), .ZN(n711) );
  OR2_X1 U811 ( .A1(n711), .A2(n871), .ZN(n720) );
  NAND2_X1 U812 ( .A1(n871), .A2(n711), .ZN(n718) );
  AND2_X1 U813 ( .A1(n731), .A2(G1996), .ZN(n713) );
  XNOR2_X1 U814 ( .A(n713), .B(n712), .ZN(n715) );
  NAND2_X1 U815 ( .A1(n753), .A2(G1341), .ZN(n714) );
  NAND2_X1 U816 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U817 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U818 ( .A1(n720), .A2(n719), .ZN(n725) );
  NAND2_X1 U819 ( .A1(n731), .A2(G2072), .ZN(n721) );
  XNOR2_X1 U820 ( .A(n721), .B(KEYINPUT27), .ZN(n723) );
  XOR2_X1 U821 ( .A(KEYINPUT96), .B(G1956), .Z(n1010) );
  NOR2_X1 U822 ( .A1(n731), .A2(n1010), .ZN(n722) );
  NOR2_X1 U823 ( .A1(n723), .A2(n722), .ZN(n726) );
  NAND2_X1 U824 ( .A1(n976), .A2(n726), .ZN(n724) );
  NAND2_X1 U825 ( .A1(n725), .A2(n724), .ZN(n729) );
  NOR2_X1 U826 ( .A1(n976), .A2(n726), .ZN(n727) );
  XOR2_X1 U827 ( .A(n727), .B(KEYINPUT28), .Z(n728) );
  NAND2_X1 U828 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U829 ( .A1(G1961), .A2(n753), .ZN(n733) );
  XOR2_X1 U830 ( .A(G2078), .B(KEYINPUT25), .Z(n931) );
  NAND2_X1 U831 ( .A1(n731), .A2(n931), .ZN(n732) );
  NAND2_X1 U832 ( .A1(n733), .A2(n732), .ZN(n742) );
  XOR2_X1 U833 ( .A(KEYINPUT31), .B(KEYINPUT100), .Z(n746) );
  OR2_X1 U834 ( .A1(G1966), .A2(n784), .ZN(n737) );
  INV_X1 U835 ( .A(G8), .ZN(n734) );
  NOR2_X1 U836 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U837 ( .A1(n737), .A2(n736), .ZN(n740) );
  NOR2_X1 U838 ( .A1(G168), .A2(n741), .ZN(n744) );
  AND2_X1 U839 ( .A1(G301), .A2(n742), .ZN(n743) );
  NOR2_X1 U840 ( .A1(n744), .A2(n743), .ZN(n745) );
  INV_X1 U841 ( .A(n752), .ZN(n748) );
  NOR2_X1 U842 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U843 ( .A1(n751), .A2(n750), .ZN(n764) );
  NAND2_X1 U844 ( .A1(n752), .A2(G286), .ZN(n759) );
  NOR2_X1 U845 ( .A1(G1971), .A2(n784), .ZN(n755) );
  NOR2_X1 U846 ( .A1(G2090), .A2(n753), .ZN(n754) );
  NOR2_X1 U847 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U848 ( .A1(n756), .A2(G303), .ZN(n757) );
  OR2_X1 U849 ( .A1(n734), .A2(n757), .ZN(n758) );
  XOR2_X1 U850 ( .A(KEYINPUT102), .B(KEYINPUT32), .Z(n760) );
  XNOR2_X1 U851 ( .A(n762), .B(n761), .ZN(n763) );
  NAND2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n781) );
  NAND2_X1 U853 ( .A1(n991), .A2(n781), .ZN(n766) );
  XNOR2_X1 U854 ( .A(n766), .B(n765), .ZN(n767) );
  NAND2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n987) );
  NAND2_X1 U856 ( .A1(n767), .A2(n987), .ZN(n768) );
  XNOR2_X1 U857 ( .A(KEYINPUT104), .B(n768), .ZN(n769) );
  INV_X1 U858 ( .A(KEYINPUT33), .ZN(n770) );
  NAND2_X1 U859 ( .A1(n526), .A2(n770), .ZN(n776) );
  NAND2_X1 U860 ( .A1(n771), .A2(KEYINPUT33), .ZN(n772) );
  NOR2_X1 U861 ( .A1(n772), .A2(n784), .ZN(n774) );
  XOR2_X1 U862 ( .A(G1981), .B(G305), .Z(n973) );
  NOR2_X1 U863 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n778) );
  INV_X1 U865 ( .A(KEYINPUT105), .ZN(n777) );
  XNOR2_X1 U866 ( .A(n778), .B(n777), .ZN(n830) );
  NOR2_X1 U867 ( .A1(G1981), .A2(G305), .ZN(n779) );
  XOR2_X1 U868 ( .A(n779), .B(KEYINPUT24), .Z(n780) );
  NOR2_X1 U869 ( .A1(n784), .A2(n780), .ZN(n787) );
  NOR2_X1 U870 ( .A1(G2090), .A2(G303), .ZN(n782) );
  NAND2_X1 U871 ( .A1(G8), .A2(n782), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n781), .A2(n783), .ZN(n785) );
  AND2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n828) );
  XNOR2_X1 U875 ( .A(KEYINPUT39), .B(KEYINPUT106), .ZN(n812) );
  NAND2_X1 U876 ( .A1(G141), .A2(n904), .ZN(n789) );
  NAND2_X1 U877 ( .A1(G129), .A2(n909), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U879 ( .A1(n905), .A2(G105), .ZN(n790) );
  XOR2_X1 U880 ( .A(KEYINPUT38), .B(n790), .Z(n791) );
  NOR2_X1 U881 ( .A1(n792), .A2(n791), .ZN(n794) );
  NAND2_X1 U882 ( .A1(n908), .A2(G117), .ZN(n793) );
  NAND2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n899) );
  NOR2_X1 U884 ( .A1(G1996), .A2(n899), .ZN(n957) );
  NAND2_X1 U885 ( .A1(G107), .A2(n908), .ZN(n796) );
  NAND2_X1 U886 ( .A1(G95), .A2(n905), .ZN(n795) );
  NAND2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n800) );
  NAND2_X1 U888 ( .A1(G131), .A2(n904), .ZN(n798) );
  NAND2_X1 U889 ( .A1(G119), .A2(n909), .ZN(n797) );
  NAND2_X1 U890 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U891 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U892 ( .A(n801), .B(KEYINPUT95), .ZN(n885) );
  AND2_X1 U893 ( .A1(n885), .A2(G1991), .ZN(n803) );
  AND2_X1 U894 ( .A1(n899), .A2(G1996), .ZN(n802) );
  NOR2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n950) );
  INV_X1 U896 ( .A(n950), .ZN(n806) );
  NOR2_X1 U897 ( .A1(n805), .A2(n804), .ZN(n834) );
  NAND2_X1 U898 ( .A1(n806), .A2(n834), .ZN(n833) );
  INV_X1 U899 ( .A(n833), .ZN(n809) );
  NOR2_X1 U900 ( .A1(G1991), .A2(n885), .ZN(n953) );
  NOR2_X1 U901 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U902 ( .A1(n953), .A2(n807), .ZN(n808) );
  NOR2_X1 U903 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U904 ( .A1(n957), .A2(n810), .ZN(n811) );
  XNOR2_X1 U905 ( .A(n812), .B(n811), .ZN(n824) );
  NAND2_X1 U906 ( .A1(n904), .A2(G140), .ZN(n813) );
  XOR2_X1 U907 ( .A(KEYINPUT93), .B(n813), .Z(n815) );
  NAND2_X1 U908 ( .A1(n905), .A2(G104), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U910 ( .A(KEYINPUT34), .B(n816), .ZN(n821) );
  NAND2_X1 U911 ( .A1(G116), .A2(n908), .ZN(n818) );
  NAND2_X1 U912 ( .A1(G128), .A2(n909), .ZN(n817) );
  NAND2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n819) );
  XOR2_X1 U914 ( .A(KEYINPUT35), .B(n819), .Z(n820) );
  NOR2_X1 U915 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U916 ( .A(KEYINPUT36), .B(n822), .ZN(n917) );
  XNOR2_X1 U917 ( .A(KEYINPUT37), .B(G2067), .ZN(n825) );
  NOR2_X1 U918 ( .A1(n917), .A2(n825), .ZN(n961) );
  NAND2_X1 U919 ( .A1(n961), .A2(n834), .ZN(n823) );
  XNOR2_X1 U920 ( .A(n823), .B(KEYINPUT94), .ZN(n832) );
  NAND2_X1 U921 ( .A1(n824), .A2(n832), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n917), .A2(n825), .ZN(n962) );
  NAND2_X1 U923 ( .A1(n826), .A2(n962), .ZN(n827) );
  NAND2_X1 U924 ( .A1(n827), .A2(n834), .ZN(n831) );
  AND2_X1 U925 ( .A1(n828), .A2(n831), .ZN(n829) );
  NAND2_X1 U926 ( .A1(n830), .A2(n829), .ZN(n840) );
  INV_X1 U927 ( .A(n831), .ZN(n838) );
  NAND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(n836) );
  XNOR2_X1 U929 ( .A(G1986), .B(G290), .ZN(n979) );
  AND2_X1 U930 ( .A1(n979), .A2(n834), .ZN(n835) );
  NOR2_X1 U931 ( .A1(n836), .A2(n835), .ZN(n837) );
  OR2_X1 U932 ( .A1(n838), .A2(n837), .ZN(n839) );
  XOR2_X1 U933 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n841) );
  XNOR2_X1 U934 ( .A(KEYINPUT40), .B(n841), .ZN(n842) );
  XNOR2_X1 U935 ( .A(n843), .B(n842), .ZN(G329) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n844), .ZN(G217) );
  AND2_X1 U937 ( .A1(G15), .A2(G2), .ZN(n845) );
  NAND2_X1 U938 ( .A1(G661), .A2(n845), .ZN(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n846) );
  NAND2_X1 U940 ( .A1(n847), .A2(n846), .ZN(G188) );
  INV_X1 U942 ( .A(G120), .ZN(G236) );
  INV_X1 U943 ( .A(G96), .ZN(G221) );
  INV_X1 U944 ( .A(G69), .ZN(G235) );
  NOR2_X1 U945 ( .A1(n849), .A2(n848), .ZN(G325) );
  INV_X1 U946 ( .A(G325), .ZN(G261) );
  INV_X1 U947 ( .A(n850), .ZN(G319) );
  XNOR2_X1 U948 ( .A(G1966), .B(G2474), .ZN(n860) );
  XOR2_X1 U949 ( .A(G1976), .B(G1961), .Z(n852) );
  XNOR2_X1 U950 ( .A(G1986), .B(G1971), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U952 ( .A(G1981), .B(G1956), .Z(n854) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1991), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U955 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U956 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(G229) );
  XOR2_X1 U959 ( .A(KEYINPUT109), .B(G2072), .Z(n862) );
  XNOR2_X1 U960 ( .A(G2090), .B(G2078), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U962 ( .A(n863), .B(G2100), .Z(n865) );
  XNOR2_X1 U963 ( .A(G2067), .B(G2084), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U965 ( .A(G2096), .B(KEYINPUT43), .Z(n867) );
  XNOR2_X1 U966 ( .A(G2678), .B(KEYINPUT42), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U968 ( .A(n869), .B(n868), .Z(G227) );
  INV_X1 U969 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U970 ( .A(n988), .B(n870), .ZN(n873) );
  XNOR2_X1 U971 ( .A(G171), .B(n871), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n874), .B(G286), .ZN(n875) );
  NOR2_X1 U974 ( .A1(G37), .A2(n875), .ZN(G397) );
  NAND2_X1 U975 ( .A1(n909), .A2(G124), .ZN(n876) );
  XNOR2_X1 U976 ( .A(n876), .B(KEYINPUT44), .ZN(n883) );
  NAND2_X1 U977 ( .A1(G112), .A2(n908), .ZN(n878) );
  NAND2_X1 U978 ( .A1(G100), .A2(n905), .ZN(n877) );
  NAND2_X1 U979 ( .A1(n878), .A2(n877), .ZN(n881) );
  NAND2_X1 U980 ( .A1(G136), .A2(n904), .ZN(n879) );
  XNOR2_X1 U981 ( .A(KEYINPUT111), .B(n879), .ZN(n880) );
  NOR2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U984 ( .A(KEYINPUT112), .B(n884), .Z(G162) );
  XNOR2_X1 U985 ( .A(G164), .B(n885), .ZN(n886) );
  XNOR2_X1 U986 ( .A(n886), .B(G162), .ZN(n903) );
  XOR2_X1 U987 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n888) );
  XNOR2_X1 U988 ( .A(KEYINPUT48), .B(KEYINPUT114), .ZN(n887) );
  XNOR2_X1 U989 ( .A(n888), .B(n887), .ZN(n898) );
  NAND2_X1 U990 ( .A1(G118), .A2(n908), .ZN(n890) );
  NAND2_X1 U991 ( .A1(G130), .A2(n909), .ZN(n889) );
  NAND2_X1 U992 ( .A1(n890), .A2(n889), .ZN(n896) );
  NAND2_X1 U993 ( .A1(G142), .A2(n904), .ZN(n892) );
  NAND2_X1 U994 ( .A1(G106), .A2(n905), .ZN(n891) );
  NAND2_X1 U995 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U996 ( .A(KEYINPUT45), .B(n893), .ZN(n894) );
  XNOR2_X1 U997 ( .A(KEYINPUT113), .B(n894), .ZN(n895) );
  NOR2_X1 U998 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U999 ( .A(n898), .B(n897), .Z(n901) );
  XOR2_X1 U1000 ( .A(G160), .B(n899), .Z(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n916) );
  NAND2_X1 U1003 ( .A1(G139), .A2(n904), .ZN(n907) );
  NAND2_X1 U1004 ( .A1(G103), .A2(n905), .ZN(n906) );
  NAND2_X1 U1005 ( .A1(n907), .A2(n906), .ZN(n914) );
  NAND2_X1 U1006 ( .A1(G115), .A2(n908), .ZN(n911) );
  NAND2_X1 U1007 ( .A1(G127), .A2(n909), .ZN(n910) );
  NAND2_X1 U1008 ( .A1(n911), .A2(n910), .ZN(n912) );
  XOR2_X1 U1009 ( .A(KEYINPUT47), .B(n912), .Z(n913) );
  NOR2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(n946) );
  XNOR2_X1 U1011 ( .A(n954), .B(n946), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(n916), .B(n915), .ZN(n918) );
  XOR2_X1 U1013 ( .A(n918), .B(n917), .Z(n919) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n919), .ZN(n920) );
  XNOR2_X1 U1015 ( .A(KEYINPUT116), .B(n920), .ZN(G395) );
  NOR2_X1 U1016 ( .A1(G229), .A2(G227), .ZN(n921) );
  XOR2_X1 U1017 ( .A(KEYINPUT49), .B(n921), .Z(n922) );
  NAND2_X1 U1018 ( .A1(G319), .A2(n922), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(G401), .A2(n923), .ZN(n924) );
  XOR2_X1 U1020 ( .A(KEYINPUT117), .B(n924), .Z(n927) );
  NOR2_X1 U1021 ( .A1(G397), .A2(G395), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(KEYINPUT118), .B(n925), .ZN(n926) );
  NAND2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1026 ( .A(G25), .B(G1991), .Z(n928) );
  NAND2_X1 U1027 ( .A1(n928), .A2(G28), .ZN(n937) );
  XNOR2_X1 U1028 ( .A(G2067), .B(G26), .ZN(n930) );
  XNOR2_X1 U1029 ( .A(G33), .B(G2072), .ZN(n929) );
  NOR2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n935) );
  XNOR2_X1 U1031 ( .A(G1996), .B(G32), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(G27), .B(n931), .ZN(n932) );
  NOR2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1036 ( .A(KEYINPUT53), .B(n938), .Z(n941) );
  XOR2_X1 U1037 ( .A(KEYINPUT54), .B(G34), .Z(n939) );
  XNOR2_X1 U1038 ( .A(G2084), .B(n939), .ZN(n940) );
  NAND2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n943) );
  XNOR2_X1 U1040 ( .A(G35), .B(G2090), .ZN(n942) );
  NOR2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(G29), .A2(n944), .ZN(n945) );
  XNOR2_X1 U1043 ( .A(n945), .B(KEYINPUT55), .ZN(n972) );
  XOR2_X1 U1044 ( .A(G2072), .B(n946), .Z(n948) );
  XOR2_X1 U1045 ( .A(G164), .B(G2078), .Z(n947) );
  NOR2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(KEYINPUT50), .B(n949), .ZN(n968) );
  XNOR2_X1 U1048 ( .A(G160), .B(G2084), .ZN(n951) );
  NAND2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n965) );
  XOR2_X1 U1052 ( .A(G2090), .B(G162), .Z(n956) );
  NOR2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1054 ( .A(n958), .B(KEYINPUT119), .Z(n959) );
  XNOR2_X1 U1055 ( .A(KEYINPUT51), .B(n959), .ZN(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(KEYINPUT120), .B(n966), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(KEYINPUT52), .B(n969), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(G29), .A2(n970), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n1027) );
  XOR2_X1 U1064 ( .A(G16), .B(KEYINPUT56), .Z(n996) );
  XNOR2_X1 U1065 ( .A(G168), .B(G1966), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(n975), .B(KEYINPUT57), .ZN(n985) );
  XNOR2_X1 U1068 ( .A(n976), .B(G1956), .ZN(n981) );
  XNOR2_X1 U1069 ( .A(G1348), .B(n977), .ZN(n978) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(G1961), .B(G301), .ZN(n982) );
  NOR2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n994) );
  NAND2_X1 U1075 ( .A1(G1971), .A2(G303), .ZN(n986) );
  NAND2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n990) );
  XNOR2_X1 U1077 ( .A(G1341), .B(n988), .ZN(n989) );
  NOR2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n992) );
  NAND2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1080 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1081 ( .A1(n996), .A2(n995), .ZN(n1024) );
  XNOR2_X1 U1082 ( .A(G1961), .B(KEYINPUT121), .ZN(n997) );
  XNOR2_X1 U1083 ( .A(n997), .B(G5), .ZN(n999) );
  XOR2_X1 U1084 ( .A(G1966), .B(G21), .Z(n998) );
  NAND2_X1 U1085 ( .A1(n999), .A2(n998), .ZN(n1020) );
  XNOR2_X1 U1086 ( .A(G1971), .B(G22), .ZN(n1001) );
  XNOR2_X1 U1087 ( .A(G1976), .B(G23), .ZN(n1000) );
  NOR2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1089 ( .A(KEYINPUT124), .B(n1002), .Z(n1004) );
  XNOR2_X1 U1090 ( .A(G1986), .B(G24), .ZN(n1003) );
  NOR2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(KEYINPUT58), .B(n1005), .ZN(n1018) );
  XOR2_X1 U1093 ( .A(G1348), .B(KEYINPUT59), .Z(n1006) );
  XNOR2_X1 U1094 ( .A(G4), .B(n1006), .ZN(n1015) );
  XNOR2_X1 U1095 ( .A(G1341), .B(G19), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(G6), .B(G1981), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1098 ( .A(KEYINPUT122), .B(n1009), .Z(n1012) );
  XOR2_X1 U1099 ( .A(n1010), .B(G20), .Z(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(n1013), .B(KEYINPUT123), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(KEYINPUT60), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1106 ( .A(KEYINPUT61), .B(n1021), .Z(n1022) );
  NOR2_X1 U1107 ( .A1(G16), .A2(n1022), .ZN(n1023) );
  NOR2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1109 ( .A(KEYINPUT125), .B(n1025), .ZN(n1026) );
  NOR2_X1 U1110 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1111 ( .A1(n1028), .A2(G11), .ZN(n1029) );
  XNOR2_X1 U1112 ( .A(n1029), .B(KEYINPUT126), .ZN(n1030) );
  XNOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1030), .ZN(G150) );
  INV_X1 U1114 ( .A(G150), .ZN(G311) );
endmodule

