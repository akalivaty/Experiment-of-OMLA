

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U558 ( .A1(n707), .A2(n540), .ZN(n754) );
  AND2_X1 U559 ( .A1(G2105), .A2(G2104), .ZN(n897) );
  XOR2_X2 U560 ( .A(n742), .B(KEYINPUT29), .Z(n524) );
  NOR2_X1 U561 ( .A1(G164), .A2(G1384), .ZN(n706) );
  OR2_X1 U562 ( .A1(n581), .A2(n580), .ZN(n583) );
  INV_X8 U563 ( .A(G2105), .ZN(n551) );
  NOR2_X1 U564 ( .A1(n791), .A2(n790), .ZN(n530) );
  NOR2_X1 U565 ( .A1(n738), .A2(G299), .ZN(n721) );
  NOR2_X1 U566 ( .A1(n786), .A2(G1966), .ZN(n747) );
  INV_X2 U567 ( .A(n754), .ZN(n722) );
  XNOR2_X1 U568 ( .A(n706), .B(KEYINPUT64), .ZN(n540) );
  XNOR2_X1 U569 ( .A(n539), .B(n538), .ZN(n537) );
  AND2_X1 U570 ( .A1(G138), .A2(n894), .ZN(n581) );
  XNOR2_X2 U571 ( .A(n583), .B(n582), .ZN(G164) );
  NOR2_X1 U572 ( .A1(n939), .A2(n724), .ZN(n725) );
  XNOR2_X1 U573 ( .A(n553), .B(KEYINPUT26), .ZN(n552) );
  NAND2_X1 U574 ( .A1(n541), .A2(n535), .ZN(n534) );
  INV_X1 U575 ( .A(n746), .ZN(n535) );
  NAND2_X1 U576 ( .A1(n524), .A2(n542), .ZN(n541) );
  INV_X1 U577 ( .A(n745), .ZN(n542) );
  NAND2_X1 U578 ( .A1(n746), .A2(n544), .ZN(n543) );
  INV_X1 U579 ( .A(n747), .ZN(n544) );
  NAND2_X1 U580 ( .A1(n754), .A2(G8), .ZN(n786) );
  NAND2_X1 U581 ( .A1(n533), .A2(n531), .ZN(n711) );
  INV_X1 U582 ( .A(n748), .ZN(n533) );
  NOR2_X1 U583 ( .A1(n747), .A2(n532), .ZN(n531) );
  NAND2_X1 U584 ( .A1(n753), .A2(n534), .ZN(n760) );
  XNOR2_X1 U585 ( .A(n547), .B(KEYINPUT96), .ZN(n750) );
  NAND2_X1 U586 ( .A1(n551), .A2(n550), .ZN(n549) );
  INV_X1 U587 ( .A(G2104), .ZN(n550) );
  INV_X1 U588 ( .A(KEYINPUT102), .ZN(n548) );
  INV_X1 U589 ( .A(KEYINPUT23), .ZN(n538) );
  NAND2_X1 U590 ( .A1(n893), .A2(G101), .ZN(n539) );
  NOR2_X1 U591 ( .A1(n567), .A2(n536), .ZN(G160) );
  AND2_X1 U592 ( .A1(n947), .A2(n839), .ZN(n526) );
  NOR2_X1 U593 ( .A1(n825), .A2(n526), .ZN(n527) );
  INV_X1 U594 ( .A(G8), .ZN(n532) );
  NAND2_X1 U595 ( .A1(n528), .A2(n841), .ZN(n842) );
  NAND2_X1 U596 ( .A1(n529), .A2(n527), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n530), .B(n548), .ZN(n529) );
  NAND2_X1 U598 ( .A1(n537), .A2(n564), .ZN(n536) );
  NOR2_X1 U599 ( .A1(n793), .A2(n540), .ZN(n839) );
  NAND2_X1 U600 ( .A1(n545), .A2(n543), .ZN(n547) );
  NAND2_X1 U601 ( .A1(n524), .A2(n546), .ZN(n545) );
  NOR2_X1 U602 ( .A1(n745), .A2(n747), .ZN(n546) );
  XNOR2_X2 U603 ( .A(n549), .B(KEYINPUT17), .ZN(n894) );
  NAND2_X1 U604 ( .A1(n552), .A2(n723), .ZN(n724) );
  NAND2_X1 U605 ( .A1(n722), .A2(G1996), .ZN(n553) );
  OR2_X1 U606 ( .A1(n722), .A2(n938), .ZN(n554) );
  INV_X1 U607 ( .A(KEYINPUT27), .ZN(n716) );
  XNOR2_X1 U608 ( .A(n717), .B(n716), .ZN(n719) );
  XNOR2_X1 U609 ( .A(KEYINPUT32), .B(KEYINPUT98), .ZN(n761) );
  XNOR2_X1 U610 ( .A(n762), .B(n761), .ZN(n763) );
  NOR2_X1 U611 ( .A1(G651), .A2(n670), .ZN(n671) );
  INV_X1 U612 ( .A(G651), .ZN(n559) );
  NOR2_X1 U613 ( .A1(G543), .A2(n559), .ZN(n556) );
  XNOR2_X1 U614 ( .A(KEYINPUT1), .B(KEYINPUT65), .ZN(n555) );
  XNOR2_X1 U615 ( .A(n556), .B(n555), .ZN(n675) );
  NAND2_X1 U616 ( .A1(G65), .A2(n675), .ZN(n558) );
  NOR2_X1 U617 ( .A1(G651), .A2(G543), .ZN(n661) );
  NAND2_X1 U618 ( .A1(G91), .A2(n661), .ZN(n557) );
  NAND2_X1 U619 ( .A1(n558), .A2(n557), .ZN(n563) );
  XOR2_X1 U620 ( .A(KEYINPUT0), .B(G543), .Z(n670) );
  NOR2_X1 U621 ( .A1(n670), .A2(n559), .ZN(n664) );
  NAND2_X1 U622 ( .A1(G78), .A2(n664), .ZN(n561) );
  NAND2_X1 U623 ( .A1(G53), .A2(n671), .ZN(n560) );
  NAND2_X1 U624 ( .A1(n561), .A2(n560), .ZN(n562) );
  OR2_X1 U625 ( .A1(n563), .A2(n562), .ZN(G299) );
  NAND2_X1 U626 ( .A1(n897), .A2(G113), .ZN(n564) );
  AND2_X2 U627 ( .A1(n551), .A2(G2104), .ZN(n893) );
  NAND2_X1 U628 ( .A1(G137), .A2(n894), .ZN(n566) );
  NOR2_X2 U629 ( .A1(G2104), .A2(n551), .ZN(n898) );
  NAND2_X1 U630 ( .A1(G125), .A2(n898), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U632 ( .A1(G64), .A2(n675), .ZN(n569) );
  NAND2_X1 U633 ( .A1(G52), .A2(n671), .ZN(n568) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(KEYINPUT66), .B(n570), .ZN(n575) );
  NAND2_X1 U636 ( .A1(G90), .A2(n661), .ZN(n572) );
  NAND2_X1 U637 ( .A1(G77), .A2(n664), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U639 ( .A(KEYINPUT9), .B(n573), .Z(n574) );
  NOR2_X1 U640 ( .A1(n575), .A2(n574), .ZN(G171) );
  AND2_X1 U641 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U642 ( .A(G69), .ZN(G235) );
  INV_X1 U643 ( .A(G120), .ZN(G236) );
  INV_X1 U644 ( .A(G132), .ZN(G219) );
  INV_X1 U645 ( .A(G82), .ZN(G220) );
  NAND2_X1 U646 ( .A1(G126), .A2(n898), .ZN(n579) );
  NAND2_X1 U647 ( .A1(G102), .A2(n893), .ZN(n577) );
  NAND2_X1 U648 ( .A1(G114), .A2(n897), .ZN(n576) );
  AND2_X1 U649 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U650 ( .A1(n579), .A2(n578), .ZN(n580) );
  INV_X1 U651 ( .A(KEYINPUT82), .ZN(n582) );
  NAND2_X1 U652 ( .A1(G63), .A2(n675), .ZN(n585) );
  NAND2_X1 U653 ( .A1(G51), .A2(n671), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U655 ( .A(KEYINPUT6), .B(n586), .ZN(n594) );
  NAND2_X1 U656 ( .A1(n664), .A2(G76), .ZN(n587) );
  XNOR2_X1 U657 ( .A(KEYINPUT70), .B(n587), .ZN(n591) );
  XOR2_X1 U658 ( .A(KEYINPUT69), .B(KEYINPUT4), .Z(n589) );
  NAND2_X1 U659 ( .A1(G89), .A2(n661), .ZN(n588) );
  XNOR2_X1 U660 ( .A(n589), .B(n588), .ZN(n590) );
  NAND2_X1 U661 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U662 ( .A(n592), .B(KEYINPUT5), .Z(n593) );
  NOR2_X1 U663 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U664 ( .A(KEYINPUT71), .B(n595), .Z(n596) );
  XOR2_X1 U665 ( .A(KEYINPUT7), .B(n596), .Z(G168) );
  XOR2_X1 U666 ( .A(G168), .B(KEYINPUT8), .Z(n597) );
  XNOR2_X1 U667 ( .A(KEYINPUT72), .B(n597), .ZN(G286) );
  NAND2_X1 U668 ( .A1(G7), .A2(G661), .ZN(n598) );
  XNOR2_X1 U669 ( .A(n598), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U670 ( .A(G223), .ZN(n843) );
  NAND2_X1 U671 ( .A1(n843), .A2(G567), .ZN(n599) );
  XOR2_X1 U672 ( .A(KEYINPUT11), .B(n599), .Z(G234) );
  NAND2_X1 U673 ( .A1(G56), .A2(n675), .ZN(n600) );
  XOR2_X1 U674 ( .A(KEYINPUT14), .B(n600), .Z(n606) );
  NAND2_X1 U675 ( .A1(n661), .A2(G81), .ZN(n601) );
  XNOR2_X1 U676 ( .A(n601), .B(KEYINPUT12), .ZN(n603) );
  NAND2_X1 U677 ( .A1(G68), .A2(n664), .ZN(n602) );
  NAND2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U679 ( .A(KEYINPUT13), .B(n604), .Z(n605) );
  NOR2_X1 U680 ( .A1(n606), .A2(n605), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n671), .A2(G43), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n608), .A2(n607), .ZN(n939) );
  INV_X1 U683 ( .A(n939), .ZN(n679) );
  NAND2_X1 U684 ( .A1(n679), .A2(G860), .ZN(G153) );
  XOR2_X1 U685 ( .A(G171), .B(KEYINPUT68), .Z(G301) );
  NAND2_X1 U686 ( .A1(G868), .A2(G301), .ZN(n617) );
  NAND2_X1 U687 ( .A1(G66), .A2(n675), .ZN(n610) );
  NAND2_X1 U688 ( .A1(G92), .A2(n661), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n614) );
  NAND2_X1 U690 ( .A1(G79), .A2(n664), .ZN(n612) );
  NAND2_X1 U691 ( .A1(G54), .A2(n671), .ZN(n611) );
  NAND2_X1 U692 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U693 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U694 ( .A(KEYINPUT15), .B(n615), .Z(n937) );
  OR2_X1 U695 ( .A1(n937), .A2(G868), .ZN(n616) );
  NAND2_X1 U696 ( .A1(n617), .A2(n616), .ZN(G284) );
  INV_X1 U697 ( .A(G868), .ZN(n688) );
  NAND2_X1 U698 ( .A1(G299), .A2(n688), .ZN(n619) );
  NAND2_X1 U699 ( .A1(G868), .A2(G286), .ZN(n618) );
  NAND2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U701 ( .A(KEYINPUT73), .B(n620), .Z(G297) );
  INV_X1 U702 ( .A(G860), .ZN(n621) );
  NAND2_X1 U703 ( .A1(n621), .A2(G559), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n622), .A2(n937), .ZN(n623) );
  XNOR2_X1 U705 ( .A(n623), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U706 ( .A1(G868), .A2(n939), .ZN(n626) );
  NAND2_X1 U707 ( .A1(G868), .A2(n937), .ZN(n624) );
  NOR2_X1 U708 ( .A1(G559), .A2(n624), .ZN(n625) );
  NOR2_X1 U709 ( .A1(n626), .A2(n625), .ZN(G282) );
  NAND2_X1 U710 ( .A1(G123), .A2(n898), .ZN(n627) );
  XNOR2_X1 U711 ( .A(n627), .B(KEYINPUT18), .ZN(n634) );
  NAND2_X1 U712 ( .A1(G111), .A2(n897), .ZN(n629) );
  NAND2_X1 U713 ( .A1(G135), .A2(n894), .ZN(n628) );
  NAND2_X1 U714 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n893), .A2(G99), .ZN(n630) );
  XOR2_X1 U716 ( .A(KEYINPUT74), .B(n630), .Z(n631) );
  NOR2_X1 U717 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U718 ( .A1(n634), .A2(n633), .ZN(n1016) );
  XOR2_X1 U719 ( .A(G2096), .B(KEYINPUT75), .Z(n635) );
  XNOR2_X1 U720 ( .A(n1016), .B(n635), .ZN(n636) );
  NOR2_X1 U721 ( .A1(G2100), .A2(n636), .ZN(n637) );
  XOR2_X1 U722 ( .A(KEYINPUT76), .B(n637), .Z(G156) );
  NAND2_X1 U723 ( .A1(G93), .A2(n661), .ZN(n639) );
  NAND2_X1 U724 ( .A1(G80), .A2(n664), .ZN(n638) );
  NAND2_X1 U725 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U726 ( .A(KEYINPUT78), .B(n640), .ZN(n644) );
  NAND2_X1 U727 ( .A1(G67), .A2(n675), .ZN(n642) );
  NAND2_X1 U728 ( .A1(G55), .A2(n671), .ZN(n641) );
  NAND2_X1 U729 ( .A1(n642), .A2(n641), .ZN(n643) );
  OR2_X1 U730 ( .A1(n644), .A2(n643), .ZN(n689) );
  NAND2_X1 U731 ( .A1(n937), .A2(G559), .ZN(n686) );
  XOR2_X1 U732 ( .A(KEYINPUT77), .B(n939), .Z(n645) );
  XNOR2_X1 U733 ( .A(n686), .B(n645), .ZN(n646) );
  NOR2_X1 U734 ( .A1(G860), .A2(n646), .ZN(n647) );
  XOR2_X1 U735 ( .A(n689), .B(n647), .Z(G145) );
  AND2_X1 U736 ( .A1(n675), .A2(G60), .ZN(n651) );
  NAND2_X1 U737 ( .A1(G85), .A2(n661), .ZN(n649) );
  NAND2_X1 U738 ( .A1(G72), .A2(n664), .ZN(n648) );
  NAND2_X1 U739 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U740 ( .A1(n651), .A2(n650), .ZN(n653) );
  NAND2_X1 U741 ( .A1(n671), .A2(G47), .ZN(n652) );
  NAND2_X1 U742 ( .A1(n653), .A2(n652), .ZN(G290) );
  NAND2_X1 U743 ( .A1(G62), .A2(n675), .ZN(n655) );
  NAND2_X1 U744 ( .A1(G88), .A2(n661), .ZN(n654) );
  NAND2_X1 U745 ( .A1(n655), .A2(n654), .ZN(n658) );
  NAND2_X1 U746 ( .A1(n664), .A2(G75), .ZN(n656) );
  XOR2_X1 U747 ( .A(KEYINPUT80), .B(n656), .Z(n657) );
  NOR2_X1 U748 ( .A1(n658), .A2(n657), .ZN(n660) );
  NAND2_X1 U749 ( .A1(n671), .A2(G50), .ZN(n659) );
  NAND2_X1 U750 ( .A1(n660), .A2(n659), .ZN(G303) );
  INV_X1 U751 ( .A(G303), .ZN(G166) );
  NAND2_X1 U752 ( .A1(G61), .A2(n675), .ZN(n663) );
  NAND2_X1 U753 ( .A1(G86), .A2(n661), .ZN(n662) );
  NAND2_X1 U754 ( .A1(n663), .A2(n662), .ZN(n667) );
  NAND2_X1 U755 ( .A1(n664), .A2(G73), .ZN(n665) );
  XOR2_X1 U756 ( .A(KEYINPUT2), .B(n665), .Z(n666) );
  NOR2_X1 U757 ( .A1(n667), .A2(n666), .ZN(n669) );
  NAND2_X1 U758 ( .A1(n671), .A2(G48), .ZN(n668) );
  NAND2_X1 U759 ( .A1(n669), .A2(n668), .ZN(G305) );
  NAND2_X1 U760 ( .A1(n670), .A2(G87), .ZN(n677) );
  NAND2_X1 U761 ( .A1(G49), .A2(n671), .ZN(n673) );
  NAND2_X1 U762 ( .A1(G74), .A2(G651), .ZN(n672) );
  NAND2_X1 U763 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U764 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U765 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U766 ( .A(KEYINPUT79), .B(n678), .Z(G288) );
  XNOR2_X1 U767 ( .A(KEYINPUT19), .B(G290), .ZN(n685) );
  XNOR2_X1 U768 ( .A(n689), .B(n679), .ZN(n680) );
  XNOR2_X1 U769 ( .A(n680), .B(G305), .ZN(n681) );
  XNOR2_X1 U770 ( .A(n681), .B(G288), .ZN(n682) );
  XNOR2_X1 U771 ( .A(G166), .B(n682), .ZN(n683) );
  XNOR2_X1 U772 ( .A(n683), .B(G299), .ZN(n684) );
  XNOR2_X1 U773 ( .A(n685), .B(n684), .ZN(n914) );
  XOR2_X1 U774 ( .A(n914), .B(n686), .Z(n687) );
  NAND2_X1 U775 ( .A1(G868), .A2(n687), .ZN(n691) );
  NAND2_X1 U776 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U777 ( .A1(n691), .A2(n690), .ZN(G295) );
  NAND2_X1 U778 ( .A1(G2078), .A2(G2084), .ZN(n692) );
  XOR2_X1 U779 ( .A(KEYINPUT20), .B(n692), .Z(n693) );
  NAND2_X1 U780 ( .A1(G2090), .A2(n693), .ZN(n694) );
  XNOR2_X1 U781 ( .A(KEYINPUT21), .B(n694), .ZN(n695) );
  NAND2_X1 U782 ( .A1(n695), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U783 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U784 ( .A(KEYINPUT67), .B(G57), .ZN(G237) );
  NOR2_X1 U785 ( .A1(G220), .A2(G219), .ZN(n696) );
  XOR2_X1 U786 ( .A(KEYINPUT22), .B(n696), .Z(n697) );
  NOR2_X1 U787 ( .A1(G218), .A2(n697), .ZN(n698) );
  NAND2_X1 U788 ( .A1(G96), .A2(n698), .ZN(n847) );
  NAND2_X1 U789 ( .A1(n847), .A2(G2106), .ZN(n703) );
  NOR2_X1 U790 ( .A1(G237), .A2(G236), .ZN(n699) );
  NAND2_X1 U791 ( .A1(G108), .A2(n699), .ZN(n700) );
  NOR2_X1 U792 ( .A1(n700), .A2(G235), .ZN(n701) );
  XNOR2_X1 U793 ( .A(n701), .B(KEYINPUT81), .ZN(n848) );
  NAND2_X1 U794 ( .A1(n848), .A2(G567), .ZN(n702) );
  NAND2_X1 U795 ( .A1(n703), .A2(n702), .ZN(n849) );
  NAND2_X1 U796 ( .A1(G661), .A2(G483), .ZN(n704) );
  NOR2_X1 U797 ( .A1(n849), .A2(n704), .ZN(n846) );
  NAND2_X1 U798 ( .A1(n846), .A2(G36), .ZN(G176) );
  NAND2_X1 U799 ( .A1(G40), .A2(G160), .ZN(n792) );
  XNOR2_X1 U800 ( .A(KEYINPUT83), .B(n792), .ZN(n707) );
  NOR2_X1 U801 ( .A1(n722), .A2(G1961), .ZN(n708) );
  XOR2_X1 U802 ( .A(KEYINPUT90), .B(n708), .Z(n710) );
  XNOR2_X1 U803 ( .A(G2078), .B(KEYINPUT25), .ZN(n990) );
  NAND2_X1 U804 ( .A1(n722), .A2(n990), .ZN(n709) );
  NAND2_X1 U805 ( .A1(n710), .A2(n709), .ZN(n743) );
  NOR2_X1 U806 ( .A1(G171), .A2(n743), .ZN(n714) );
  NOR2_X1 U807 ( .A1(G2084), .A2(n754), .ZN(n748) );
  XNOR2_X1 U808 ( .A(KEYINPUT30), .B(n711), .ZN(n712) );
  NOR2_X1 U809 ( .A1(G168), .A2(n712), .ZN(n713) );
  NOR2_X1 U810 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U811 ( .A(n715), .B(KEYINPUT31), .ZN(n746) );
  NAND2_X1 U812 ( .A1(n722), .A2(G2072), .ZN(n717) );
  NAND2_X1 U813 ( .A1(n754), .A2(G1956), .ZN(n718) );
  NAND2_X1 U814 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U815 ( .A(n720), .B(KEYINPUT92), .ZN(n738) );
  XNOR2_X1 U816 ( .A(n721), .B(KEYINPUT95), .ZN(n737) );
  NAND2_X1 U817 ( .A1(n754), .A2(G1341), .ZN(n723) );
  OR2_X1 U818 ( .A1(n937), .A2(n725), .ZN(n735) );
  NAND2_X1 U819 ( .A1(n937), .A2(n725), .ZN(n733) );
  NAND2_X1 U820 ( .A1(G2067), .A2(n722), .ZN(n726) );
  XNOR2_X1 U821 ( .A(KEYINPUT94), .B(n726), .ZN(n727) );
  INV_X1 U822 ( .A(G1348), .ZN(n938) );
  NAND2_X1 U823 ( .A1(n727), .A2(n554), .ZN(n728) );
  NOR2_X1 U824 ( .A1(KEYINPUT93), .A2(n728), .ZN(n731) );
  NAND2_X1 U825 ( .A1(KEYINPUT94), .A2(KEYINPUT93), .ZN(n729) );
  NOR2_X1 U826 ( .A1(n729), .A2(n554), .ZN(n730) );
  NOR2_X1 U827 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U828 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U829 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U830 ( .A1(n737), .A2(n736), .ZN(n741) );
  NAND2_X1 U831 ( .A1(n738), .A2(G299), .ZN(n739) );
  XNOR2_X1 U832 ( .A(n739), .B(KEYINPUT28), .ZN(n740) );
  NAND2_X1 U833 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U834 ( .A1(G171), .A2(n743), .ZN(n744) );
  XNOR2_X1 U835 ( .A(KEYINPUT91), .B(n744), .ZN(n745) );
  NAND2_X1 U836 ( .A1(G8), .A2(n748), .ZN(n749) );
  NAND2_X1 U837 ( .A1(n750), .A2(n749), .ZN(n752) );
  INV_X1 U838 ( .A(KEYINPUT97), .ZN(n751) );
  XNOR2_X1 U839 ( .A(n752), .B(n751), .ZN(n764) );
  AND2_X1 U840 ( .A1(G286), .A2(G8), .ZN(n753) );
  NOR2_X1 U841 ( .A1(G2090), .A2(n754), .ZN(n756) );
  NOR2_X1 U842 ( .A1(G1971), .A2(n786), .ZN(n755) );
  NOR2_X1 U843 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U844 ( .A1(n757), .A2(G303), .ZN(n758) );
  OR2_X1 U845 ( .A1(n532), .A2(n758), .ZN(n759) );
  AND2_X1 U846 ( .A1(n760), .A2(n759), .ZN(n762) );
  NAND2_X1 U847 ( .A1(n764), .A2(n763), .ZN(n783) );
  NOR2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n950) );
  NOR2_X1 U849 ( .A1(G1971), .A2(G303), .ZN(n765) );
  NOR2_X1 U850 ( .A1(n950), .A2(n765), .ZN(n766) );
  XOR2_X1 U851 ( .A(KEYINPUT99), .B(n766), .Z(n768) );
  INV_X1 U852 ( .A(KEYINPUT33), .ZN(n767) );
  AND2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U854 ( .A1(n783), .A2(n769), .ZN(n773) );
  INV_X1 U855 ( .A(n786), .ZN(n770) );
  NAND2_X1 U856 ( .A1(G1976), .A2(G288), .ZN(n951) );
  AND2_X1 U857 ( .A1(n770), .A2(n951), .ZN(n771) );
  OR2_X1 U858 ( .A1(KEYINPUT33), .A2(n771), .ZN(n772) );
  NAND2_X1 U859 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U860 ( .A(n774), .B(KEYINPUT100), .ZN(n779) );
  XOR2_X1 U861 ( .A(G1981), .B(G305), .Z(n934) );
  NAND2_X1 U862 ( .A1(n950), .A2(KEYINPUT33), .ZN(n775) );
  NOR2_X1 U863 ( .A1(n786), .A2(n775), .ZN(n776) );
  XNOR2_X1 U864 ( .A(n776), .B(KEYINPUT101), .ZN(n777) );
  NAND2_X1 U865 ( .A1(n934), .A2(n777), .ZN(n778) );
  NOR2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n791) );
  NOR2_X1 U867 ( .A1(G1981), .A2(G305), .ZN(n780) );
  XOR2_X1 U868 ( .A(n780), .B(KEYINPUT24), .Z(n781) );
  NOR2_X1 U869 ( .A1(n786), .A2(n781), .ZN(n782) );
  XNOR2_X1 U870 ( .A(n782), .B(KEYINPUT89), .ZN(n789) );
  NOR2_X1 U871 ( .A1(G2090), .A2(G303), .ZN(n784) );
  NAND2_X1 U872 ( .A1(G8), .A2(n784), .ZN(n785) );
  NAND2_X1 U873 ( .A1(n783), .A2(n785), .ZN(n787) );
  NAND2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U876 ( .A(KEYINPUT83), .B(n792), .Z(n793) );
  XOR2_X1 U877 ( .A(KEYINPUT36), .B(KEYINPUT86), .Z(n805) );
  XNOR2_X1 U878 ( .A(KEYINPUT34), .B(KEYINPUT84), .ZN(n797) );
  NAND2_X1 U879 ( .A1(G104), .A2(n893), .ZN(n795) );
  NAND2_X1 U880 ( .A1(G140), .A2(n894), .ZN(n794) );
  NAND2_X1 U881 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U882 ( .A(n797), .B(n796), .ZN(n802) );
  NAND2_X1 U883 ( .A1(G116), .A2(n897), .ZN(n799) );
  NAND2_X1 U884 ( .A1(G128), .A2(n898), .ZN(n798) );
  NAND2_X1 U885 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U886 ( .A(KEYINPUT35), .B(n800), .Z(n801) );
  NOR2_X1 U887 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U888 ( .A(n803), .B(KEYINPUT85), .ZN(n804) );
  XNOR2_X1 U889 ( .A(n805), .B(n804), .ZN(n912) );
  XNOR2_X1 U890 ( .A(KEYINPUT37), .B(G2067), .ZN(n837) );
  NOR2_X1 U891 ( .A1(n912), .A2(n837), .ZN(n1022) );
  NAND2_X1 U892 ( .A1(n839), .A2(n1022), .ZN(n834) );
  NAND2_X1 U893 ( .A1(G95), .A2(n893), .ZN(n807) );
  NAND2_X1 U894 ( .A1(G131), .A2(n894), .ZN(n806) );
  NAND2_X1 U895 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U896 ( .A(KEYINPUT88), .B(n808), .ZN(n811) );
  NAND2_X1 U897 ( .A1(G107), .A2(n897), .ZN(n809) );
  XNOR2_X1 U898 ( .A(KEYINPUT87), .B(n809), .ZN(n810) );
  NOR2_X1 U899 ( .A1(n811), .A2(n810), .ZN(n813) );
  NAND2_X1 U900 ( .A1(n898), .A2(G119), .ZN(n812) );
  NAND2_X1 U901 ( .A1(n813), .A2(n812), .ZN(n906) );
  AND2_X1 U902 ( .A1(n906), .A2(G1991), .ZN(n822) );
  NAND2_X1 U903 ( .A1(G117), .A2(n897), .ZN(n815) );
  NAND2_X1 U904 ( .A1(G141), .A2(n894), .ZN(n814) );
  NAND2_X1 U905 ( .A1(n815), .A2(n814), .ZN(n818) );
  NAND2_X1 U906 ( .A1(n893), .A2(G105), .ZN(n816) );
  XOR2_X1 U907 ( .A(KEYINPUT38), .B(n816), .Z(n817) );
  NOR2_X1 U908 ( .A1(n818), .A2(n817), .ZN(n820) );
  NAND2_X1 U909 ( .A1(n898), .A2(G129), .ZN(n819) );
  NAND2_X1 U910 ( .A1(n820), .A2(n819), .ZN(n908) );
  AND2_X1 U911 ( .A1(G1996), .A2(n908), .ZN(n821) );
  NOR2_X1 U912 ( .A1(n822), .A2(n821), .ZN(n1021) );
  INV_X1 U913 ( .A(n839), .ZN(n823) );
  NOR2_X1 U914 ( .A1(n1021), .A2(n823), .ZN(n829) );
  INV_X1 U915 ( .A(n829), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n834), .A2(n824), .ZN(n825) );
  XNOR2_X1 U917 ( .A(G1986), .B(G290), .ZN(n947) );
  XOR2_X1 U918 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n833) );
  NOR2_X1 U919 ( .A1(G1996), .A2(n908), .ZN(n826) );
  XOR2_X1 U920 ( .A(KEYINPUT103), .B(n826), .Z(n1028) );
  NOR2_X1 U921 ( .A1(G1991), .A2(n906), .ZN(n1019) );
  NOR2_X1 U922 ( .A1(G1986), .A2(G290), .ZN(n827) );
  NOR2_X1 U923 ( .A1(n1019), .A2(n827), .ZN(n828) );
  NOR2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n830) );
  NOR2_X1 U925 ( .A1(n1028), .A2(n830), .ZN(n831) );
  XNOR2_X1 U926 ( .A(n831), .B(KEYINPUT39), .ZN(n832) );
  XNOR2_X1 U927 ( .A(n833), .B(n832), .ZN(n835) );
  NAND2_X1 U928 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U929 ( .A(n836), .B(KEYINPUT106), .ZN(n838) );
  NAND2_X1 U930 ( .A1(n912), .A2(n837), .ZN(n1026) );
  NAND2_X1 U931 ( .A1(n838), .A2(n1026), .ZN(n840) );
  NAND2_X1 U932 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U933 ( .A(KEYINPUT40), .B(n842), .ZN(G329) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n843), .ZN(G217) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n844) );
  NAND2_X1 U936 ( .A1(G661), .A2(n844), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n845) );
  NAND2_X1 U938 ( .A1(n846), .A2(n845), .ZN(G188) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  NOR2_X1 U941 ( .A1(n848), .A2(n847), .ZN(G325) );
  INV_X1 U942 ( .A(G325), .ZN(G261) );
  INV_X1 U943 ( .A(n849), .ZN(G319) );
  XOR2_X1 U944 ( .A(KEYINPUT110), .B(G1956), .Z(n851) );
  XNOR2_X1 U945 ( .A(G1986), .B(G1976), .ZN(n850) );
  XNOR2_X1 U946 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U947 ( .A(n852), .B(KEYINPUT41), .Z(n854) );
  XNOR2_X1 U948 ( .A(G1996), .B(G1991), .ZN(n853) );
  XNOR2_X1 U949 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U950 ( .A(G1966), .B(G1961), .Z(n856) );
  XNOR2_X1 U951 ( .A(G1981), .B(G1971), .ZN(n855) );
  XNOR2_X1 U952 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U953 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U954 ( .A(KEYINPUT109), .B(G2474), .ZN(n859) );
  XNOR2_X1 U955 ( .A(n860), .B(n859), .ZN(G229) );
  XOR2_X1 U956 ( .A(KEYINPUT43), .B(G2678), .Z(n862) );
  XNOR2_X1 U957 ( .A(KEYINPUT108), .B(KEYINPUT107), .ZN(n861) );
  XNOR2_X1 U958 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U959 ( .A(KEYINPUT42), .B(G2072), .Z(n864) );
  XNOR2_X1 U960 ( .A(G2067), .B(G2090), .ZN(n863) );
  XNOR2_X1 U961 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U962 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U963 ( .A(G2096), .B(G2100), .ZN(n867) );
  XNOR2_X1 U964 ( .A(n868), .B(n867), .ZN(n870) );
  XOR2_X1 U965 ( .A(G2078), .B(G2084), .Z(n869) );
  XNOR2_X1 U966 ( .A(n870), .B(n869), .ZN(G227) );
  NAND2_X1 U967 ( .A1(G100), .A2(n893), .ZN(n871) );
  XNOR2_X1 U968 ( .A(n871), .B(KEYINPUT112), .ZN(n874) );
  NAND2_X1 U969 ( .A1(G112), .A2(n897), .ZN(n872) );
  XOR2_X1 U970 ( .A(KEYINPUT111), .B(n872), .Z(n873) );
  NAND2_X1 U971 ( .A1(n874), .A2(n873), .ZN(n879) );
  NAND2_X1 U972 ( .A1(G124), .A2(n898), .ZN(n875) );
  XNOR2_X1 U973 ( .A(n875), .B(KEYINPUT44), .ZN(n877) );
  NAND2_X1 U974 ( .A1(n894), .A2(G136), .ZN(n876) );
  NAND2_X1 U975 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U976 ( .A1(n879), .A2(n878), .ZN(G162) );
  NAND2_X1 U977 ( .A1(G118), .A2(n897), .ZN(n881) );
  NAND2_X1 U978 ( .A1(G130), .A2(n898), .ZN(n880) );
  NAND2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n886) );
  NAND2_X1 U980 ( .A1(G106), .A2(n893), .ZN(n883) );
  NAND2_X1 U981 ( .A1(G142), .A2(n894), .ZN(n882) );
  NAND2_X1 U982 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U983 ( .A(KEYINPUT45), .B(n884), .Z(n885) );
  NOR2_X1 U984 ( .A1(n886), .A2(n885), .ZN(n892) );
  XOR2_X1 U985 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n887) );
  XNOR2_X1 U986 ( .A(n1016), .B(n887), .ZN(n888) );
  XNOR2_X1 U987 ( .A(KEYINPUT114), .B(n888), .ZN(n890) );
  XNOR2_X1 U988 ( .A(G164), .B(KEYINPUT48), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U990 ( .A(n892), .B(n891), .Z(n905) );
  NAND2_X1 U991 ( .A1(G103), .A2(n893), .ZN(n896) );
  NAND2_X1 U992 ( .A1(G139), .A2(n894), .ZN(n895) );
  NAND2_X1 U993 ( .A1(n896), .A2(n895), .ZN(n903) );
  NAND2_X1 U994 ( .A1(G115), .A2(n897), .ZN(n900) );
  NAND2_X1 U995 ( .A1(G127), .A2(n898), .ZN(n899) );
  NAND2_X1 U996 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U997 ( .A(KEYINPUT47), .B(n901), .Z(n902) );
  NOR2_X1 U998 ( .A1(n903), .A2(n902), .ZN(n1012) );
  XNOR2_X1 U999 ( .A(G162), .B(n1012), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(n905), .B(n904), .ZN(n907) );
  XNOR2_X1 U1001 ( .A(n907), .B(n906), .ZN(n910) );
  XOR2_X1 U1002 ( .A(G160), .B(n908), .Z(n909) );
  XNOR2_X1 U1003 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1004 ( .A(n912), .B(n911), .Z(n913) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n913), .ZN(G395) );
  XNOR2_X1 U1006 ( .A(n937), .B(n914), .ZN(n916) );
  XNOR2_X1 U1007 ( .A(G286), .B(G171), .ZN(n915) );
  XNOR2_X1 U1008 ( .A(n916), .B(n915), .ZN(n917) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n917), .ZN(G397) );
  XOR2_X1 U1010 ( .A(G2451), .B(G2430), .Z(n919) );
  XNOR2_X1 U1011 ( .A(G2438), .B(G2443), .ZN(n918) );
  XNOR2_X1 U1012 ( .A(n919), .B(n918), .ZN(n925) );
  XOR2_X1 U1013 ( .A(G2435), .B(G2454), .Z(n921) );
  XNOR2_X1 U1014 ( .A(G1348), .B(G1341), .ZN(n920) );
  XNOR2_X1 U1015 ( .A(n921), .B(n920), .ZN(n923) );
  XOR2_X1 U1016 ( .A(G2446), .B(G2427), .Z(n922) );
  XNOR2_X1 U1017 ( .A(n923), .B(n922), .ZN(n924) );
  XOR2_X1 U1018 ( .A(n925), .B(n924), .Z(n926) );
  NAND2_X1 U1019 ( .A1(G14), .A2(n926), .ZN(n932) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n932), .ZN(n929) );
  NOR2_X1 U1021 ( .A1(G229), .A2(G227), .ZN(n927) );
  XNOR2_X1 U1022 ( .A(KEYINPUT49), .B(n927), .ZN(n928) );
  NOR2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(n931) );
  NOR2_X1 U1024 ( .A1(G395), .A2(G397), .ZN(n930) );
  NAND2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(G225) );
  INV_X1 U1026 ( .A(G225), .ZN(G308) );
  INV_X1 U1027 ( .A(G108), .ZN(G238) );
  INV_X1 U1028 ( .A(n932), .ZN(G401) );
  XNOR2_X1 U1029 ( .A(KEYINPUT56), .B(G16), .ZN(n959) );
  XOR2_X1 U1030 ( .A(G168), .B(G1966), .Z(n933) );
  XNOR2_X1 U1031 ( .A(KEYINPUT121), .B(n933), .ZN(n935) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(n936), .B(KEYINPUT57), .ZN(n957) );
  XNOR2_X1 U1034 ( .A(n938), .B(n937), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(n939), .B(G1341), .ZN(n940) );
  NOR2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n949) );
  XNOR2_X1 U1037 ( .A(G171), .B(G1961), .ZN(n945) );
  XNOR2_X1 U1038 ( .A(G303), .B(G1971), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(G299), .B(G1956), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n955) );
  INV_X1 U1044 ( .A(n950), .ZN(n952) );
  NAND2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(KEYINPUT122), .B(n953), .ZN(n954) );
  NOR2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1048 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1049 ( .A1(n959), .A2(n958), .ZN(n987) );
  XNOR2_X1 U1050 ( .A(G16), .B(KEYINPUT123), .ZN(n985) );
  XOR2_X1 U1051 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n983) );
  XNOR2_X1 U1052 ( .A(KEYINPUT125), .B(G1966), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(n960), .B(G21), .ZN(n973) );
  XNOR2_X1 U1054 ( .A(G1348), .B(KEYINPUT59), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(n961), .B(G4), .ZN(n965) );
  XNOR2_X1 U1056 ( .A(G1341), .B(G19), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(G20), .B(G1956), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(KEYINPUT124), .B(G1981), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(G6), .B(n966), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1063 ( .A(KEYINPUT60), .B(n969), .Z(n971) );
  XNOR2_X1 U1064 ( .A(G1961), .B(G5), .ZN(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n980) );
  XNOR2_X1 U1067 ( .A(G1976), .B(G23), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(G1971), .B(G22), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n977) );
  XOR2_X1 U1070 ( .A(G1986), .B(G24), .Z(n976) );
  NAND2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(KEYINPUT58), .B(n978), .ZN(n979) );
  NOR2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(n981), .B(KEYINPUT61), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(n983), .B(n982), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n1011) );
  XOR2_X1 U1078 ( .A(G1991), .B(G25), .Z(n988) );
  NAND2_X1 U1079 ( .A1(n988), .A2(G28), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(n989), .B(KEYINPUT119), .ZN(n998) );
  XNOR2_X1 U1081 ( .A(G27), .B(n990), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(G1996), .B(G32), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(G2072), .B(G33), .ZN(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(G26), .B(G2067), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(n999), .B(KEYINPUT53), .ZN(n1002) );
  XOR2_X1 U1090 ( .A(G2084), .B(G34), .Z(n1000) );
  XNOR2_X1 U1091 ( .A(KEYINPUT54), .B(n1000), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G35), .B(G2090), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(n1005), .B(KEYINPUT55), .ZN(n1007) );
  INV_X1 U1096 ( .A(G29), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(G11), .A2(n1008), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(KEYINPUT120), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1042) );
  INV_X1 U1101 ( .A(KEYINPUT55), .ZN(n1038) );
  XOR2_X1 U1102 ( .A(G2072), .B(n1012), .Z(n1014) );
  XOR2_X1 U1103 ( .A(G164), .B(G2078), .Z(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(KEYINPUT50), .B(n1015), .ZN(n1035) );
  XNOR2_X1 U1106 ( .A(G160), .B(G2084), .ZN(n1017) );
  NAND2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1023) );
  NOR2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1111 ( .A(KEYINPUT115), .B(n1024), .Z(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1033) );
  XOR2_X1 U1113 ( .A(G2090), .B(G162), .Z(n1027) );
  NOR2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1115 ( .A(KEYINPUT51), .B(n1029), .Z(n1031) );
  XNOR2_X1 U1116 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n1030) );
  XNOR2_X1 U1117 ( .A(n1031), .B(n1030), .ZN(n1032) );
  NOR2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1119 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XOR2_X1 U1120 ( .A(KEYINPUT52), .B(n1036), .Z(n1037) );
  NAND2_X1 U1121 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NAND2_X1 U1122 ( .A1(n1039), .A2(G29), .ZN(n1040) );
  XNOR2_X1 U1123 ( .A(n1040), .B(KEYINPUT118), .ZN(n1041) );
  NAND2_X1 U1124 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  XOR2_X1 U1125 ( .A(KEYINPUT62), .B(n1043), .Z(G311) );
  INV_X1 U1126 ( .A(G311), .ZN(G150) );
endmodule

