//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(new_n203), .A2(G50), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G1), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n211), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  OR3_X1    g0016(.A1(new_n216), .A2(KEYINPUT64), .A3(G13), .ZN(new_n217));
  OAI21_X1  g0017(.A(KEYINPUT64), .B1(new_n216), .B2(G13), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT0), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n213), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(new_n221), .B2(new_n220), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT65), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  INV_X1    g0025(.A(G238), .ZN(new_n226));
  INV_X1    g0026(.A(G87), .ZN(new_n227));
  INV_X1    g0027(.A(G250), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n225), .B1(new_n202), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n230));
  INV_X1    g0030(.A(G77), .ZN(new_n231));
  INV_X1    g0031(.A(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G107), .ZN(new_n233));
  INV_X1    g0033(.A(G264), .ZN(new_n234));
  OAI221_X1 g0034(.A(new_n230), .B1(new_n231), .B2(new_n232), .C1(new_n233), .C2(new_n234), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n216), .B1(new_n229), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT1), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n224), .A2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G358));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT67), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G68), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(new_n201), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT66), .B(G50), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n250), .B(new_n254), .ZN(G351));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n210), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n257), .B(KEYINPUT68), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n214), .A2(G13), .A3(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT8), .B(G58), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n211), .A2(G1), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n261), .A2(new_n264), .B1(new_n260), .B2(new_n262), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT73), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT16), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT7), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT3), .B(G33), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n268), .B1(new_n269), .B2(G20), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n274));
  OAI211_X1 g0074(.A(KEYINPUT7), .B(new_n211), .C1(new_n272), .C2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n202), .B1(new_n270), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n211), .A2(new_n273), .A3(KEYINPUT69), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT69), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(G20), .B2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G159), .ZN(new_n281));
  XNOR2_X1  g0081(.A(G58), .B(G68), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n266), .B(new_n267), .C1(new_n276), .C2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n271), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(KEYINPUT7), .B1(new_n288), .B2(new_n211), .ZN(new_n289));
  AOI211_X1 g0089(.A(new_n268), .B(G20), .C1(new_n286), .C2(new_n287), .ZN(new_n290));
  OAI21_X1  g0090(.A(G68), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n281), .A2(new_n283), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(KEYINPUT16), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n285), .A2(new_n293), .A3(new_n257), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(new_n292), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n266), .B1(new_n295), .B2(new_n267), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n265), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G200), .ZN(new_n298));
  INV_X1    g0098(.A(G41), .ZN(new_n299));
  OAI211_X1 g0099(.A(G1), .B(G13), .C1(new_n273), .C2(new_n299), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n286), .A2(new_n287), .A3(G226), .A4(G1698), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT74), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n269), .A2(KEYINPUT74), .A3(G226), .A4(G1698), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G1698), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n286), .A2(new_n287), .A3(G223), .A4(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G33), .A2(G87), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n300), .B1(new_n305), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n312));
  INV_X1    g0112(.A(G274), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n214), .B1(G41), .B2(G45), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n300), .A2(new_n314), .ZN(new_n317));
  INV_X1    g0117(.A(G232), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n298), .B1(new_n311), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n317), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n315), .B1(G232), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G190), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n309), .B1(new_n303), .B2(new_n304), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n322), .B(new_n323), .C1(new_n324), .C2(new_n300), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT17), .B1(new_n297), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT75), .ZN(new_n328));
  INV_X1    g0128(.A(new_n257), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n270), .A2(new_n275), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n284), .B1(G68), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n329), .B1(new_n331), .B2(KEYINPUT16), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n267), .B1(new_n276), .B2(new_n284), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT73), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n334), .A3(new_n285), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n320), .A2(new_n325), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(new_n265), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT75), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT17), .ZN(new_n339));
  INV_X1    g0139(.A(new_n265), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n285), .A2(new_n293), .A3(new_n257), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n340), .B1(new_n341), .B2(new_n334), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT17), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n342), .A2(KEYINPUT76), .A3(new_n343), .A4(new_n336), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n335), .A2(new_n343), .A3(new_n336), .A4(new_n265), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT76), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n328), .A2(new_n339), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n322), .B1(new_n324), .B2(new_n300), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G169), .ZN(new_n350));
  INV_X1    g0150(.A(G179), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n350), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n297), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n353), .B(KEYINPUT18), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  XOR2_X1   g0155(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n269), .A2(G1698), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT71), .B1(new_n358), .B2(new_n318), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT71), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n269), .A2(new_n360), .A3(G232), .A4(G1698), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(G33), .A2(G97), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n269), .A2(new_n306), .ZN(new_n364));
  INV_X1    g0164(.A(G226), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n300), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n315), .B1(G238), .B2(new_n321), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n357), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n366), .B1(new_n361), .B2(new_n359), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n369), .B(new_n356), .C1(new_n372), .C2(new_n300), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G200), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n211), .A2(G33), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n376), .A2(new_n231), .B1(new_n211), .B2(G68), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(G50), .B2(new_n280), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT68), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n257), .B(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n381), .A2(KEYINPUT11), .ZN(new_n382));
  INV_X1    g0182(.A(G13), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(G1), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n384), .A2(KEYINPUT70), .A3(G20), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT70), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n259), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n257), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n263), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(G68), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n381), .A2(KEYINPUT11), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n385), .A2(new_n387), .ZN(new_n392));
  OAI21_X1  g0192(.A(KEYINPUT12), .B1(new_n392), .B2(G68), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT12), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n384), .A2(new_n394), .A3(G20), .A4(new_n202), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n382), .A2(new_n390), .A3(new_n391), .A4(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n368), .A2(new_n370), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT13), .ZN(new_n400));
  OAI211_X1 g0200(.A(G190), .B(new_n373), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n375), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT14), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(new_n374), .B2(G169), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  OAI211_X1 g0206(.A(G179), .B(new_n373), .C1(new_n399), .C2(new_n400), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n374), .A2(new_n404), .A3(G169), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n403), .B1(new_n409), .B2(new_n397), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n316), .B1(new_n317), .B2(new_n365), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n288), .A2(new_n306), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n412), .A2(G223), .B1(G77), .B2(new_n288), .ZN(new_n413));
  INV_X1    g0213(.A(G222), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n413), .B1(new_n414), .B2(new_n364), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n411), .B1(new_n415), .B2(new_n312), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n351), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n261), .A2(G50), .A3(new_n389), .ZN(new_n418));
  INV_X1    g0218(.A(new_n280), .ZN(new_n419));
  INV_X1    g0219(.A(G150), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n262), .B2(new_n376), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n258), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G50), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n260), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n418), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n417), .B(new_n427), .C1(G169), .C2(new_n416), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n316), .B1(new_n317), .B2(new_n232), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n412), .A2(G238), .B1(G107), .B2(new_n288), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n318), .B2(new_n364), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n430), .B1(new_n432), .B2(new_n312), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(G190), .ZN(new_n434));
  XNOR2_X1  g0234(.A(KEYINPUT15), .B(G87), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(new_n376), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(G20), .B2(G77), .ZN(new_n437));
  INV_X1    g0237(.A(new_n262), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n280), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n329), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n388), .A2(G77), .A3(new_n389), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n392), .A2(G77), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n434), .B(new_n443), .C1(new_n298), .C2(new_n433), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n433), .A2(new_n351), .ZN(new_n445));
  OR3_X1    g0245(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n445), .B(new_n446), .C1(G169), .C2(new_n433), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT9), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n427), .A2(new_n449), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n416), .A2(new_n298), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n416), .A2(G190), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n427), .A2(new_n449), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT10), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n453), .A2(new_n452), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT10), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n456), .A2(new_n457), .A3(new_n450), .A4(new_n451), .ZN(new_n458));
  AOI211_X1 g0258(.A(new_n429), .B(new_n448), .C1(new_n455), .C2(new_n458), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n355), .A2(new_n410), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT80), .ZN(new_n461));
  XNOR2_X1  g0261(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n461), .B1(new_n462), .B2(G41), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n312), .A2(new_n313), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT79), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(KEYINPUT5), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT5), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(KEYINPUT79), .ZN(new_n468));
  OAI211_X1 g0268(.A(KEYINPUT80), .B(new_n299), .C1(new_n466), .C2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G45), .ZN(new_n470));
  AOI211_X1 g0270(.A(G1), .B(new_n470), .C1(new_n467), .C2(G41), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n463), .A2(new_n464), .A3(new_n469), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n467), .A2(KEYINPUT79), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n465), .A2(KEYINPUT5), .ZN(new_n474));
  AOI21_X1  g0274(.A(G41), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n470), .A2(G1), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(KEYINPUT5), .B2(new_n299), .ZN(new_n477));
  OAI211_X1 g0277(.A(G257), .B(new_n300), .C1(new_n475), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n286), .A2(new_n287), .A3(G244), .A4(new_n306), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT4), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G250), .A2(G1698), .ZN(new_n483));
  NAND2_X1  g0283(.A1(KEYINPUT4), .A2(G244), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(G1698), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n269), .A2(new_n485), .B1(G33), .B2(G283), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n300), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(G200), .B1(new_n479), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT81), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n479), .A2(new_n487), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G190), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT6), .ZN(new_n494));
  INV_X1    g0294(.A(G97), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n494), .A2(new_n495), .A3(G107), .ZN(new_n496));
  XNOR2_X1  g0296(.A(G97), .B(G107), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n496), .B1(new_n497), .B2(new_n494), .ZN(new_n498));
  OAI22_X1  g0298(.A1(new_n498), .A2(new_n211), .B1(new_n231), .B2(new_n419), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n233), .B1(new_n270), .B2(new_n275), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n257), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n273), .A2(G1), .ZN(new_n502));
  XNOR2_X1  g0302(.A(new_n502), .B(KEYINPUT77), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n380), .A2(G97), .A3(new_n259), .A4(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n259), .A2(G97), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n501), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT78), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n501), .A2(KEYINPUT78), .A3(new_n504), .A4(new_n506), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n491), .A2(new_n489), .A3(G190), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n493), .A2(new_n509), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(G169), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n479), .B2(new_n487), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n482), .A2(new_n486), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n312), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n516), .A2(new_n351), .A3(new_n472), .A4(new_n478), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(KEYINPUT82), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT82), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n491), .A2(new_n519), .A3(new_n351), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n507), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n512), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT21), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n269), .A2(G257), .A3(new_n306), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT85), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n269), .A2(KEYINPUT85), .A3(G257), .A4(new_n306), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n412), .A2(G264), .B1(G303), .B2(new_n288), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n300), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(G270), .B(new_n300), .C1(new_n475), .C2(new_n477), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n472), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n388), .A2(new_n503), .A3(G116), .ZN(new_n535));
  INV_X1    g0335(.A(new_n392), .ZN(new_n536));
  INV_X1    g0336(.A(G116), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n256), .A2(new_n210), .B1(G20), .B2(new_n537), .ZN(new_n539));
  AOI21_X1  g0339(.A(G20), .B1(G33), .B2(G283), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(G33), .B2(new_n495), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT20), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n539), .A2(KEYINPUT20), .A3(new_n541), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n535), .B(new_n538), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G169), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n524), .B1(new_n534), .B2(new_n545), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n531), .A2(new_n533), .A3(new_n351), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n544), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n472), .A2(new_n532), .ZN(new_n549));
  INV_X1    g0349(.A(G303), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n358), .A2(new_n234), .B1(new_n550), .B2(new_n269), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n527), .B2(new_n528), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n549), .B1(new_n552), .B2(new_n300), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n553), .A2(KEYINPUT21), .A3(G169), .A4(new_n544), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n546), .A2(new_n548), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n534), .A2(G190), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n553), .A2(G200), .ZN(new_n557));
  INV_X1    g0357(.A(new_n544), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n476), .A2(new_n313), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n228), .B1(new_n470), .B2(G1), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n300), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n269), .A2(G244), .A3(G1698), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n269), .A2(G238), .A3(new_n306), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G33), .A2(G116), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n564), .B1(new_n568), .B2(new_n312), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n351), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT83), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n569), .A2(G169), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT83), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n569), .A2(new_n574), .A3(new_n351), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n571), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT84), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n380), .A2(new_n259), .A3(new_n503), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n577), .B1(new_n578), .B2(new_n435), .ZN(new_n579));
  INV_X1    g0379(.A(new_n435), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n261), .A2(KEYINPUT84), .A3(new_n580), .A4(new_n503), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n269), .A2(new_n211), .A3(G68), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT19), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n211), .B1(new_n363), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(G87), .B2(new_n206), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n584), .B1(new_n376), .B2(new_n495), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n583), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n257), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n536), .A2(new_n435), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n582), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n261), .A2(G87), .A3(new_n503), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n593), .A2(new_n589), .A3(new_n590), .ZN(new_n594));
  AOI211_X1 g0394(.A(new_n323), .B(new_n564), .C1(new_n568), .C2(new_n312), .ZN(new_n595));
  INV_X1    g0395(.A(new_n569), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n595), .B1(G200), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n576), .A2(new_n592), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n523), .A2(new_n560), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n260), .A2(new_n233), .ZN(new_n600));
  XNOR2_X1  g0400(.A(new_n600), .B(KEYINPUT25), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n578), .B2(new_n233), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT87), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT22), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(new_n211), .A3(G87), .ZN(new_n607));
  OAI21_X1  g0407(.A(KEYINPUT86), .B1(new_n288), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT86), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n227), .A2(KEYINPUT22), .A3(G20), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n269), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n286), .A2(new_n287), .A3(new_n211), .A4(G87), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n608), .A2(new_n611), .B1(KEYINPUT22), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n567), .A2(G20), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT23), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n211), .B2(G107), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n233), .A2(KEYINPUT23), .A3(G20), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n605), .B1(new_n613), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n612), .A2(KEYINPUT22), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n288), .A2(KEYINPUT86), .A3(new_n607), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n609), .B1(new_n269), .B2(new_n610), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(KEYINPUT87), .A3(new_n618), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n620), .A2(KEYINPUT24), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n257), .B1(new_n620), .B2(KEYINPUT24), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n604), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n228), .A2(new_n306), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(G257), .B2(new_n306), .ZN(new_n630));
  INV_X1    g0430(.A(G294), .ZN(new_n631));
  OAI22_X1  g0431(.A1(new_n630), .A2(new_n288), .B1(new_n273), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n312), .ZN(new_n633));
  OAI211_X1 g0433(.A(G264), .B(new_n300), .C1(new_n475), .C2(new_n477), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(new_n472), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n513), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(G179), .B2(new_n635), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT88), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n628), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(KEYINPUT87), .B1(new_n624), .B2(new_n618), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT24), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n329), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n620), .A2(new_n625), .A3(KEYINPUT24), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n603), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT88), .B1(new_n645), .B2(new_n637), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n635), .A2(new_n323), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n647), .B1(G200), .B2(new_n635), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n640), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n599), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n460), .A2(new_n651), .ZN(G372));
  XOR2_X1   g0452(.A(new_n353), .B(KEYINPUT18), .Z(new_n653));
  INV_X1    g0453(.A(new_n447), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n409), .A2(new_n397), .B1(new_n402), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n653), .B1(new_n655), .B2(new_n348), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n455), .A2(new_n458), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n429), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n460), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n572), .B1(new_n351), .B2(new_n569), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n661), .A2(new_n592), .B1(new_n597), .B2(new_n594), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n509), .A2(new_n510), .B1(new_n518), .B2(new_n520), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n662), .B1(new_n663), .B2(KEYINPUT89), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n509), .A2(new_n510), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n665), .A2(KEYINPUT89), .A3(new_n521), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n660), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n597), .A2(new_n594), .ZN(new_n668));
  INV_X1    g0468(.A(new_n592), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n571), .A2(new_n573), .A3(new_n575), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n671), .A2(new_n522), .A3(new_n660), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n661), .A2(new_n592), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  AND4_X1   g0476(.A1(new_n649), .A2(new_n512), .A3(new_n662), .A4(new_n522), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n645), .A2(new_n637), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n555), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n676), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n674), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n658), .B1(new_n659), .B2(new_n683), .ZN(G369));
  AND3_X1   g0484(.A1(new_n640), .A2(new_n646), .A3(new_n649), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n384), .A2(new_n211), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G213), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n628), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n678), .A2(new_n691), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n691), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n558), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n555), .A2(new_n698), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n546), .A2(new_n548), .A3(new_n554), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n699), .B1(new_n702), .B2(new_n698), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n696), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n700), .A2(new_n691), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n685), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n691), .B(KEYINPUT90), .Z(new_n709));
  NAND2_X1  g0509(.A1(new_n678), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n706), .A2(new_n711), .ZN(G399));
  INV_X1    g0512(.A(new_n219), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G41), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n205), .A2(new_n227), .A3(new_n537), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n714), .A2(new_n214), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n716), .B1(new_n209), .B2(new_n714), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT91), .ZN(new_n718));
  XOR2_X1   g0518(.A(new_n718), .B(KEYINPUT28), .Z(new_n719));
  INV_X1    g0519(.A(new_n522), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT26), .B1(new_n598), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n664), .A2(new_n666), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(KEYINPUT26), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n700), .A2(new_n640), .A3(new_n646), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n512), .A2(new_n662), .A3(new_n522), .A4(new_n649), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n675), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI211_X1 g0526(.A(KEYINPUT29), .B(new_n697), .C1(new_n723), .C2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n709), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n728), .B1(new_n674), .B2(new_n681), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n727), .B1(new_n729), .B2(KEYINPUT29), .ZN(new_n730));
  INV_X1    g0530(.A(G330), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n512), .A2(new_n522), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n702), .A2(new_n732), .A3(new_n671), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(new_n685), .A3(new_n709), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n534), .A2(G179), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n491), .A2(new_n634), .A3(new_n633), .A4(new_n569), .ZN(new_n736));
  OAI21_X1  g0536(.A(KEYINPUT30), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n633), .A2(new_n634), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n739), .A2(new_n479), .A3(new_n487), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n547), .A2(new_n738), .A3(new_n569), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n596), .A2(new_n635), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n351), .B1(new_n479), .B2(new_n487), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n534), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(KEYINPUT31), .A3(new_n728), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT31), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n745), .B1(new_n737), .B2(new_n741), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n749), .B1(new_n750), .B2(new_n697), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n731), .B1(new_n734), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n730), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n719), .B1(new_n756), .B2(G1), .ZN(G364));
  NOR2_X1   g0557(.A1(new_n383), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n214), .B1(new_n758), .B2(G45), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OR3_X1    g0560(.A1(new_n714), .A2(KEYINPUT92), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(KEYINPUT92), .B1(new_n714), .B2(new_n760), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n703), .A2(G330), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n705), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT93), .Z(new_n767));
  NAND3_X1  g0567(.A1(new_n219), .A2(G355), .A3(new_n269), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G116), .B2(new_n219), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n269), .B(new_n713), .C1(new_n470), .C2(new_n209), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n254), .A2(G45), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT94), .Z(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n210), .B1(G20), .B2(new_n513), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n764), .B1(new_n772), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n703), .A2(new_n776), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n323), .A2(G20), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n783), .A2(KEYINPUT96), .ZN(new_n784));
  AOI21_X1  g0584(.A(G179), .B1(new_n783), .B2(KEYINPUT96), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G200), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G159), .ZN(new_n789));
  OR3_X1    g0589(.A1(new_n788), .A2(KEYINPUT32), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(KEYINPUT32), .B1(new_n788), .B2(new_n789), .ZN(new_n791));
  NAND2_X1  g0591(.A1(G20), .A2(G179), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT95), .Z(new_n793));
  NOR2_X1   g0593(.A1(new_n323), .A2(G200), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G58), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n323), .A2(new_n298), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n797), .A2(G20), .A3(new_n351), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n227), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n793), .A2(new_n797), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n288), .B(new_n799), .C1(new_n800), .C2(G50), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n790), .A2(new_n791), .A3(new_n796), .A4(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n793), .A2(new_n323), .A3(G200), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n793), .A2(new_n323), .A3(new_n298), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(G68), .A2(new_n804), .B1(new_n806), .B2(G77), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n211), .B1(new_n794), .B2(new_n351), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT97), .Z(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G97), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n784), .A2(G200), .A3(new_n785), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n807), .B(new_n810), .C1(new_n233), .C2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(KEYINPUT33), .B(G317), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n804), .A2(new_n813), .B1(G329), .B2(new_n787), .ZN(new_n814));
  INV_X1    g0614(.A(G283), .ZN(new_n815));
  INV_X1    g0615(.A(G311), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n814), .B1(new_n815), .B2(new_n811), .C1(new_n816), .C2(new_n805), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n288), .B1(new_n798), .B2(new_n550), .ZN(new_n818));
  INV_X1    g0618(.A(new_n808), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n818), .B1(G294), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n795), .ZN(new_n821));
  INV_X1    g0621(.A(G322), .ZN(new_n822));
  INV_X1    g0622(.A(G326), .ZN(new_n823));
  INV_X1    g0623(.A(new_n800), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n820), .B1(new_n821), .B2(new_n822), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n802), .A2(new_n812), .B1(new_n817), .B2(new_n825), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n781), .B(new_n782), .C1(new_n778), .C2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n767), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G396));
  OAI21_X1  g0629(.A(new_n444), .B1(new_n443), .B2(new_n697), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n830), .A2(new_n447), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n654), .A2(new_n697), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n729), .B(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n764), .B1(new_n835), .B2(new_n754), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n754), .B2(new_n835), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n778), .A2(new_n773), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n763), .B1(new_n231), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n778), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n811), .A2(new_n227), .ZN(new_n841));
  INV_X1    g0641(.A(new_n798), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n269), .B1(new_n842), .B2(G107), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n810), .B(new_n843), .C1(new_n631), .C2(new_n821), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n841), .B(new_n844), .C1(G311), .C2(new_n787), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n800), .A2(G303), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n846), .B1(new_n537), .B2(new_n805), .C1(new_n815), .C2(new_n803), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT98), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G137), .A2(new_n800), .B1(new_n795), .B2(G143), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n849), .B1(new_n420), .B2(new_n803), .C1(new_n789), .C2(new_n805), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT34), .ZN(new_n851));
  OR2_X1    g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n787), .A2(G132), .ZN(new_n853));
  INV_X1    g0653(.A(new_n811), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(G68), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n819), .A2(G58), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n288), .B1(new_n842), .B2(G50), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n853), .A2(new_n855), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n850), .B2(new_n851), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n845), .A2(new_n848), .B1(new_n852), .B2(new_n859), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n839), .B1(new_n840), .B2(new_n860), .C1(new_n834), .C2(new_n774), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n837), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(G384));
  INV_X1    g0663(.A(new_n498), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n864), .A2(KEYINPUT35), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(KEYINPUT35), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n865), .A2(G116), .A3(new_n212), .A4(new_n866), .ZN(new_n867));
  XOR2_X1   g0667(.A(KEYINPUT99), .B(KEYINPUT36), .Z(new_n868));
  XNOR2_X1  g0668(.A(new_n867), .B(new_n868), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n209), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n425), .A2(G68), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n214), .B(G13), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n397), .B(new_n691), .C1(new_n409), .C2(new_n403), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n408), .A2(new_n407), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n397), .B1(new_n875), .B2(new_n405), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n397), .A2(new_n691), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n402), .A3(new_n877), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n665), .A2(new_n521), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT89), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n663), .A2(KEYINPUT89), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(new_n883), .A3(new_n662), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n672), .B1(new_n884), .B2(new_n660), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n675), .B1(new_n725), .B2(new_n679), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n709), .B(new_n834), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n879), .B1(new_n887), .B2(new_n832), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT38), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n293), .A2(new_n333), .A3(new_n258), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n265), .ZN(new_n891));
  INV_X1    g0691(.A(new_n689), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n344), .A2(new_n347), .ZN(new_n894));
  INV_X1    g0694(.A(new_n339), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n338), .B1(new_n337), .B2(KEYINPUT17), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n893), .B1(new_n897), .B2(new_n653), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n891), .B1(new_n352), .B2(new_n892), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n899), .A2(new_n337), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT37), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n297), .A2(new_n892), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n353), .A2(new_n337), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n889), .B1(new_n898), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n893), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n348), .B2(new_n354), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n905), .A2(new_n906), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n901), .B2(new_n900), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n910), .A2(KEYINPUT38), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n908), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n888), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n653), .B2(new_n892), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n409), .A2(new_n397), .A3(new_n697), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT39), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n910), .A2(KEYINPUT38), .A3(new_n912), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT100), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n901), .B1(new_n903), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n353), .A2(new_n903), .A3(new_n337), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n906), .A2(new_n922), .A3(new_n903), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n904), .B1(new_n348), .B2(new_n354), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT38), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n919), .B1(new_n920), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n908), .A2(KEYINPUT39), .A3(new_n913), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n916), .B1(new_n918), .B2(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n727), .B(new_n460), .C1(KEYINPUT29), .C2(new_n729), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n658), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n934), .B(new_n936), .Z(new_n937));
  INV_X1    g0737(.A(KEYINPUT101), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n874), .A2(new_n878), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n834), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n747), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n751), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n651), .B2(new_n709), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n938), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n903), .B1(new_n897), .B2(new_n653), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n925), .A2(new_n926), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n889), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n913), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n831), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n832), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n874), .B2(new_n878), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n734), .A2(new_n751), .A3(new_n941), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n938), .A2(KEYINPUT40), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT40), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n908), .A2(new_n957), .A3(new_n913), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n949), .A2(KEYINPUT40), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n659), .B2(new_n943), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n956), .A2(new_n958), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n957), .B1(new_n944), .B2(new_n948), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n460), .B(new_n953), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n960), .A2(new_n963), .A3(G330), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n937), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(KEYINPUT102), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n966), .B1(new_n214), .B2(new_n758), .C1(new_n937), .C2(new_n964), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n965), .A2(KEYINPUT102), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n873), .B1(new_n967), .B2(new_n968), .ZN(G367));
  NOR2_X1   g0769(.A1(new_n594), .A2(new_n697), .ZN(new_n970));
  MUX2_X1   g0770(.A(new_n662), .B(new_n676), .S(new_n970), .Z(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n728), .A2(new_n665), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n523), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n663), .A2(new_n728), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n640), .A2(new_n646), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n522), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n977), .A2(new_n685), .A3(new_n707), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n980), .A2(new_n709), .B1(KEYINPUT42), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(KEYINPUT42), .B2(new_n981), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n973), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n983), .A2(new_n973), .A3(new_n984), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n706), .A2(new_n978), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n988), .B(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n714), .B(KEYINPUT41), .Z(new_n991));
  NAND2_X1  g0791(.A1(new_n711), .A2(new_n977), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT45), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n708), .A2(new_n710), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n978), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT44), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n705), .B(new_n696), .C1(new_n993), .C2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n707), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n695), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(KEYINPUT103), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT103), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n695), .A2(new_n1001), .A3(new_n998), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(new_n708), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n705), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1000), .A2(new_n704), .A3(new_n708), .A4(new_n1002), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n996), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT45), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n992), .B(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1007), .A2(new_n1009), .A3(new_n706), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n997), .A2(new_n1006), .A3(new_n1010), .A4(new_n756), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n991), .B1(new_n1011), .B2(new_n756), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n759), .B1(new_n1012), .B2(KEYINPUT104), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT104), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1014), .B(new_n991), .C1(new_n1011), .C2(new_n756), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n990), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n779), .B1(new_n219), .B2(new_n435), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n713), .A2(new_n269), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1017), .B1(new_n245), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1019), .A2(new_n763), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n550), .A2(new_n821), .B1(new_n824), .B2(new_n816), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n288), .B1(new_n808), .B2(new_n233), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n798), .A2(new_n537), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT46), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n811), .A2(new_n495), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n804), .B2(G294), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n806), .A2(G283), .B1(G317), .B2(new_n787), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1025), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G50), .A2(new_n806), .B1(new_n804), .B2(G159), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n288), .B1(new_n854), .B2(G77), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1031), .A2(KEYINPUT105), .B1(KEYINPUT106), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(KEYINPUT106), .B2(new_n1032), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n809), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1035), .A2(new_n202), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G137), .B2(new_n787), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n795), .A2(G150), .B1(G58), .B2(new_n842), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n800), .A2(G143), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1037), .B(new_n1040), .C1(KEYINPUT105), .C2(new_n1031), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1029), .B1(new_n1034), .B2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT47), .Z(new_n1043));
  OAI221_X1 g0843(.A(new_n1020), .B1(new_n776), .B2(new_n971), .C1(new_n1043), .C2(new_n840), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1016), .A2(new_n1044), .ZN(G387));
  AOI22_X1  g0845(.A1(G317), .A2(new_n795), .B1(new_n800), .B2(G322), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n550), .B2(new_n805), .C1(new_n816), .C2(new_n803), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT48), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n819), .A2(G283), .B1(new_n842), .B2(G294), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT49), .Z(new_n1053));
  OAI221_X1 g0853(.A(new_n288), .B1(new_n537), .B2(new_n811), .C1(new_n788), .C2(new_n823), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT111), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n288), .B(new_n1026), .C1(new_n800), .C2(G159), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G68), .A2(new_n806), .B1(new_n804), .B2(new_n438), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT108), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n842), .A2(G77), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n788), .B2(new_n420), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1057), .B(new_n1058), .C1(new_n1059), .C2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n809), .A2(new_n580), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n425), .B2(new_n821), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT109), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1062), .B(new_n1065), .C1(new_n1059), .C2(new_n1061), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT110), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n778), .B1(new_n1056), .B2(new_n1067), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n242), .A2(new_n470), .A3(new_n269), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n1070));
  OR3_X1    g0870(.A1(new_n262), .A2(new_n1070), .A3(G50), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1070), .B1(new_n262), .B2(G50), .ZN(new_n1072));
  AOI21_X1  g0872(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n715), .B1(new_n1074), .B2(new_n288), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n219), .B1(new_n1069), .B2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1076), .B(new_n779), .C1(new_n233), .C2(new_n219), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1068), .A2(new_n764), .A3(new_n1077), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT112), .Z(new_n1079));
  NAND2_X1  g0879(.A1(new_n695), .A2(new_n777), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1079), .A2(new_n1080), .B1(new_n760), .B2(new_n1006), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1006), .A2(new_n756), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1006), .A2(new_n756), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n714), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1081), .B1(new_n1082), .B2(new_n1084), .ZN(G393));
  OAI21_X1  g0885(.A(new_n779), .B1(new_n495), .B2(new_n219), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n250), .B2(new_n1018), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(G311), .A2(new_n795), .B1(new_n800), .B2(G317), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT52), .Z(new_n1089));
  OAI221_X1 g0889(.A(new_n288), .B1(new_n798), .B2(new_n815), .C1(new_n537), .C2(new_n808), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G107), .B2(new_n854), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n788), .A2(new_n822), .B1(new_n631), .B2(new_n805), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G303), .B2(new_n804), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1089), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(G150), .A2(new_n800), .B1(new_n795), .B2(G159), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT51), .Z(new_n1096));
  AOI211_X1 g0896(.A(new_n288), .B(new_n841), .C1(G68), .C2(new_n842), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n787), .A2(G143), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n809), .A2(G77), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n425), .A2(new_n803), .B1(new_n805), .B2(new_n262), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT113), .Z(new_n1102));
  OAI21_X1  g0902(.A(new_n1094), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n763), .B(new_n1087), .C1(new_n1103), .C2(new_n778), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n776), .B2(new_n977), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n997), .A2(new_n1010), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1105), .B1(new_n1106), .B2(new_n759), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1011), .A2(new_n714), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1083), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(G390));
  AOI21_X1  g0911(.A(KEYINPUT38), .B1(new_n910), .B2(new_n912), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n920), .A2(new_n1112), .A3(new_n919), .ZN(new_n1113));
  AOI21_X1  g0913(.A(KEYINPUT39), .B1(new_n947), .B2(new_n913), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n1113), .A2(new_n1114), .B1(new_n918), .B2(new_n888), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n918), .B1(new_n947), .B2(new_n913), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n700), .A2(new_n640), .A3(new_n646), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n676), .B1(new_n677), .B2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n882), .A2(KEYINPUT26), .A3(new_n883), .A4(new_n662), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n660), .B1(new_n671), .B2(new_n522), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n691), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n833), .B1(new_n1122), .B2(new_n950), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1116), .B1(new_n879), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n753), .A2(new_n834), .A3(new_n939), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1115), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n460), .A2(new_n953), .A3(G330), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n935), .A2(new_n658), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n887), .A2(new_n832), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n939), .B1(new_n753), .B2(new_n834), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n599), .A2(new_n650), .A3(new_n728), .ZN(new_n1131));
  OAI21_X1  g0931(.A(G330), .B1(new_n1131), .B2(new_n942), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1132), .A2(new_n940), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1129), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n879), .B1(new_n1132), .B2(new_n951), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1135), .A2(new_n1125), .A3(new_n1123), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1128), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1129), .A2(new_n939), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n917), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n1122), .A2(new_n950), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n939), .B1(new_n1140), .B2(new_n833), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1139), .A2(new_n932), .B1(new_n1141), .B2(new_n1116), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1133), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1126), .B(new_n1137), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT114), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1143), .B1(new_n1115), .B2(new_n1124), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1148), .A2(KEYINPUT114), .A3(new_n1126), .A4(new_n1137), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1128), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1115), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1153), .B1(new_n1154), .B2(new_n1147), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1150), .A2(new_n714), .A3(new_n1155), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1126), .B(new_n760), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT115), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1148), .A2(KEYINPUT115), .A3(new_n760), .A4(new_n1126), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n932), .A2(new_n773), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n288), .B1(new_n227), .B2(new_n798), .C1(new_n821), .C2(new_n537), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G283), .B2(new_n800), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n495), .A2(new_n805), .B1(new_n803), .B2(new_n233), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G294), .B2(new_n787), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1163), .A2(new_n855), .A3(new_n1099), .A4(new_n1165), .ZN(new_n1166));
  OR3_X1    g0966(.A1(new_n798), .A2(KEYINPUT53), .A3(new_n420), .ZN(new_n1167));
  OAI21_X1  g0967(.A(KEYINPUT53), .B1(new_n798), .B2(new_n420), .ZN(new_n1168));
  INV_X1    g0968(.A(G128), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1167), .B(new_n1168), .C1(new_n824), .C2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(G132), .B2(new_n795), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n809), .A2(G159), .B1(new_n804), .B2(G137), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT54), .B(G143), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n806), .A2(new_n1174), .B1(G125), .B2(new_n787), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n269), .B1(new_n811), .B2(new_n425), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT116), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1171), .A2(new_n1172), .A3(new_n1175), .A4(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n840), .B1(new_n1166), .B2(new_n1178), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n763), .B(new_n1179), .C1(new_n262), .C2(new_n838), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT117), .Z(new_n1181));
  AOI22_X1  g0981(.A1(new_n1159), .A2(new_n1160), .B1(new_n1161), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1156), .A2(new_n1182), .ZN(G378));
  NAND2_X1  g0983(.A1(new_n657), .A2(new_n428), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n427), .A2(new_n892), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1184), .B(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1186), .B(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n773), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n838), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n764), .B1(G50), .B2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n269), .A2(G41), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n1060), .A2(new_n1193), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1194), .B1(new_n821), .B2(new_n233), .C1(new_n537), .C2(new_n824), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G283), .A2(new_n787), .B1(new_n854), .B2(G58), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n495), .B2(new_n803), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n805), .A2(new_n435), .ZN(new_n1198));
  NOR4_X1   g0998(.A1(new_n1195), .A2(new_n1197), .A3(new_n1036), .A4(new_n1198), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT118), .Z(new_n1200));
  AOI22_X1  g1000(.A1(new_n800), .A2(G125), .B1(new_n842), .B2(new_n1174), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n1169), .B2(new_n821), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n804), .A2(G132), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n1035), .B2(new_n420), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1202), .B(new_n1204), .C1(G137), .C2(new_n806), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n854), .A2(G159), .ZN(new_n1208));
  AOI211_X1 g1008(.A(G33), .B(G41), .C1(new_n787), .C2(G124), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1200), .A2(KEYINPUT58), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n425), .B1(G33), .B2(G41), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1212), .B1(KEYINPUT58), .B2(new_n1200), .C1(new_n1193), .C2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1192), .B1(new_n1214), .B2(new_n778), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1190), .A2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1189), .B1(new_n959), .B2(new_n731), .ZN(new_n1217));
  OAI211_X1 g1017(.A(G330), .B(new_n1188), .C1(new_n961), .C2(new_n962), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1217), .A2(new_n934), .A3(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n934), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1216), .B1(new_n1221), .B2(new_n759), .ZN(new_n1222));
  OAI21_X1  g1022(.A(KEYINPUT57), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1128), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n714), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT57), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1224), .B2(new_n1221), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1222), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(G375));
  NAND2_X1  g1030(.A1(new_n879), .A2(new_n773), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n764), .B1(G68), .B2(new_n1191), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n824), .A2(new_n631), .B1(new_n495), .B2(new_n798), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(G283), .B2(new_n795), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n804), .A2(G116), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n806), .A2(G107), .B1(G303), .B2(new_n787), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1234), .A2(new_n1063), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n288), .B1(new_n811), .B2(new_n231), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1238), .B(KEYINPUT119), .Z(new_n1239));
  NAND2_X1  g1039(.A1(new_n800), .A2(G132), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT120), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n269), .B1(new_n798), .B2(new_n789), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n795), .B2(G137), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1241), .B(new_n1243), .C1(new_n201), .C2(new_n811), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n806), .A2(G150), .B1(G128), .B2(new_n787), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1245), .B1(new_n803), .B2(new_n1173), .C1(new_n1035), .C2(new_n425), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n1237), .A2(new_n1239), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1232), .B1(new_n1247), .B2(new_n778), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1151), .A2(new_n760), .B1(new_n1231), .B2(new_n1248), .ZN(new_n1249));
  OR2_X1    g1049(.A1(new_n1137), .A2(new_n991), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1249), .B1(new_n1250), .B2(new_n1251), .ZN(G381));
  OR3_X1    g1052(.A1(G393), .A2(G396), .A3(G381), .ZN(new_n1253));
  NOR4_X1   g1053(.A1(G387), .A2(new_n1253), .A3(G384), .A4(G390), .ZN(new_n1254));
  XOR2_X1   g1054(.A(new_n1254), .B(KEYINPUT121), .Z(new_n1255));
  INV_X1    g1055(.A(KEYINPUT122), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1155), .A2(new_n714), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1161), .A2(new_n1181), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1256), .B1(new_n1258), .B2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1156), .A2(KEYINPUT122), .A3(new_n1182), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1255), .A2(new_n1229), .A3(new_n1265), .ZN(G407));
  NAND3_X1  g1066(.A1(new_n1265), .A2(new_n1229), .A3(new_n690), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(G407), .A2(G213), .A3(new_n1267), .ZN(G409));
  NOR3_X1   g1068(.A1(new_n1224), .A2(new_n1221), .A3(new_n991), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1262), .B(new_n1263), .C1(new_n1222), .C2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1222), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1272));
  OR2_X1    g1072(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT57), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(G378), .B(new_n1271), .C1(new_n1274), .C2(new_n1225), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1270), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n690), .A2(G213), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1153), .A2(KEYINPUT60), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n1152), .B2(new_n1151), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1251), .A2(KEYINPUT60), .A3(new_n1153), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1279), .A2(new_n714), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1249), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n862), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1281), .A2(G384), .A3(new_n1249), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1276), .A2(new_n1277), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(KEYINPUT62), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1277), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(G2897), .ZN(new_n1291));
  XOR2_X1   g1091(.A(new_n1291), .B(KEYINPUT124), .Z(new_n1292));
  NAND2_X1  g1092(.A1(new_n1285), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1292), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1283), .A2(new_n1284), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1289), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1290), .B1(new_n1270), .B2(new_n1275), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT62), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1299), .A2(new_n1300), .A3(new_n1286), .ZN(new_n1301));
  XOR2_X1   g1101(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1302));
  NAND4_X1  g1102(.A1(new_n1288), .A2(new_n1298), .A3(new_n1301), .A4(new_n1302), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(G393), .B(new_n828), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1016), .A2(new_n1044), .A3(G390), .ZN(new_n1306));
  AOI21_X1  g1106(.A(G390), .B1(new_n1016), .B2(new_n1044), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1305), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(G387), .A2(new_n1110), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1016), .A2(new_n1044), .A3(G390), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1309), .A2(new_n1304), .A3(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1308), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1303), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT125), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1289), .A2(new_n1314), .A3(new_n1297), .ZN(new_n1315));
  OAI21_X1  g1115(.A(KEYINPUT125), .B1(new_n1299), .B2(new_n1296), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT61), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1308), .A2(new_n1311), .A3(new_n1318), .ZN(new_n1319));
  AOI211_X1 g1119(.A(new_n1290), .B(new_n1285), .C1(new_n1270), .C2(new_n1275), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1319), .B1(new_n1320), .B2(KEYINPUT63), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT123), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1322), .B1(new_n1320), .B2(KEYINPUT63), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1287), .A2(KEYINPUT123), .A3(new_n1324), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1317), .A2(new_n1321), .A3(new_n1323), .A4(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1313), .A2(new_n1326), .ZN(G405));
  OAI21_X1  g1127(.A(new_n1275), .B1(new_n1229), .B2(new_n1264), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1329), .A2(KEYINPUT127), .A3(new_n1286), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1312), .ZN(new_n1331));
  OR2_X1    g1131(.A1(new_n1286), .A2(KEYINPUT127), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1286), .A2(KEYINPUT127), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1328), .A2(new_n1332), .A3(new_n1333), .ZN(new_n1334));
  AND3_X1   g1134(.A1(new_n1330), .A2(new_n1331), .A3(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1331), .B1(new_n1330), .B2(new_n1334), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1335), .A2(new_n1336), .ZN(G402));
endmodule


