//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT1), .B1(new_n187), .B2(G146), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(G146), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  OAI211_X1 g005(.A(G128), .B(new_n188), .C1(new_n189), .C2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n187), .A2(G146), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n193), .B(new_n194), .C1(KEYINPUT1), .C2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n192), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G125), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT0), .A2(G128), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n193), .A2(new_n194), .A3(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G143), .B(G146), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT0), .B(G128), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n201), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n199), .B1(new_n198), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G953), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n207), .A2(G224), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT7), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n199), .B(new_n210), .C1(new_n198), .C2(new_n205), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G119), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT69), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT69), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G119), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n218), .A3(G116), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n215), .A2(G116), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(KEYINPUT5), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT5), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n216), .A2(new_n218), .A3(new_n223), .A4(G116), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(G113), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G104), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT3), .B1(new_n226), .B2(G107), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n228));
  INV_X1    g042(.A(G107), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n229), .A3(G104), .ZN(new_n230));
  INV_X1    g044(.A(G101), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n226), .A2(G107), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n227), .A2(new_n230), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n226), .A2(G107), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n229), .A2(G104), .ZN(new_n235));
  OAI21_X1  g049(.A(G101), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT69), .B(G119), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n220), .B1(new_n238), .B2(G116), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT2), .ZN(new_n241));
  INV_X1    g055(.A(G113), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n243), .A2(new_n244), .B1(new_n241), .B2(new_n242), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n239), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n225), .A2(new_n237), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT84), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT84), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n225), .A2(new_n237), .A3(new_n249), .A4(new_n246), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n219), .A2(new_n221), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n243), .A2(new_n244), .ZN(new_n252));
  NOR2_X1   g066(.A1(KEYINPUT2), .A2(G113), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n227), .A2(new_n230), .A3(new_n232), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G101), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n254), .A2(new_n246), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT78), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n260), .B1(new_n255), .B2(G101), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n233), .A2(KEYINPUT4), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n255), .A2(new_n260), .A3(G101), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n248), .A2(new_n250), .B1(new_n259), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(G110), .B(G122), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n214), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(KEYINPUT8), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT86), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n225), .A2(new_n237), .A3(new_n271), .A4(new_n246), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n224), .A2(G113), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n273), .A2(new_n222), .B1(new_n245), .B2(new_n239), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n272), .B1(new_n237), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n271), .B1(new_n274), .B2(new_n237), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n270), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(G902), .B1(new_n269), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n259), .A2(new_n266), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n249), .B1(new_n274), .B2(new_n237), .ZN(new_n280));
  INV_X1    g094(.A(new_n250), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XOR2_X1   g096(.A(new_n268), .B(KEYINPUT85), .Z(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(KEYINPUT6), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT6), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(new_n267), .B2(new_n268), .ZN(new_n286));
  INV_X1    g100(.A(new_n283), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n267), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n284), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n206), .B(new_n208), .ZN(new_n290));
  AOI22_X1  g104(.A1(KEYINPUT87), .A2(new_n278), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT88), .ZN(new_n292));
  OAI21_X1  g106(.A(G210), .B1(G237), .B2(G902), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n279), .B(new_n268), .C1(new_n280), .C2(new_n281), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n212), .A2(new_n213), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n277), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT87), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n291), .A2(new_n292), .A3(new_n293), .A4(new_n300), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n294), .A2(KEYINPUT6), .B1(new_n282), .B2(new_n283), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n267), .A2(new_n285), .A3(new_n287), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n290), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n296), .A2(KEYINPUT87), .A3(new_n297), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n300), .A2(new_n304), .A3(new_n293), .A4(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT88), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n300), .A2(new_n304), .A3(new_n305), .ZN(new_n308));
  INV_X1    g122(.A(new_n293), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n301), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(G214), .B1(G237), .B2(G902), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT82), .ZN(new_n313));
  XOR2_X1   g127(.A(new_n313), .B(KEYINPUT83), .Z(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT9), .B(G234), .ZN(new_n315));
  OAI21_X1  g129(.A(G221), .B1(new_n315), .B2(G902), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT77), .ZN(new_n317));
  INV_X1    g131(.A(G469), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(new_n297), .ZN(new_n319));
  XNOR2_X1  g133(.A(G110), .B(G140), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n207), .A2(G227), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n320), .B(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n197), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n323), .A2(new_n237), .A3(KEYINPUT79), .A4(KEYINPUT10), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT79), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n192), .A2(new_n233), .A3(new_n236), .A4(new_n196), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT10), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n326), .A2(new_n327), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n255), .A2(new_n260), .A3(G101), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n331), .A2(new_n261), .A3(new_n263), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n204), .A2(KEYINPUT70), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n255), .A2(new_n258), .A3(G101), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT70), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n201), .B(new_n335), .C1(new_n202), .C2(new_n203), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n333), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n330), .B1(new_n332), .B2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n329), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G134), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT64), .B1(new_n340), .B2(G137), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT11), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT65), .B(G131), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT11), .ZN(new_n344));
  OAI211_X1 g158(.A(KEYINPUT64), .B(new_n344), .C1(new_n340), .C2(G137), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n340), .A2(G137), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n342), .A2(new_n343), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n342), .A2(KEYINPUT66), .A3(new_n345), .A4(new_n346), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G131), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n341), .A2(KEYINPUT11), .B1(new_n340), .B2(G137), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT66), .B1(new_n350), .B2(new_n345), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n347), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT80), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n342), .A2(new_n345), .A3(new_n346), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT66), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(G131), .A3(new_n348), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT80), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(new_n347), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n353), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n322), .B1(new_n339), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT81), .B1(new_n329), .B2(new_n338), .ZN(new_n363));
  INV_X1    g177(.A(new_n336), .ZN(new_n364));
  INV_X1    g178(.A(new_n200), .ZN(new_n365));
  OR2_X1    g179(.A1(KEYINPUT0), .A2(G128), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n365), .B(new_n366), .C1(new_n189), .C2(new_n191), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n335), .B1(new_n367), .B2(new_n201), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n266), .A2(new_n369), .A3(new_n334), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n324), .A2(new_n328), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT81), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n370), .A2(new_n371), .A3(new_n372), .A4(new_n330), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n363), .A2(new_n352), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n370), .A2(new_n371), .A3(new_n330), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n233), .A2(new_n236), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n197), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n326), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n352), .A2(KEYINPUT12), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT12), .B1(new_n352), .B2(new_n378), .ZN(new_n380));
  OAI22_X1  g194(.A1(new_n375), .A2(new_n360), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n362), .A2(new_n374), .B1(new_n381), .B2(new_n322), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n319), .B1(new_n382), .B2(G469), .ZN(new_n383));
  INV_X1    g197(.A(new_n322), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n339), .A2(new_n361), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n384), .B1(new_n374), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n375), .A2(new_n360), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n379), .A2(new_n380), .ZN(new_n388));
  NOR3_X1   g202(.A1(new_n387), .A2(new_n388), .A3(new_n322), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n318), .B(new_n297), .C1(new_n386), .C2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n317), .B1(new_n383), .B2(new_n390), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n311), .A2(new_n314), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT25), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT23), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n394), .B1(new_n238), .B2(G128), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n215), .A2(new_n195), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n396), .B1(new_n238), .B2(new_n195), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n395), .B1(new_n397), .B2(new_n394), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G110), .ZN(new_n399));
  XOR2_X1   g213(.A(KEYINPUT24), .B(G110), .Z(new_n400));
  NAND2_X1  g214(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G140), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G125), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n198), .A2(G140), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT75), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n405), .B(KEYINPUT16), .C1(KEYINPUT75), .C2(new_n403), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT16), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n190), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n190), .B1(new_n406), .B2(new_n408), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n399), .B(new_n401), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G125), .B(G140), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n413), .A2(new_n190), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  OAI22_X1  g229(.A1(new_n398), .A2(G110), .B1(new_n400), .B2(new_n397), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n207), .A2(G221), .A3(G234), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(KEYINPUT76), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT22), .B(G137), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n419), .B(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n412), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n421), .B1(new_n412), .B2(new_n417), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n393), .B(new_n297), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(G217), .A2(G902), .ZN(new_n426));
  INV_X1    g240(.A(G217), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n426), .B1(new_n427), .B2(G234), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n428), .B(KEYINPUT74), .Z(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n423), .A2(new_n424), .ZN(new_n433));
  OAI21_X1  g247(.A(KEYINPUT25), .B1(new_n433), .B2(G902), .ZN(new_n434));
  OR2_X1    g248(.A1(new_n423), .A2(new_n424), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n430), .A2(G902), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n432), .A2(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(G472), .A2(G902), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT32), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT30), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n204), .B1(new_n357), .B2(new_n347), .ZN(new_n442));
  OAI21_X1  g256(.A(KEYINPUT67), .B1(new_n340), .B2(G137), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT67), .ZN(new_n444));
  INV_X1    g258(.A(G137), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n445), .A3(G134), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n443), .A2(new_n446), .A3(new_n346), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G131), .ZN(new_n448));
  AND4_X1   g262(.A1(new_n196), .A2(new_n347), .A3(new_n192), .A4(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n441), .B1(new_n442), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n254), .A2(new_n246), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n352), .A2(new_n369), .ZN(new_n452));
  INV_X1    g266(.A(new_n449), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(KEYINPUT30), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n450), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n449), .B1(new_n352), .B2(new_n369), .ZN(new_n456));
  INV_X1    g270(.A(new_n451), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(G237), .A2(G953), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G210), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT27), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT26), .B(G101), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n455), .A2(new_n458), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT31), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT31), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n455), .A2(new_n466), .A3(new_n458), .A4(new_n463), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n449), .B1(new_n352), .B2(new_n205), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT71), .B1(new_n469), .B2(new_n457), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT71), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n471), .B(new_n451), .C1(new_n442), .C2(new_n449), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(new_n472), .A3(new_n458), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT28), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT28), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT72), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n457), .B1(new_n456), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n333), .A2(new_n336), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n478), .B1(new_n357), .B2(new_n347), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n479), .A2(KEYINPUT72), .A3(new_n449), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n475), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n474), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n463), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n440), .B1(new_n468), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G472), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT72), .B1(new_n479), .B2(new_n449), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n452), .A2(new_n476), .A3(new_n453), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n457), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n483), .B1(new_n489), .B2(new_n475), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n474), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n455), .A2(new_n458), .ZN(new_n492));
  AOI21_X1  g306(.A(KEYINPUT29), .B1(new_n492), .B2(new_n483), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT29), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n457), .B1(new_n452), .B2(new_n453), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n458), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n495), .B1(new_n498), .B2(KEYINPUT28), .ZN(new_n499));
  AOI21_X1  g313(.A(G902), .B1(new_n499), .B2(new_n490), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n486), .B1(new_n494), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n485), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n465), .A2(new_n467), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n463), .B1(new_n474), .B2(new_n481), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n439), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  XOR2_X1   g319(.A(KEYINPUT73), .B(KEYINPUT32), .Z(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n438), .B1(new_n502), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n187), .A2(G128), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n195), .A2(G143), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT91), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n512), .B1(new_n510), .B2(new_n511), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n340), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n510), .A2(new_n511), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT91), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(G134), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G122), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(G116), .ZN(new_n522));
  INV_X1    g336(.A(G116), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G122), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(new_n524), .A3(new_n229), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT14), .B1(new_n521), .B2(G116), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n521), .A2(G116), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT92), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT14), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n529), .B1(new_n523), .B2(G122), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT92), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n524), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n527), .A2(new_n529), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n528), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(G107), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n520), .A2(new_n525), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n510), .A2(KEYINPUT13), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(new_n340), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT13), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n522), .A2(new_n524), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G107), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n538), .A2(new_n539), .B1(new_n541), .B2(new_n525), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n515), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n315), .A2(new_n427), .A3(G953), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n536), .A2(KEYINPUT93), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n525), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n515), .B2(new_n519), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n547), .A2(new_n535), .B1(new_n515), .B2(new_n542), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n545), .B1(new_n548), .B2(new_n544), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT93), .B1(new_n548), .B2(new_n544), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n297), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT94), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n536), .A2(new_n543), .A3(new_n544), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT93), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n536), .A2(new_n543), .ZN(new_n557));
  INV_X1    g371(.A(new_n544), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(new_n559), .A3(new_n545), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(KEYINPUT94), .A3(new_n297), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n553), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(G478), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(KEYINPUT15), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n561), .A2(new_n564), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n207), .A2(G952), .ZN(new_n568));
  NAND2_X1  g382(.A1(G234), .A2(G237), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g384(.A(KEYINPUT21), .B(G898), .Z(new_n571));
  NAND3_X1  g385(.A1(new_n569), .A2(G902), .A3(G953), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(G475), .A2(G902), .ZN(new_n574));
  INV_X1    g388(.A(new_n343), .ZN(new_n575));
  INV_X1    g389(.A(G237), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n207), .A3(G214), .ZN(new_n577));
  OR2_X1    g391(.A1(KEYINPUT90), .A2(G143), .ZN(new_n578));
  NAND2_X1  g392(.A1(KEYINPUT90), .A2(G143), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n577), .A2(new_n579), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n575), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n578), .A2(new_n579), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n583), .A2(G214), .A3(new_n459), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n577), .A2(new_n579), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n343), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT17), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n582), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n406), .A2(new_n408), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G146), .ZN(new_n590));
  OAI211_X1 g404(.A(KEYINPUT17), .B(new_n575), .C1(new_n580), .C2(new_n581), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n588), .A2(new_n590), .A3(new_n409), .A4(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(G113), .B(G122), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(new_n226), .ZN(new_n594));
  AND4_X1   g408(.A1(KEYINPUT18), .A2(new_n584), .A3(G131), .A4(new_n585), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n584), .A2(new_n585), .B1(KEYINPUT18), .B2(G131), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n405), .B1(KEYINPUT75), .B2(new_n403), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(new_n190), .ZN(new_n598));
  OAI22_X1  g412(.A1(new_n595), .A2(new_n596), .B1(new_n414), .B2(new_n598), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n592), .A2(new_n594), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n582), .A2(new_n586), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n413), .A2(KEYINPUT19), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(new_n597), .B2(KEYINPUT19), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n590), .B(new_n601), .C1(G146), .C2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n594), .B1(new_n604), .B2(new_n599), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n574), .B1(new_n600), .B2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n601), .B1(G146), .B2(new_n603), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n599), .B1(new_n610), .B2(new_n411), .ZN(new_n611));
  INV_X1    g425(.A(new_n594), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n592), .A2(new_n594), .A3(new_n599), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT20), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n616), .A3(new_n574), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n594), .B1(new_n592), .B2(new_n599), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n297), .B1(new_n600), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n609), .A2(new_n617), .B1(G475), .B2(new_n619), .ZN(new_n620));
  AND4_X1   g434(.A1(new_n566), .A2(new_n567), .A3(new_n573), .A4(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n392), .A2(new_n509), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G101), .ZN(G3));
  AOI21_X1  g437(.A(new_n313), .B1(new_n310), .B2(new_n306), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n619), .A2(G475), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n607), .B1(new_n615), .B2(new_n574), .ZN(new_n626));
  INV_X1    g440(.A(new_n574), .ZN(new_n627));
  AOI211_X1 g441(.A(KEYINPUT20), .B(new_n627), .C1(new_n613), .C2(new_n614), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n625), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n549), .B2(new_n550), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n630), .B1(new_n557), .B2(new_n558), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n554), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n563), .A2(G902), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n631), .A2(KEYINPUT95), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n551), .A2(new_n563), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n560), .A2(new_n630), .B1(new_n554), .B2(new_n632), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT95), .B1(new_n638), .B2(new_n634), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n629), .B(KEYINPUT96), .C1(new_n637), .C2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n631), .A2(new_n633), .A3(new_n634), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT95), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(new_n636), .A3(new_n635), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT96), .B1(new_n645), .B2(new_n629), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n624), .B(new_n573), .C1(new_n641), .C2(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n297), .B1(new_n503), .B2(new_n504), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(G472), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n649), .A2(new_n391), .A3(new_n505), .A4(new_n437), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT34), .B(G104), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  NAND4_X1  g467(.A1(new_n615), .A2(KEYINPUT97), .A3(new_n607), .A4(new_n574), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n615), .A2(new_n607), .A3(new_n574), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT97), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n609), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n564), .B1(new_n553), .B2(new_n561), .ZN(new_n658));
  INV_X1    g472(.A(new_n567), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n654), .B(new_n657), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n573), .B(KEYINPUT98), .Z(new_n661));
  NAND2_X1  g475(.A1(new_n625), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n624), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n650), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(new_n229), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT99), .B(KEYINPUT35), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  NAND2_X1  g482(.A1(new_n432), .A2(new_n434), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n412), .A2(new_n417), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n421), .A2(KEYINPUT36), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n436), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  AND4_X1   g488(.A1(new_n621), .A2(new_n649), .A3(new_n505), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n392), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT37), .B(G110), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G12));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n570), .B(KEYINPUT100), .Z(new_n680));
  OAI21_X1  g494(.A(new_n680), .B1(G900), .B2(new_n572), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n625), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n679), .B1(new_n660), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n566), .A2(new_n567), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n657), .A2(new_n654), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n685), .A2(new_n686), .A3(KEYINPUT101), .A4(new_n682), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n674), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n502), .B2(new_n508), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n624), .A2(new_n391), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n688), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G128), .ZN(G30));
  XNOR2_X1  g507(.A(new_n681), .B(KEYINPUT39), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n391), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(KEYINPUT40), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n696), .A2(new_n313), .A3(new_n674), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n311), .B(KEYINPUT38), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n685), .A2(new_n629), .ZN(new_n699));
  INV_X1    g513(.A(new_n498), .ZN(new_n700));
  AOI21_X1  g514(.A(G902), .B1(new_n700), .B2(new_n483), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n492), .A2(new_n463), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n486), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n484), .A2(new_n465), .A3(new_n467), .ZN(new_n704));
  INV_X1    g518(.A(new_n440), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n699), .B1(new_n706), .B2(new_n508), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n695), .A2(KEYINPUT40), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n697), .A2(new_n698), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G143), .ZN(G45));
  NAND3_X1  g524(.A1(new_n645), .A2(new_n629), .A3(new_n681), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n690), .A2(new_n691), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G146), .ZN(G48));
  OAI21_X1  g528(.A(new_n297), .B1(new_n386), .B2(new_n389), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(G469), .ZN(new_n716));
  INV_X1    g530(.A(new_n317), .ZN(new_n717));
  AND3_X1   g531(.A1(new_n716), .A2(new_n717), .A3(new_n390), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n705), .B1(new_n503), .B2(new_n504), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n479), .A2(new_n451), .A3(new_n449), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT28), .B1(new_n720), .B2(new_n496), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n481), .A2(new_n721), .A3(KEYINPUT29), .A4(new_n463), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n297), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(new_n491), .B2(new_n493), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n719), .B1(new_n724), .B2(new_n486), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n506), .B1(new_n704), .B2(new_n439), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n437), .B(new_n718), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n647), .ZN(new_n728));
  XOR2_X1   g542(.A(KEYINPUT41), .B(G113), .Z(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G15));
  INV_X1    g544(.A(KEYINPUT102), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n731), .B1(new_n727), .B2(new_n664), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n663), .A2(new_n624), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n509), .A2(new_n733), .A3(KEYINPUT102), .A4(new_n718), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT103), .B(G116), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G18));
  NAND2_X1  g551(.A1(new_n494), .A2(new_n500), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(G472), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n508), .A2(new_n739), .A3(new_n719), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n674), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n718), .A2(new_n621), .A3(new_n624), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(new_n215), .ZN(G21));
  OAI211_X1 g558(.A(new_n629), .B(new_n661), .C1(new_n658), .C2(new_n659), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n718), .A2(new_n624), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n463), .B1(new_n481), .B2(new_n721), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n439), .B1(new_n503), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n649), .A2(new_n437), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n521), .ZN(G24));
  AND3_X1   g566(.A1(new_n649), .A2(new_n674), .A3(new_n749), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n753), .A2(new_n624), .A3(new_n712), .A4(new_n718), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G125), .ZN(G27));
  INV_X1    g569(.A(KEYINPUT32), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n505), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n438), .B1(new_n502), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n313), .B1(new_n308), .B2(new_n309), .ZN(new_n759));
  AND4_X1   g573(.A1(new_n307), .A2(new_n391), .A3(new_n301), .A4(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n758), .A2(KEYINPUT42), .A3(new_n760), .A4(new_n712), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n760), .A2(new_n740), .A3(new_n437), .A4(new_n712), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT104), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT42), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n763), .B1(new_n762), .B2(new_n764), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n761), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G131), .ZN(G33));
  NAND3_X1  g582(.A1(new_n688), .A2(new_n509), .A3(new_n760), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  INV_X1    g584(.A(new_n390), .ZN(new_n771));
  OAI21_X1  g585(.A(G469), .B1(new_n382), .B2(KEYINPUT45), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n772), .B1(KEYINPUT45), .B2(new_n382), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n773), .A2(new_n319), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT46), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n771), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n776), .B1(new_n775), .B2(new_n774), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n717), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n694), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT105), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n645), .A2(new_n620), .ZN(new_n782));
  XOR2_X1   g596(.A(new_n782), .B(KEYINPUT43), .Z(new_n783));
  AOI21_X1  g597(.A(new_n689), .B1(new_n505), .B2(new_n649), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XOR2_X1   g601(.A(new_n787), .B(KEYINPUT106), .Z(new_n788));
  INV_X1    g602(.A(KEYINPUT105), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n779), .A2(new_n789), .A3(new_n694), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n301), .A2(new_n307), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n759), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n792), .B1(new_n785), .B2(new_n786), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n781), .A2(new_n788), .A3(new_n790), .A4(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G137), .ZN(G39));
  NOR4_X1   g609(.A1(new_n792), .A2(new_n740), .A3(new_n437), .A4(new_n711), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n779), .A2(KEYINPUT47), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n777), .A2(KEYINPUT47), .A3(new_n717), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  INV_X1    g614(.A(new_n698), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n716), .A2(new_n390), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n802), .A2(KEYINPUT49), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(KEYINPUT49), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n437), .A2(new_n314), .A3(new_n717), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n803), .A2(new_n804), .A3(new_n782), .A4(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n801), .A2(new_n806), .A3(new_n508), .A4(new_n706), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n802), .A2(new_n717), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n797), .A2(new_n798), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n680), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n783), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n750), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OR3_X1    g627(.A1(new_n809), .A2(new_n792), .A3(new_n813), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n792), .A2(new_n317), .A3(new_n802), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT114), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n817), .A2(new_n753), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n801), .A2(new_n313), .A3(new_n718), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT113), .B1(new_n813), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n706), .A2(new_n508), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n823), .A2(new_n570), .A3(new_n438), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n815), .A2(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n825), .A2(new_n629), .A3(new_n645), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n818), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n814), .B(new_n827), .C1(new_n821), .C2(new_n820), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n817), .A2(new_n758), .ZN(new_n832));
  XOR2_X1   g646(.A(new_n832), .B(KEYINPUT48), .Z(new_n833));
  NOR2_X1   g647(.A1(new_n641), .A2(new_n646), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n718), .A2(new_n624), .ZN(new_n835));
  OAI221_X1 g649(.A(new_n568), .B1(new_n825), .B2(new_n834), .C1(new_n813), .C2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n831), .A2(new_n837), .ZN(new_n838));
  OAI22_X1  g652(.A1(new_n741), .A2(new_n742), .B1(new_n747), .B2(new_n750), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n728), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n840), .A2(new_n735), .ZN(new_n841));
  INV_X1    g655(.A(new_n661), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n629), .B1(new_n637), .B2(new_n639), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n620), .B1(new_n658), .B2(new_n659), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n845), .A2(new_n311), .A3(new_n314), .ZN(new_n846));
  INV_X1    g660(.A(new_n650), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n622), .A2(new_n848), .A3(new_n676), .ZN(new_n849));
  INV_X1    g663(.A(new_n769), .ZN(new_n850));
  INV_X1    g664(.A(new_n760), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT107), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n682), .A2(new_n657), .A3(new_n654), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n852), .B1(new_n685), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n658), .A2(new_n659), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n686), .A2(new_n855), .A3(KEYINPUT107), .A4(new_n682), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n740), .A2(new_n674), .A3(new_n854), .A4(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n712), .A2(new_n649), .A3(new_n674), .A4(new_n749), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n851), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n849), .A2(new_n850), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n767), .A2(new_n841), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT108), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n690), .B(new_n691), .C1(new_n688), .C2(new_n712), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n393), .B1(new_n435), .B2(new_n297), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n673), .B(new_n681), .C1(new_n864), .C2(new_n431), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n391), .A2(new_n866), .A3(KEYINPUT109), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT109), .B1(new_n391), .B2(new_n866), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n707), .B(new_n624), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n863), .A2(new_n754), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT52), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n863), .A2(KEYINPUT52), .A3(new_n754), .A4(new_n869), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT108), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n767), .A2(new_n841), .A3(new_n860), .A4(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n862), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n854), .A2(new_n856), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n690), .A2(new_n881), .B1(new_n753), .B2(new_n712), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n769), .B1(new_n882), .B2(new_n851), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT110), .B1(new_n883), .B2(new_n849), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n311), .A2(new_n314), .A3(new_n391), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n740), .A2(new_n621), .A3(new_n437), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n621), .A2(new_n649), .A3(new_n505), .A4(new_n674), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n845), .A2(new_n311), .A3(new_n314), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n650), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT110), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n857), .A2(new_n858), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n760), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n891), .A2(new_n892), .A3(new_n769), .A4(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n884), .A2(new_n767), .A3(new_n895), .A4(new_n841), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n874), .A2(KEYINPUT53), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT111), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n884), .A2(new_n895), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n767), .A2(new_n841), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT111), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n878), .B1(new_n872), .B2(new_n873), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n899), .A2(new_n900), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n879), .A2(new_n880), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n862), .A2(new_n876), .A3(new_n902), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n880), .B1(new_n879), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT112), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n879), .A2(new_n904), .A3(new_n880), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT112), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n862), .A2(new_n876), .ZN(new_n911));
  AOI22_X1  g725(.A1(new_n911), .A2(new_n902), .B1(new_n877), .B2(new_n878), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n909), .B(new_n910), .C1(new_n912), .C2(new_n880), .ZN(new_n913));
  AOI211_X1 g727(.A(new_n830), .B(new_n838), .C1(new_n908), .C2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(G952), .A2(G953), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n807), .B1(new_n914), .B2(new_n915), .ZN(G75));
  NOR2_X1   g730(.A1(new_n207), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n297), .B1(new_n879), .B2(new_n904), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT56), .B1(new_n919), .B2(G210), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n289), .B(new_n290), .Z(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT55), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n918), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n923), .B1(new_n920), .B2(new_n922), .ZN(G51));
  NAND2_X1  g738(.A1(new_n879), .A2(new_n904), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(KEYINPUT54), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n909), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n319), .B(KEYINPUT57), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(new_n386), .B2(new_n389), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n919), .A2(new_n773), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n917), .B1(new_n930), .B2(new_n931), .ZN(G54));
  AND3_X1   g746(.A1(new_n919), .A2(KEYINPUT58), .A3(G475), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n918), .B1(new_n933), .B2(new_n615), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n615), .B2(new_n933), .ZN(G60));
  NAND2_X1  g749(.A1(G478), .A2(G902), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT59), .Z(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n908), .A2(new_n913), .A3(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT115), .ZN(new_n940));
  INV_X1    g754(.A(new_n638), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n940), .B1(new_n939), .B2(new_n941), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n927), .A2(new_n638), .A3(new_n938), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n918), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n942), .A2(new_n943), .A3(new_n945), .ZN(G63));
  XOR2_X1   g760(.A(new_n426), .B(KEYINPUT60), .Z(new_n947));
  NAND2_X1  g761(.A1(new_n925), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n435), .B(KEYINPUT118), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n917), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n672), .B(KEYINPUT117), .Z(new_n951));
  OAI21_X1  g765(.A(new_n950), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT116), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n952), .A2(new_n953), .A3(KEYINPUT61), .ZN(new_n954));
  AOI21_X1  g768(.A(KEYINPUT61), .B1(new_n952), .B2(new_n953), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n954), .A2(new_n955), .ZN(G66));
  AOI21_X1  g770(.A(new_n207), .B1(new_n571), .B2(G224), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n841), .A2(new_n891), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n957), .B1(new_n958), .B2(new_n207), .ZN(new_n959));
  INV_X1    g773(.A(new_n289), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(G898), .B2(new_n207), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT119), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n959), .B(new_n962), .ZN(G69));
  NAND2_X1  g777(.A1(new_n450), .A2(new_n454), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(new_n603), .ZN(new_n965));
  NAND2_X1  g779(.A1(G900), .A2(G953), .ZN(new_n966));
  AND4_X1   g780(.A1(new_n685), .A2(new_n758), .A3(new_n629), .A4(new_n624), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n781), .A2(new_n790), .A3(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n968), .A2(new_n769), .A3(new_n799), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n863), .A2(new_n754), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT120), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n969), .A2(new_n767), .A3(new_n794), .A4(new_n971), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n965), .B(new_n966), .C1(new_n972), .C2(G953), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT122), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n207), .B1(G227), .B2(G900), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT123), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n695), .B1(new_n843), .B2(new_n844), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n979), .A2(new_n509), .A3(new_n791), .A4(new_n759), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT121), .Z(new_n981));
  AND2_X1   g795(.A1(new_n799), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n971), .A2(new_n709), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n983), .A2(KEYINPUT62), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(KEYINPUT62), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n982), .A2(new_n984), .A3(new_n794), .A4(new_n985), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n986), .A2(new_n207), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n973), .B1(new_n987), .B2(new_n965), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n978), .B(new_n988), .ZN(G72));
  XNOR2_X1  g803(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n486), .A2(new_n297), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n972), .B2(new_n958), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n455), .A2(new_n458), .A3(new_n483), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT126), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n917), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n992), .B1(new_n986), .B2(new_n958), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT125), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n463), .B(new_n492), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n997), .A2(new_n998), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n996), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n702), .A2(new_n994), .A3(new_n992), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n912), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(KEYINPUT127), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1001), .A2(new_n1004), .ZN(G57));
endmodule


