//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193, new_n1194;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT65), .B(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT66), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  XNOR2_X1  g013(.A(KEYINPUT68), .B(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  XNOR2_X1  g016(.A(KEYINPUT69), .B(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  AND2_X1   g018(.A1(G2072), .A2(G2078), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g027(.A1(G218), .A2(G220), .A3(G219), .A4(G221), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(G325));
  XOR2_X1   g032(.A(new_n456), .B(KEYINPUT70), .Z(G261));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n454), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(G2106), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT71), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n469), .B1(new_n465), .B2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G137), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n466), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n468), .A2(G101), .A3(G2104), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n473), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n467), .A2(G2105), .A3(new_n470), .ZN(new_n485));
  INV_X1    g060(.A(G124), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n487), .B1(G136), .B2(new_n472), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OR2_X1    g067(.A1(new_n492), .A2(new_n476), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n470), .A2(new_n464), .A3(new_n490), .A4(new_n466), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT75), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT4), .B1(new_n494), .B2(KEYINPUT75), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT73), .ZN(new_n499));
  OAI21_X1  g074(.A(G2105), .B1(KEYINPUT72), .B2(G114), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT72), .A2(G114), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OR2_X1    g079(.A1(KEYINPUT72), .A2(G114), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT72), .A2(G114), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(G2105), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n503), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(KEYINPUT73), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n467), .A2(G126), .A3(G2105), .A4(new_n470), .ZN(new_n512));
  AND3_X1   g087(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n511), .B1(new_n510), .B2(new_n512), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n498), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT76), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n518), .B(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT77), .ZN(new_n522));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(KEYINPUT77), .A2(KEYINPUT5), .A3(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n517), .A2(KEYINPUT6), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n520), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G88), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n520), .A2(G543), .A3(new_n527), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G50), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n526), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n517), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n530), .A2(new_n533), .A3(KEYINPUT78), .A4(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT78), .ZN(new_n538));
  INV_X1    g113(.A(G50), .ZN(new_n539));
  INV_X1    g114(.A(G88), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n539), .A2(new_n531), .B1(new_n528), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n538), .B1(new_n541), .B2(new_n535), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n537), .A2(new_n542), .ZN(G166));
  NAND2_X1  g118(.A1(new_n532), .A2(G51), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n529), .A2(G89), .ZN(new_n545));
  AND2_X1   g120(.A1(G63), .A2(G651), .ZN(new_n546));
  NAND3_X1  g121(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(KEYINPUT7), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(KEYINPUT7), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n526), .A2(new_n546), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n544), .A2(new_n545), .A3(new_n550), .ZN(G286));
  INV_X1    g126(.A(G286), .ZN(G168));
  INV_X1    g127(.A(G52), .ZN(new_n553));
  INV_X1    g128(.A(G90), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n553), .A2(new_n531), .B1(new_n528), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n517), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n555), .A2(new_n557), .ZN(G171));
  XNOR2_X1  g133(.A(KEYINPUT79), .B(G43), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n532), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n529), .A2(G81), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n562));
  OR2_X1    g137(.A1(new_n562), .A2(new_n517), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(new_n566));
  XOR2_X1   g141(.A(new_n566), .B(KEYINPUT80), .Z(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(KEYINPUT81), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n520), .A2(G543), .A3(new_n527), .A4(new_n573), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT9), .ZN(new_n575));
  XOR2_X1   g150(.A(KEYINPUT82), .B(G65), .Z(new_n576));
  AOI22_X1  g151(.A1(new_n526), .A2(new_n576), .B1(G78), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(new_n517), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n529), .B2(G91), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n575), .A2(new_n579), .ZN(G299));
  INV_X1    g155(.A(G171), .ZN(G301));
  INV_X1    g156(.A(G166), .ZN(G303));
  OAI21_X1  g157(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n583));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  INV_X1    g159(.A(G49), .ZN(new_n585));
  OAI221_X1 g160(.A(new_n583), .B1(new_n528), .B2(new_n584), .C1(new_n585), .C2(new_n531), .ZN(G288));
  NAND4_X1  g161(.A1(new_n520), .A2(G86), .A3(new_n526), .A4(new_n527), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n520), .A2(G48), .A3(G543), .A4(new_n527), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n524), .B2(new_n525), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT83), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT84), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g171(.A(KEYINPUT84), .B(G651), .C1(new_n591), .C2(new_n593), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n589), .A2(new_n596), .A3(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(new_n532), .A2(G47), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n529), .A2(G85), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n599), .B(new_n600), .C1(new_n517), .C2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n529), .A2(G92), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n526), .A2(G66), .ZN(new_n607));
  INV_X1    g182(.A(G79), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n523), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n532), .A2(G54), .B1(new_n609), .B2(G651), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n603), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n603), .B1(new_n612), .B2(G868), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(G299), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G280));
  XOR2_X1   g192(.A(G280), .B(KEYINPUT85), .Z(G297));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(G148));
  OAI21_X1  g195(.A(KEYINPUT86), .B1(new_n565), .B2(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n612), .A2(new_n619), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  MUX2_X1   g198(.A(KEYINPUT86), .B(new_n621), .S(new_n623), .Z(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n472), .A2(G135), .ZN(new_n626));
  INV_X1    g201(.A(G123), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n468), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  OAI221_X1 g204(.A(new_n626), .B1(new_n627), .B2(new_n485), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT88), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT89), .B(G2096), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n468), .A2(G2104), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n476), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT87), .B(KEYINPUT12), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT13), .B(G2100), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n634), .A2(new_n640), .ZN(G156));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n644), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT91), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT90), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n647), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(G14), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n652), .A2(new_n655), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(G401));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT92), .Z(new_n662));
  NOR2_X1   g237(.A1(G2072), .A2(G2078), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n444), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n660), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(KEYINPUT17), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n665), .B1(new_n662), .B2(new_n666), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n660), .B(new_n661), .C1(new_n444), .C2(new_n663), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT18), .Z(new_n669));
  NAND3_X1  g244(.A1(new_n662), .A2(new_n666), .A3(new_n660), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2096), .B(G2100), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1956), .B(G2474), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1961), .B(G1966), .ZN(new_n678));
  OR3_X1    g253(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT93), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n677), .A2(new_n678), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n677), .A2(new_n678), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n683), .B1(new_n676), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n676), .A2(KEYINPUT94), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n680), .A2(new_n681), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n682), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1981), .B(G1986), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(G229));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G20), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT23), .Z(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G299), .B2(G16), .ZN(new_n699));
  INV_X1    g274(.A(G1956), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n696), .A2(G21), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G168), .B2(new_n696), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT105), .Z(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(G1966), .ZN(new_n706));
  INV_X1    g281(.A(G2090), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G35), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G162), .B2(new_n708), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT29), .Z(new_n711));
  AOI211_X1 g286(.A(new_n701), .B(new_n706), .C1(new_n707), .C2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n612), .A2(G16), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G4), .B2(G16), .ZN(new_n714));
  INV_X1    g289(.A(G1348), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n708), .A2(G26), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT28), .ZN(new_n719));
  INV_X1    g294(.A(G128), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n468), .A2(G116), .ZN(new_n721));
  OAI21_X1  g296(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n722));
  OAI22_X1  g297(.A1(new_n485), .A2(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G140), .B2(new_n472), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n719), .B1(new_n724), .B2(new_n708), .ZN(new_n725));
  INV_X1    g300(.A(G2067), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n716), .A2(new_n717), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n708), .A2(G33), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT25), .Z(new_n731));
  AND2_X1   g306(.A1(new_n475), .A2(new_n466), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n732), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT100), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n472), .B2(G139), .ZN(new_n735));
  INV_X1    g310(.A(G139), .ZN(new_n736));
  NOR3_X1   g311(.A1(new_n471), .A2(KEYINPUT100), .A3(new_n736), .ZN(new_n737));
  OAI221_X1 g312(.A(new_n731), .B1(new_n468), .B2(new_n733), .C1(new_n735), .C2(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT101), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n729), .B1(new_n739), .B2(new_n708), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n740), .A2(G2072), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n740), .A2(G2072), .ZN(new_n742));
  NOR3_X1   g317(.A1(new_n728), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n708), .A2(G32), .ZN(new_n744));
  NAND3_X1  g319(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT103), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT26), .Z(new_n747));
  INV_X1    g322(.A(G141), .ZN(new_n748));
  INV_X1    g323(.A(G105), .ZN(new_n749));
  OAI22_X1  g324(.A1(new_n471), .A2(new_n748), .B1(new_n749), .B2(new_n635), .ZN(new_n750));
  INV_X1    g325(.A(G129), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n485), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n747), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT104), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n744), .B1(new_n755), .B2(new_n708), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT27), .B(G1996), .Z(new_n757));
  AND2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G1966), .ZN(new_n759));
  OAI22_X1  g334(.A1(new_n704), .A2(new_n759), .B1(new_n707), .B2(new_n711), .ZN(new_n760));
  INV_X1    g335(.A(G2078), .ZN(new_n761));
  NOR2_X1   g336(.A1(G164), .A2(new_n708), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G27), .B2(new_n708), .ZN(new_n763));
  AOI211_X1 g338(.A(new_n758), .B(new_n760), .C1(new_n761), .C2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n565), .A2(new_n696), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n696), .B2(G19), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G171), .A2(new_n696), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G5), .B2(new_n696), .ZN(new_n769));
  INV_X1    g344(.A(G1961), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n767), .A2(G1341), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT31), .B(G11), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT106), .B(G28), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(KEYINPUT30), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(KEYINPUT30), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n775), .A2(new_n708), .ZN(new_n776));
  INV_X1    g351(.A(G34), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(KEYINPUT24), .ZN(new_n778));
  AOI21_X1  g353(.A(G29), .B1(new_n777), .B2(KEYINPUT24), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(KEYINPUT102), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(KEYINPUT102), .B2(new_n779), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n481), .B2(new_n708), .ZN(new_n782));
  INV_X1    g357(.A(G2084), .ZN(new_n783));
  OAI221_X1 g358(.A(new_n772), .B1(new_n774), .B2(new_n776), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n783), .B2(new_n782), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n771), .A2(new_n785), .ZN(new_n786));
  OAI22_X1  g361(.A1(new_n756), .A2(new_n757), .B1(new_n763), .B2(new_n761), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n769), .A2(new_n770), .ZN(new_n788));
  OAI22_X1  g363(.A1(new_n767), .A2(G1341), .B1(new_n632), .B2(new_n708), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n786), .A2(new_n787), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n712), .A2(new_n743), .A3(new_n764), .A4(new_n790), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n696), .A2(G23), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G288), .B2(G16), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT33), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n793), .A2(new_n794), .ZN(new_n797));
  OAI21_X1  g372(.A(G1976), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n797), .ZN(new_n799));
  INV_X1    g374(.A(G1976), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n799), .A2(new_n800), .A3(new_n795), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  MUX2_X1   g377(.A(G6), .B(G305), .S(G16), .Z(new_n803));
  XOR2_X1   g378(.A(KEYINPUT32), .B(G1981), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT97), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n696), .B1(new_n537), .B2(new_n542), .ZN(new_n809));
  NOR2_X1   g384(.A1(G16), .A2(G22), .ZN(new_n810));
  OR3_X1    g385(.A1(new_n809), .A2(G1971), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(G1971), .B1(new_n809), .B2(new_n810), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n808), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n811), .A2(new_n808), .A3(new_n812), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n806), .A2(new_n807), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n802), .A2(new_n815), .A3(new_n805), .ZN(new_n817));
  OAI21_X1  g392(.A(KEYINPUT97), .B1(new_n817), .B2(new_n813), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n816), .A2(new_n818), .A3(KEYINPUT34), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT98), .ZN(new_n820));
  AOI21_X1  g395(.A(KEYINPUT34), .B1(new_n816), .B2(new_n818), .ZN(new_n821));
  MUX2_X1   g396(.A(G24), .B(G290), .S(G16), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1986), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n708), .A2(G25), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n472), .A2(G131), .ZN(new_n825));
  INV_X1    g400(.A(G119), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n468), .A2(G107), .ZN(new_n827));
  OAI21_X1  g402(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n485), .A2(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n824), .B1(new_n830), .B2(new_n708), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT35), .B(G1991), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT95), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n831), .B(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n823), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n820), .B1(new_n821), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n821), .A2(new_n820), .A3(new_n835), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n819), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT36), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n821), .ZN(new_n844));
  INV_X1    g419(.A(new_n835), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n844), .A2(KEYINPUT98), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(new_n836), .ZN(new_n847));
  INV_X1    g422(.A(new_n842), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n847), .A2(new_n819), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n791), .B1(new_n843), .B2(new_n849), .ZN(G311));
  INV_X1    g425(.A(new_n791), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n848), .B1(new_n847), .B2(new_n819), .ZN(new_n852));
  INV_X1    g427(.A(new_n819), .ZN(new_n853));
  AOI211_X1 g428(.A(new_n853), .B(new_n842), .C1(new_n846), .C2(new_n836), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n851), .B1(new_n852), .B2(new_n854), .ZN(G150));
  NOR2_X1   g430(.A1(new_n611), .A2(new_n619), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT38), .ZN(new_n857));
  INV_X1    g432(.A(G55), .ZN(new_n858));
  INV_X1    g433(.A(G93), .ZN(new_n859));
  OAI22_X1  g434(.A1(new_n858), .A2(new_n531), .B1(new_n528), .B2(new_n859), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n861), .A2(new_n517), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n565), .B(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n857), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n866));
  AOI21_X1  g441(.A(G860), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n866), .B2(new_n865), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n863), .A2(G860), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT37), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(G145));
  XNOR2_X1  g446(.A(new_n632), .B(new_n481), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(G162), .Z(new_n873));
  INV_X1    g448(.A(new_n739), .ZN(new_n874));
  OAI21_X1  g449(.A(KEYINPUT107), .B1(new_n874), .B2(KEYINPUT104), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT107), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n739), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n753), .B(new_n724), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n502), .A2(new_n499), .A3(new_n503), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT73), .B1(new_n507), .B2(new_n508), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n512), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n497), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n495), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n882), .B1(new_n884), .B2(new_n493), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n879), .B(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n878), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(G130), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n468), .A2(G118), .ZN(new_n890));
  OAI21_X1  g465(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n891));
  OAI22_X1  g466(.A1(new_n485), .A2(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n892), .B1(G142), .B2(new_n472), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n830), .B(new_n893), .Z(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n638), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n875), .A2(new_n886), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n888), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n895), .B1(new_n888), .B2(new_n896), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n873), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(G37), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n873), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT108), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n903), .B(new_n897), .C1(new_n899), .C2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n886), .B1(new_n875), .B2(new_n877), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n906), .B1(new_n886), .B2(new_n875), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n907), .A2(KEYINPUT108), .A3(new_n895), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT109), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT108), .B1(new_n907), .B2(new_n895), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n873), .B1(new_n907), .B2(new_n895), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT109), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n899), .A2(new_n904), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n910), .A2(new_n911), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n902), .B1(new_n909), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT40), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n915), .B(new_n916), .ZN(G395));
  INV_X1    g492(.A(KEYINPUT111), .ZN(new_n918));
  INV_X1    g493(.A(new_n863), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n918), .B1(new_n919), .B2(G868), .ZN(new_n920));
  XNOR2_X1  g495(.A(G166), .B(G288), .ZN(new_n921));
  XOR2_X1   g496(.A(G290), .B(G305), .Z(new_n922));
  XNOR2_X1  g497(.A(new_n921), .B(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n923), .B(KEYINPUT110), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(new_n924), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n612), .A2(new_n616), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n611), .A2(G299), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT41), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT41), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n928), .A2(new_n932), .A3(new_n929), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n622), .B(new_n864), .ZN(new_n936));
  MUX2_X1   g511(.A(new_n930), .B(new_n935), .S(new_n936), .Z(new_n937));
  OR2_X1    g512(.A1(new_n927), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G868), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n939), .B1(new_n927), .B2(new_n937), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n920), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n938), .A2(new_n940), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n941), .B1(KEYINPUT111), .B2(new_n942), .ZN(G295));
  AOI21_X1  g518(.A(new_n941), .B1(KEYINPUT111), .B2(new_n942), .ZN(G331));
  NAND3_X1  g519(.A1(new_n930), .A2(KEYINPUT113), .A3(KEYINPUT41), .ZN(new_n945));
  XNOR2_X1  g520(.A(G286), .B(G171), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n864), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n864), .A2(KEYINPUT112), .A3(new_n946), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n864), .A2(new_n946), .ZN(new_n952));
  OAI221_X1 g527(.A(new_n945), .B1(new_n951), .B2(new_n952), .C1(new_n934), .C2(KEYINPUT113), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n930), .A2(new_n952), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n947), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n923), .B(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n864), .B(new_n946), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n934), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n954), .A2(new_n949), .A3(new_n950), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(G37), .B1(new_n964), .B2(new_n926), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n959), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n964), .A2(new_n926), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n901), .B1(new_n958), .B2(new_n963), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT43), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n967), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n926), .B1(new_n953), .B2(new_n955), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT43), .B1(new_n973), .B2(new_n969), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT114), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT114), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n976), .B(KEYINPUT43), .C1(new_n973), .C2(new_n969), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n965), .B(new_n966), .C1(new_n926), .C2(new_n964), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n972), .B1(new_n979), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g555(.A(new_n724), .B(G2067), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT116), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n753), .ZN(new_n983));
  XNOR2_X1  g558(.A(KEYINPUT115), .B(G1384), .ZN(new_n984));
  INV_X1    g559(.A(new_n882), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n984), .B1(new_n985), .B2(new_n498), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n473), .A2(G40), .A3(new_n479), .A4(new_n480), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n986), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1996), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT46), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g568(.A(new_n993), .B(KEYINPUT47), .Z(new_n994));
  INV_X1    g569(.A(new_n988), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n982), .A2(new_n990), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n983), .A2(new_n996), .A3(new_n988), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n755), .A2(new_n990), .A3(new_n988), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n830), .ZN(new_n1000));
  OR3_X1    g575(.A1(new_n999), .A2(new_n833), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n724), .A2(new_n726), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n995), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(new_n830), .B(new_n833), .Z(new_n1004));
  AOI21_X1  g579(.A(new_n999), .B1(new_n988), .B2(new_n1004), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n995), .A2(G1986), .A3(G290), .ZN(new_n1006));
  XOR2_X1   g581(.A(new_n1006), .B(KEYINPUT48), .Z(new_n1007));
  AOI211_X1 g582(.A(new_n994), .B(new_n1003), .C1(new_n1005), .C2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G8), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n885), .A2(G1384), .ZN(new_n1010));
  INV_X1    g585(.A(new_n987), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(G288), .A2(new_n800), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT52), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT52), .B1(G288), .B2(new_n800), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1012), .B(new_n1016), .C1(new_n800), .C2(G288), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1981), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n589), .A2(new_n1019), .A3(new_n596), .A4(new_n597), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n587), .A2(new_n588), .A3(new_n597), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n594), .A2(new_n595), .ZN(new_n1022));
  OAI21_X1  g597(.A(G1981), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1020), .A2(new_n1023), .A3(KEYINPUT119), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n1025));
  NAND3_X1  g600(.A1(G305), .A2(new_n1025), .A3(G1981), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT49), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1028), .B(KEYINPUT120), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1027), .A2(KEYINPUT49), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(new_n1013), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1018), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n537), .A2(new_n542), .A3(G8), .ZN(new_n1034));
  XOR2_X1   g609(.A(new_n1034), .B(KEYINPUT55), .Z(new_n1035));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n1036));
  INV_X1    g611(.A(G1384), .ZN(new_n1037));
  AOI211_X1 g612(.A(KEYINPUT118), .B(new_n1036), .C1(new_n515), .C2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n515), .A2(new_n1037), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1039), .B1(new_n1040), .B2(KEYINPUT50), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n985), .A2(new_n498), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1042), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1038), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n1044), .A2(G2090), .A3(new_n987), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT45), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1040), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n987), .B1(new_n986), .B2(KEYINPUT45), .ZN(new_n1048));
  AOI21_X1  g623(.A(G1971), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT117), .ZN(new_n1050));
  INV_X1    g625(.A(G1971), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n986), .A2(KEYINPUT45), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n1011), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT45), .B1(new_n515), .B2(new_n1037), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1050), .A2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(G8), .B(new_n1035), .C1(new_n1045), .C2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1020), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1028), .A2(KEYINPUT120), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1028), .A2(KEYINPUT120), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1031), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(G288), .A2(G1976), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1060), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI22_X1  g640(.A1(new_n1033), .A2(new_n1059), .B1(new_n1065), .B2(new_n1013), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n515), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT50), .B1(new_n885), .B2(G1384), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(new_n707), .A4(new_n1011), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(G8), .B1(new_n1070), .B2(new_n1049), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n1034), .B(KEYINPUT55), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1009), .B1(new_n1055), .B2(new_n1069), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT121), .B1(new_n1075), .B2(new_n1035), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1011), .A2(new_n783), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n882), .A2(KEYINPUT74), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(G1384), .B1(new_n1081), .B2(new_n498), .ZN(new_n1082));
  OAI211_X1 g657(.A(KEYINPUT118), .B(new_n1043), .C1(new_n1082), .C2(new_n1036), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1040), .A2(new_n1039), .A3(KEYINPUT50), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1078), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1082), .A2(KEYINPUT45), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1042), .A2(new_n1037), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n987), .B1(new_n1087), .B2(new_n1046), .ZN(new_n1088));
  AOI21_X1  g663(.A(G1966), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g664(.A(G8), .B(G168), .C1(new_n1085), .C2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1077), .A2(new_n1059), .A3(new_n1032), .A4(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT63), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(G8), .B1(new_n1045), .B2(new_n1058), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1073), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1096), .A2(new_n1059), .A3(new_n1032), .A4(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1066), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1067), .A2(new_n1068), .A3(new_n1011), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n700), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n1102));
  XNOR2_X1  g677(.A(G299), .B(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT56), .B(G2072), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1047), .A2(new_n1048), .A3(new_n1104), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1101), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n715), .B1(new_n1044), .B2(new_n987), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1010), .A2(new_n726), .A3(new_n1011), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n612), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1103), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1106), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1107), .A2(KEYINPUT60), .A3(new_n611), .A4(new_n1108), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1048), .B(new_n990), .C1(new_n1082), .C2(KEYINPUT45), .ZN(new_n1116));
  XOR2_X1   g691(.A(KEYINPUT58), .B(G1341), .Z(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n1087), .B2(new_n987), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n564), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1119), .B(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1101), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1113), .A2(KEYINPUT61), .A3(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1115), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1113), .A2(new_n1122), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT123), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1103), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1128));
  OAI211_X1 g703(.A(KEYINPUT123), .B(new_n1126), .C1(new_n1106), .C2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1124), .A2(new_n1127), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT60), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1109), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1107), .A2(KEYINPUT60), .A3(new_n1108), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1133), .A2(new_n612), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1114), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1047), .A2(new_n761), .A3(new_n1048), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT53), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(G2078), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1048), .B(new_n1140), .C1(KEYINPUT45), .C2(new_n986), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n987), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1139), .B(new_n1141), .C1(new_n1142), .C2(G1961), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT126), .B1(new_n1144), .B2(G301), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1086), .A2(new_n1088), .A3(new_n1140), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1139), .B(new_n1147), .C1(new_n1142), .C2(G1961), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1146), .B1(new_n1149), .B2(G301), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1143), .A2(new_n1151), .A3(G171), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1145), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(G8), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT51), .ZN(new_n1155));
  NAND2_X1  g730(.A1(G286), .A2(G8), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1154), .A2(KEYINPUT125), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1160), .B(G8), .C1(new_n1085), .C2(new_n1089), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1159), .A2(new_n1156), .A3(new_n1161), .ZN(new_n1162));
  OAI211_X1 g737(.A(G8), .B(G286), .C1(new_n1085), .C2(new_n1089), .ZN(new_n1163));
  XNOR2_X1  g738(.A(KEYINPUT124), .B(KEYINPUT51), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1158), .B1(new_n1162), .B2(new_n1166), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1077), .A2(new_n1059), .A3(new_n1032), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1148), .A2(G171), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1143), .A2(G171), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1146), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1153), .A2(new_n1167), .A3(new_n1168), .A4(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1099), .B1(new_n1136), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT127), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n1175));
  AND2_X1   g750(.A1(new_n1161), .A2(new_n1156), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1165), .B1(new_n1176), .B2(new_n1159), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1175), .B1(new_n1177), .B2(new_n1158), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1162), .A2(new_n1166), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1179), .A2(KEYINPUT62), .A3(new_n1157), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1077), .A2(new_n1169), .A3(new_n1059), .A4(new_n1032), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1181), .ZN(new_n1182));
  AND4_X1   g757(.A1(new_n1174), .A2(new_n1178), .A3(new_n1180), .A4(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1181), .B1(new_n1167), .B2(KEYINPUT62), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1174), .B1(new_n1184), .B2(new_n1178), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1173), .A2(new_n1183), .A3(new_n1185), .ZN(new_n1186));
  XOR2_X1   g761(.A(G290), .B(G1986), .Z(new_n1187));
  OAI21_X1  g762(.A(new_n1005), .B1(new_n995), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1008), .B1(new_n1186), .B2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g764(.A1(new_n967), .A2(new_n970), .ZN(new_n1191));
  OAI211_X1 g765(.A(G319), .B(new_n673), .C1(new_n657), .C2(new_n658), .ZN(new_n1192));
  NOR2_X1   g766(.A1(G229), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g768(.A1(new_n1194), .A2(new_n915), .ZN(G308));
  OR2_X1    g769(.A1(new_n1194), .A2(new_n915), .ZN(G225));
endmodule


