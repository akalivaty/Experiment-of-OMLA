//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n568, new_n570, new_n571, new_n572, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n632, new_n633, new_n636, new_n638, new_n639, new_n640,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT67), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT69), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n463));
  AND3_X1   g038(.A1(new_n462), .A2(G137), .A3(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n465), .B1(new_n466), .B2(KEYINPUT70), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT70), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n466), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G125), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n474), .A2(new_n481), .ZN(G160));
  INV_X1    g057(.A(new_n470), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n483), .A2(new_n477), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  OAI221_X1 g062(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n477), .C2(G112), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(new_n467), .B2(new_n469), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n475), .A2(new_n476), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n462), .A2(G138), .A3(new_n463), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n465), .A2(G2104), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n491), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n461), .A2(G114), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT71), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OR2_X1    g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(G114), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n504), .A2(new_n506), .A3(new_n507), .A4(G2104), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(G126), .A2(G2105), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n470), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n495), .A2(new_n500), .A3(new_n509), .A4(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  AND2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n520), .A2(new_n521), .B1(new_n514), .B2(new_n515), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  OR2_X1    g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n526), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n523), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(G51), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n517), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n521), .A2(new_n520), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n516), .A2(G89), .ZN(new_n537));
  NAND2_X1  g112(.A1(G63), .A2(G651), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n535), .A2(new_n539), .ZN(G168));
  AOI22_X1  g115(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(new_n528), .ZN(new_n542));
  INV_X1    g117(.A(new_n522), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n514), .A2(new_n515), .ZN(new_n544));
  INV_X1    g119(.A(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(G90), .A2(new_n543), .B1(new_n546), .B2(G52), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G52), .ZN(new_n550));
  INV_X1    g125(.A(G90), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n517), .A2(new_n550), .B1(new_n551), .B2(new_n522), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(KEYINPUT72), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n542), .B1(new_n549), .B2(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  AOI22_X1  g130(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n528), .ZN(new_n557));
  XNOR2_X1  g132(.A(KEYINPUT73), .B(G81), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n543), .A2(new_n558), .B1(new_n546), .B2(G43), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n557), .A2(new_n559), .A3(KEYINPUT74), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(G860), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT75), .ZN(G153));
  AND3_X1   g142(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G36), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT76), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G188));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  INV_X1    g149(.A(G78), .ZN(new_n575));
  OAI22_X1  g150(.A1(new_n536), .A2(new_n574), .B1(new_n575), .B2(new_n545), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT78), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n578));
  OAI221_X1 g153(.A(new_n578), .B1(new_n575), .B2(new_n545), .C1(new_n536), .C2(new_n574), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(G651), .A3(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(G53), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n581), .B1(new_n582), .B2(KEYINPUT9), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n546), .B(new_n583), .C1(new_n582), .C2(KEYINPUT9), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n582), .A2(KEYINPUT9), .ZN(new_n585));
  INV_X1    g160(.A(new_n583), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n517), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n543), .A2(G91), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n580), .A2(new_n584), .A3(new_n587), .A4(new_n588), .ZN(G299));
  OR2_X1    g164(.A1(new_n535), .A2(new_n539), .ZN(G286));
  NAND2_X1  g165(.A1(new_n543), .A2(G87), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n546), .A2(G49), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(G288));
  OAI211_X1 g169(.A(G48), .B(G543), .C1(new_n514), .C2(new_n515), .ZN(new_n595));
  INV_X1    g170(.A(G86), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n522), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(KEYINPUT79), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n601), .A2(G73), .A3(G543), .ZN(new_n602));
  INV_X1    g177(.A(G61), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n600), .B(new_n602), .C1(new_n536), .C2(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(KEYINPUT80), .B1(new_n604), .B2(G651), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n603), .B1(new_n524), .B2(new_n525), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n600), .A2(new_n602), .ZN(new_n607));
  OAI211_X1 g182(.A(KEYINPUT80), .B(G651), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n598), .B1(new_n605), .B2(new_n609), .ZN(G305));
  NAND2_X1  g185(.A1(new_n543), .A2(G85), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n546), .A2(G47), .ZN(new_n613));
  AND3_X1   g188(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n612), .B1(new_n611), .B2(new_n613), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n616));
  OAI22_X1  g191(.A1(new_n614), .A2(new_n615), .B1(new_n528), .B2(new_n616), .ZN(G290));
  NAND2_X1  g192(.A1(G301), .A2(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n543), .A2(G92), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT10), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n526), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n622));
  INV_X1    g197(.A(G54), .ZN(new_n623));
  OAI22_X1  g198(.A1(new_n622), .A2(new_n528), .B1(new_n517), .B2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT82), .ZN(new_n625));
  AND2_X1   g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n621), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n618), .B1(new_n629), .B2(G868), .ZN(G284));
  OAI21_X1  g205(.A(new_n618), .B1(new_n629), .B2(G868), .ZN(G321));
  NAND2_X1  g206(.A1(G286), .A2(G868), .ZN(new_n632));
  AND4_X1   g207(.A1(new_n580), .A2(new_n584), .A3(new_n587), .A4(new_n588), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(G868), .ZN(G297));
  OAI21_X1  g209(.A(new_n632), .B1(new_n633), .B2(G868), .ZN(G280));
  AOI21_X1  g210(.A(new_n628), .B1(G559), .B2(new_n565), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT83), .Z(G148));
  INV_X1    g212(.A(G868), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n564), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n628), .A2(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(new_n638), .ZN(G323));
  XNOR2_X1  g216(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g217(.A1(new_n478), .A2(new_n472), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT12), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT13), .ZN(new_n646));
  AOI22_X1  g221(.A1(new_n645), .A2(new_n646), .B1(KEYINPUT84), .B2(G2100), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n646), .B2(new_n645), .ZN(new_n648));
  OR3_X1    g223(.A1(new_n648), .A2(KEYINPUT84), .A3(G2100), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n648), .B1(KEYINPUT84), .B2(G2100), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n484), .A2(G135), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n486), .A2(G123), .ZN(new_n652));
  OAI221_X1 g227(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n477), .C2(G111), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(G2096), .Z(new_n655));
  NAND3_X1  g230(.A1(new_n649), .A2(new_n650), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT85), .Z(G156));
  INV_X1    g232(.A(KEYINPUT14), .ZN(new_n658));
  XOR2_X1   g233(.A(KEYINPUT15), .B(G2435), .Z(new_n659));
  XOR2_X1   g234(.A(KEYINPUT86), .B(G2438), .Z(new_n660));
  XOR2_X1   g235(.A(new_n659), .B(new_n660), .Z(new_n661));
  XNOR2_X1  g236(.A(G2427), .B(G2430), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n658), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT87), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n662), .B2(new_n661), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1341), .B(G1348), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2451), .B(G2454), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT16), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(new_n669), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(G14), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n672), .B1(new_n670), .B2(new_n673), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(G401));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  XNOR2_X1  g253(.A(G2067), .B(G2678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n680), .A2(KEYINPUT17), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n678), .A2(new_n679), .ZN(new_n682));
  AOI21_X1  g257(.A(KEYINPUT18), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2072), .B(G2078), .Z(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n680), .B2(KEYINPUT18), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G2096), .B(G2100), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G227));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT89), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1956), .B(G2474), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1971), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT20), .Z(new_n698));
  OR2_X1    g273(.A1(new_n690), .A2(new_n692), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n699), .A2(new_n693), .A3(new_n696), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n698), .B(new_n700), .C1(new_n696), .C2(new_n699), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1991), .B(G1996), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1981), .B(G1986), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n705), .B(new_n706), .Z(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(G229));
  XNOR2_X1  g283(.A(KEYINPUT98), .B(KEYINPUT23), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G20), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n709), .B(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G299), .B2(G16), .ZN(new_n713));
  INV_X1    g288(.A(G1956), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT24), .B(G34), .ZN(new_n716));
  MUX2_X1   g291(.A(new_n716), .B(G160), .S(G29), .Z(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(G2084), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(G2084), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n720), .A2(G32), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n484), .A2(G141), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n486), .A2(G129), .ZN(new_n723));
  NAND3_X1  g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT26), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n726), .A2(new_n727), .B1(G105), .B2(new_n472), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n722), .A2(new_n723), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n721), .B1(new_n729), .B2(G29), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT27), .B(G1996), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n718), .A2(new_n719), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G2078), .ZN(new_n733));
  NAND2_X1  g308(.A1(G164), .A2(G29), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G27), .B2(G29), .ZN(new_n735));
  INV_X1    g310(.A(G2090), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n720), .A2(G35), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT97), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n489), .B2(G29), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT29), .ZN(new_n740));
  OAI221_X1 g315(.A(new_n732), .B1(new_n733), .B2(new_n735), .C1(new_n736), .C2(new_n740), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n715), .B(new_n741), .C1(new_n736), .C2(new_n740), .ZN(new_n742));
  INV_X1    g317(.A(new_n564), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(new_n710), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n710), .B2(G19), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT93), .B(G1341), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n710), .A2(G5), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G171), .B2(new_n710), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n745), .A2(new_n746), .B1(G1961), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT30), .B(G28), .ZN(new_n750));
  OR2_X1    g325(.A1(KEYINPUT31), .A2(G11), .ZN(new_n751));
  NAND2_X1  g326(.A1(KEYINPUT31), .A2(G11), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n750), .A2(new_n720), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n710), .A2(G21), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G168), .B2(new_n710), .ZN(new_n755));
  OAI221_X1 g330(.A(new_n753), .B1(new_n720), .B2(new_n654), .C1(new_n755), .C2(G1966), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G1966), .B2(new_n755), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n730), .A2(new_n731), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n733), .B2(new_n735), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n749), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n720), .A2(G26), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT28), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n484), .A2(G140), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n486), .A2(G128), .ZN(new_n764));
  OAI221_X1 g339(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n477), .C2(G116), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n762), .B1(new_n766), .B2(G29), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G2067), .ZN(new_n768));
  OAI221_X1 g343(.A(new_n768), .B1(G1961), .B2(new_n748), .C1(new_n745), .C2(new_n746), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n760), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n710), .A2(G4), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n629), .B2(new_n710), .ZN(new_n772));
  INV_X1    g347(.A(G1348), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G29), .A2(G33), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT94), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n484), .A2(G139), .ZN(new_n777));
  AND2_X1   g352(.A1(G103), .A2(G2104), .ZN(new_n778));
  AOI21_X1  g353(.A(KEYINPUT25), .B1(new_n477), .B2(new_n778), .ZN(new_n779));
  AND3_X1   g354(.A1(new_n477), .A2(KEYINPUT25), .A3(new_n778), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n777), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n781), .A2(KEYINPUT95), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(KEYINPUT95), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n478), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n784), .A2(new_n477), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT96), .Z(new_n786));
  NAND3_X1  g361(.A1(new_n782), .A2(new_n783), .A3(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n776), .B1(new_n787), .B2(new_n720), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G2072), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n742), .A2(new_n770), .A3(new_n774), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n710), .A2(G6), .ZN(new_n791));
  OAI21_X1  g366(.A(G651), .B1(new_n606), .B2(new_n607), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT80), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n597), .B1(new_n794), .B2(new_n608), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n791), .B1(new_n795), .B2(new_n710), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT92), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT32), .B(G1981), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n710), .A2(G22), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G166), .B2(new_n710), .ZN(new_n802));
  INV_X1    g377(.A(G1971), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n710), .A2(G23), .ZN(new_n805));
  INV_X1    g380(.A(G288), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(new_n710), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT33), .B(G1976), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n799), .A2(new_n800), .A3(new_n804), .A4(new_n809), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n810), .A2(KEYINPUT34), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n810), .A2(KEYINPUT34), .ZN(new_n812));
  NAND2_X1  g387(.A1(G290), .A2(G16), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n710), .A2(G24), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n815), .A2(G1986), .ZN(new_n816));
  NOR2_X1   g391(.A1(G25), .A2(G29), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n477), .A2(G107), .ZN(new_n818));
  OAI21_X1  g393(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n486), .A2(G119), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n484), .A2(G131), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n822), .A2(KEYINPUT90), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n822), .A2(KEYINPUT90), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n817), .B1(new_n826), .B2(G29), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT35), .B(G1991), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT91), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n816), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n815), .A2(G1986), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n830), .B(new_n831), .C1(new_n827), .C2(new_n829), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n811), .A2(new_n812), .A3(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n790), .B1(new_n835), .B2(new_n836), .ZN(G311));
  XOR2_X1   g412(.A(G311), .B(KEYINPUT99), .Z(G150));
  INV_X1    g413(.A(G55), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT100), .B(G93), .ZN(new_n840));
  OAI22_X1  g415(.A1(new_n517), .A2(new_n839), .B1(new_n522), .B2(new_n840), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(new_n528), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n562), .B2(new_n563), .ZN(new_n845));
  INV_X1    g420(.A(new_n844), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(new_n560), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n629), .A2(G559), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n852), .A2(new_n565), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n844), .A2(new_n565), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(G145));
  XNOR2_X1  g432(.A(new_n766), .B(G164), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n729), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n787), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n825), .B(new_n645), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n486), .A2(G130), .ZN(new_n862));
  OAI221_X1 g437(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n477), .C2(G118), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(G142), .B2(new_n484), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n861), .B(new_n865), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n860), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n654), .B(G160), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(G162), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(KEYINPUT101), .B1(new_n860), .B2(new_n866), .ZN(new_n871));
  OR3_X1    g446(.A1(new_n860), .A2(KEYINPUT101), .A3(new_n866), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(G37), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n860), .A2(new_n866), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n869), .B1(new_n867), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n873), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g453(.A1(new_n846), .A2(new_n638), .ZN(new_n879));
  XNOR2_X1  g454(.A(G290), .B(new_n795), .ZN(new_n880));
  XNOR2_X1  g455(.A(G303), .B(G288), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT42), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n848), .B(new_n640), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n633), .B(new_n621), .C1(new_n627), .C2(new_n626), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n628), .A2(G299), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT102), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT102), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT41), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT41), .B1(new_n885), .B2(new_n886), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n889), .B1(new_n893), .B2(new_n884), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n883), .B(new_n894), .Z(new_n895));
  OAI21_X1  g470(.A(new_n879), .B1(new_n895), .B2(new_n638), .ZN(G295));
  OAI21_X1  g471(.A(new_n879), .B1(new_n895), .B2(new_n638), .ZN(G331));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n552), .B(KEYINPUT72), .ZN(new_n899));
  AOI21_X1  g474(.A(G168), .B1(new_n899), .B2(new_n542), .ZN(new_n900));
  OAI211_X1 g475(.A(G168), .B(new_n542), .C1(new_n549), .C2(new_n553), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OAI22_X1  g477(.A1(new_n900), .A2(new_n902), .B1(new_n845), .B2(new_n847), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n564), .A2(new_n846), .ZN(new_n904));
  INV_X1    g479(.A(new_n847), .ZN(new_n905));
  NAND2_X1  g480(.A1(G301), .A2(G286), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .A4(new_n901), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n903), .A2(new_n907), .A3(KEYINPUT103), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT103), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n848), .A2(new_n909), .A3(new_n906), .A4(new_n901), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n888), .A2(new_n887), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n903), .A2(new_n907), .ZN(new_n913));
  OAI22_X1  g488(.A1(new_n893), .A2(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n882), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n885), .A2(new_n886), .ZN(new_n916));
  AOI22_X1  g491(.A1(new_n911), .A2(new_n916), .B1(new_n892), .B2(new_n913), .ZN(new_n917));
  INV_X1    g492(.A(new_n882), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n915), .A2(new_n919), .A3(new_n874), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n920), .A2(KEYINPUT43), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n921), .B(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  OAI211_X1 g499(.A(KEYINPUT104), .B(new_n874), .C1(new_n917), .C2(new_n918), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n925), .A2(new_n919), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n874), .B1(new_n917), .B2(new_n918), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n924), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n898), .B1(new_n923), .B2(new_n930), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n929), .A2(new_n924), .A3(new_n925), .A4(new_n919), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT106), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n926), .A2(new_n934), .A3(new_n924), .A4(new_n929), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n915), .A2(new_n919), .A3(KEYINPUT107), .A4(new_n874), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n920), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n898), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n936), .A2(KEYINPUT108), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT108), .B1(new_n936), .B2(new_n941), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n931), .B1(new_n942), .B2(new_n943), .ZN(G397));
  INV_X1    g519(.A(KEYINPUT55), .ZN(new_n945));
  INV_X1    g520(.A(G8), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n945), .B1(G166), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n949), .A2(KEYINPUT111), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n951), .B1(new_n947), .B2(new_n948), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G1384), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n512), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT50), .ZN(new_n956));
  INV_X1    g531(.A(G40), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n474), .A2(new_n481), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n512), .A2(new_n959), .A3(new_n954), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n956), .A2(new_n736), .A3(new_n958), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT109), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n955), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n512), .A2(KEYINPUT45), .A3(new_n954), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n958), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n803), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n959), .B1(new_n512), .B2(new_n954), .ZN(new_n968));
  AOI22_X1  g543(.A1(new_n464), .A2(new_n470), .B1(G101), .B2(new_n472), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n479), .A2(new_n480), .ZN(new_n970));
  OAI211_X1 g545(.A(G40), .B(new_n969), .C1(new_n970), .C2(new_n477), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n972), .A2(new_n973), .A3(new_n736), .A4(new_n960), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n962), .A2(new_n967), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT110), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n962), .A2(new_n967), .A3(new_n974), .A4(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n953), .A2(new_n976), .A3(G8), .A4(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT115), .B1(new_n968), .B2(new_n971), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT115), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n477), .A2(new_n478), .A3(G138), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n982), .A2(new_n491), .B1(new_n492), .B2(new_n494), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n503), .A2(new_n508), .B1(new_n470), .B2(new_n510), .ZN(new_n984));
  AOI21_X1  g559(.A(G1384), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n958), .B(new_n981), .C1(new_n985), .C2(new_n959), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n980), .A2(new_n986), .A3(new_n736), .A4(new_n960), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n967), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n946), .B1(new_n988), .B2(KEYINPUT116), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n987), .A2(new_n990), .A3(new_n967), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n949), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n958), .B1(new_n985), .B2(KEYINPUT45), .ZN(new_n993));
  INV_X1    g568(.A(new_n965), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT117), .B1(new_n995), .B2(G1966), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n997));
  INV_X1    g572(.A(G1966), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n997), .B(new_n998), .C1(new_n993), .C2(new_n994), .ZN(new_n999));
  INV_X1    g574(.A(G2084), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n972), .A2(new_n1000), .A3(new_n960), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n996), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT63), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n1002), .A2(new_n1003), .A3(G8), .A4(G168), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n979), .B1(new_n992), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n946), .B1(new_n958), .B2(new_n985), .ZN(new_n1006));
  INV_X1    g581(.A(G1976), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1006), .B1(new_n1007), .B2(G288), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT52), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n806), .B2(G1976), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n1013));
  INV_X1    g588(.A(G1981), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n795), .A2(new_n1014), .ZN(new_n1015));
  AOI211_X1 g590(.A(G1981), .B(new_n597), .C1(new_n794), .C2(new_n608), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(G305), .A2(G1981), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n795), .A2(new_n1014), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(KEYINPUT112), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT49), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1017), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT113), .B1(new_n1023), .B2(KEYINPUT49), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1018), .A2(KEYINPUT49), .A3(new_n1019), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1022), .B(new_n1006), .C1(new_n1024), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1025), .B(new_n1026), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1031), .A2(KEYINPUT114), .A3(new_n1022), .A4(new_n1006), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1012), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1005), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n806), .A2(new_n1007), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1035), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1006), .B1(new_n1036), .B2(new_n1016), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n999), .A2(new_n1001), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n997), .B1(new_n966), .B2(new_n998), .ZN(new_n1040));
  OAI211_X1 g615(.A(G8), .B(G168), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  AOI211_X1 g616(.A(new_n1012), .B(new_n1041), .C1(new_n1030), .C2(new_n1032), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n975), .A2(KEYINPUT110), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n978), .A2(G8), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT118), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n949), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n976), .A2(new_n1047), .A3(G8), .A4(new_n978), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1003), .B1(new_n1042), .B2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1038), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(G168), .A2(new_n946), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT123), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1054), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n996), .A2(KEYINPUT123), .A3(new_n999), .A4(new_n1001), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1053), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n946), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1053), .B1(new_n1058), .B2(KEYINPUT124), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT124), .ZN(new_n1060));
  AOI211_X1 g635(.A(new_n1060), .B(new_n946), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT51), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1002), .A2(G8), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1063), .A2(KEYINPUT51), .A3(new_n1052), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1057), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1067), .A2(KEYINPUT57), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(KEYINPUT57), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n633), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(G299), .A2(new_n1067), .A3(KEYINPUT57), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n980), .A2(new_n960), .A3(new_n986), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n714), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT56), .B(G2072), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n995), .A2(new_n1075), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1072), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1072), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n958), .A2(new_n985), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(G2067), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n972), .A2(new_n960), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n1085), .B2(new_n773), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1082), .B1(new_n628), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1081), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1078), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1086), .A2(KEYINPUT60), .A3(new_n628), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n628), .B1(new_n1086), .B2(KEYINPUT60), .ZN(new_n1091));
  OAI22_X1  g666(.A1(new_n1090), .A2(new_n1091), .B1(KEYINPUT60), .B2(new_n1086), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT61), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1073), .A2(new_n714), .B1(new_n995), .B2(new_n1075), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1093), .B1(new_n1094), .B2(new_n1072), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1095), .A2(new_n1077), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1079), .A2(new_n1080), .A3(new_n1093), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1092), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT58), .B(G1341), .Z(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1101), .B1(new_n958), .B2(new_n985), .ZN(new_n1102));
  INV_X1    g677(.A(G1996), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n964), .A2(new_n1103), .A3(new_n958), .A4(new_n965), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1102), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n971), .B1(new_n955), .B2(new_n963), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1107), .A2(KEYINPUT121), .A3(new_n1103), .A4(new_n965), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n564), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1099), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1102), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(new_n1108), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n743), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT122), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(KEYINPUT122), .A3(new_n1099), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1089), .B1(new_n1098), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n992), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n966), .A2(G2078), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1122), .A2(KEYINPUT53), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1107), .A2(KEYINPUT53), .A3(new_n733), .A4(new_n965), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n956), .A2(new_n958), .A3(new_n960), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1124), .B1(new_n1125), .B2(G1961), .ZN(new_n1126));
  XNOR2_X1  g701(.A(G301), .B(KEYINPUT54), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1123), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(KEYINPUT125), .ZN(new_n1129));
  OR2_X1    g704(.A1(new_n1122), .A2(KEYINPUT53), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1124), .B(new_n1131), .C1(new_n1125), .C2(G1961), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1129), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1128), .B1(new_n1133), .B2(new_n1127), .ZN(new_n1134));
  AND4_X1   g709(.A1(new_n1121), .A2(new_n1033), .A3(new_n1134), .A4(new_n979), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1120), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1051), .B1(new_n1066), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(G8), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n1060), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1058), .A2(KEYINPUT124), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1142), .A2(new_n1143), .A3(new_n1053), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1064), .B1(new_n1144), .B2(KEYINPUT51), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT62), .B1(new_n1145), .B2(new_n1057), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1066), .A2(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1133), .A2(G171), .ZN(new_n1149));
  AND4_X1   g724(.A1(new_n1121), .A2(new_n1033), .A3(new_n1149), .A4(new_n979), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1146), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1051), .B(KEYINPUT126), .C1(new_n1066), .C2(new_n1136), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1139), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n964), .A2(new_n971), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n826), .A2(new_n828), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n766), .B(G2067), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n729), .B(G1996), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n826), .A2(new_n828), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1155), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(G290), .B(G1986), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1154), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1153), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1154), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1158), .A2(new_n826), .A3(new_n828), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n766), .A2(G2067), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT46), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1168), .B1(new_n1164), .B2(G1996), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1154), .B1(new_n1156), .B2(new_n729), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1154), .A2(KEYINPUT46), .A3(new_n1103), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  XOR2_X1   g747(.A(new_n1172), .B(KEYINPUT47), .Z(new_n1173));
  NAND2_X1  g748(.A1(new_n1160), .A2(new_n1154), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1164), .A2(G1986), .A3(G290), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n1175), .B(KEYINPUT48), .Z(new_n1176));
  AOI211_X1 g751(.A(new_n1167), .B(new_n1173), .C1(new_n1174), .C2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1163), .A2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g753(.A1(new_n923), .A2(new_n930), .ZN(new_n1180));
  INV_X1    g754(.A(G319), .ZN(new_n1181));
  NOR2_X1   g755(.A1(G227), .A2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g756(.A(new_n1182), .B1(new_n675), .B2(new_n676), .ZN(new_n1183));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n1184));
  NAND2_X1  g758(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g759(.A(KEYINPUT127), .B(new_n1182), .C1(new_n675), .C2(new_n676), .ZN(new_n1186));
  NAND4_X1  g760(.A1(new_n707), .A2(new_n1185), .A3(new_n877), .A4(new_n1186), .ZN(new_n1187));
  NOR2_X1   g761(.A1(new_n1180), .A2(new_n1187), .ZN(G308));
  OR2_X1    g762(.A1(new_n1180), .A2(new_n1187), .ZN(G225));
endmodule


