//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n547, new_n548, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1166,
    new_n1167, new_n1168;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT66), .ZN(new_n447));
  XNOR2_X1  g022(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT68), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  OR2_X1    g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(G2105), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n463), .A2(G137), .B1(G101), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n467), .B1(new_n461), .B2(new_n462), .ZN(new_n468));
  AND2_X1   g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n466), .A2(new_n470), .ZN(G160));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n472), .B1(new_n461), .B2(new_n462), .ZN(new_n473));
  MUX2_X1   g048(.A(G100), .B(G112), .S(G2105), .Z(new_n474));
  AOI22_X1  g049(.A1(G124), .A2(new_n473), .B1(new_n474), .B2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(G136), .ZN(new_n476));
  INV_X1    g051(.A(new_n463), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT69), .ZN(G162));
  AND2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  OAI211_X1 g056(.A(G138), .B(new_n472), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT4), .ZN(new_n483));
  XNOR2_X1  g058(.A(KEYINPUT3), .B(G2104), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n484), .A2(new_n485), .A3(G138), .A4(new_n472), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(G114), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G102), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n473), .A2(G126), .B1(G2104), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G164));
  INV_X1    g068(.A(G50), .ZN(new_n494));
  AND2_X1   g069(.A1(KEYINPUT6), .A2(G651), .ZN(new_n495));
  NOR2_X1   g070(.A1(KEYINPUT6), .A2(G651), .ZN(new_n496));
  OR2_X1    g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G543), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G88), .ZN(new_n505));
  OAI22_X1  g080(.A1(new_n494), .A2(new_n498), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n506), .A2(new_n509), .ZN(G166));
  NAND3_X1  g085(.A1(new_n503), .A2(G63), .A3(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n495), .A2(new_n496), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n512), .A2(new_n500), .ZN(new_n513));
  AOI22_X1  g088(.A1(KEYINPUT70), .A2(new_n511), .B1(new_n513), .B2(G51), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n511), .A2(KEYINPUT70), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n514), .A2(KEYINPUT71), .A3(new_n515), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n520), .B(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n503), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n512), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n522), .B1(G89), .B2(new_n524), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n518), .A2(new_n519), .A3(new_n525), .ZN(G168));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n527));
  INV_X1    g102(.A(G52), .ZN(new_n528));
  INV_X1    g103(.A(G90), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n528), .A2(new_n498), .B1(new_n504), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n508), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n527), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n524), .A2(G90), .B1(G52), .B2(new_n513), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n531), .A2(new_n508), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT73), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n533), .A2(new_n536), .ZN(G171));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n538), .A2(new_n498), .B1(new_n504), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n508), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  AND3_X1   g119(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G36), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n545), .A2(new_n548), .ZN(G188));
  NAND2_X1  g124(.A1(new_n513), .A2(G53), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT9), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n503), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n508), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(G91), .B2(new_n524), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n551), .A2(new_n554), .A3(KEYINPUT74), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(KEYINPUT74), .B1(new_n551), .B2(new_n554), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n556), .A2(new_n557), .ZN(G299));
  INV_X1    g133(.A(KEYINPUT75), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n559), .B1(new_n533), .B2(new_n536), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n533), .A2(new_n536), .A3(new_n559), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(G301));
  NAND3_X1  g139(.A1(new_n518), .A2(new_n519), .A3(new_n525), .ZN(G286));
  INV_X1    g140(.A(G166), .ZN(G303));
  NAND2_X1  g141(.A1(new_n524), .A2(G87), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n513), .A2(G49), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n503), .B2(G74), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(G288));
  NAND2_X1  g145(.A1(new_n513), .A2(G48), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n497), .A2(G86), .A3(new_n503), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n501), .B2(new_n502), .ZN(new_n575));
  AND2_X1   g150(.A1(G73), .A2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G305));
  NAND2_X1  g155(.A1(G72), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G60), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n523), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n508), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n585), .B1(new_n584), .B2(new_n583), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT77), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n586), .B(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n524), .A2(G85), .B1(G47), .B2(new_n513), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(new_n524), .A2(G92), .ZN(new_n591));
  XOR2_X1   g166(.A(new_n591), .B(KEYINPUT10), .Z(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n523), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(new_n513), .B2(G54), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(new_n563), .B2(new_n598), .ZN(G284));
  OAI21_X1  g175(.A(new_n599), .B1(new_n563), .B2(new_n598), .ZN(G321));
  NAND2_X1  g176(.A1(G286), .A2(G868), .ZN(new_n602));
  XNOR2_X1  g177(.A(G299), .B(KEYINPUT78), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(G297));
  OAI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(G280));
  AND2_X1   g180(.A1(new_n592), .A2(new_n596), .ZN(new_n606));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G860), .ZN(G148));
  NOR2_X1   g183(.A1(new_n597), .A2(G559), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n543), .A2(new_n598), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT11), .Z(G282));
  INV_X1    g188(.A(new_n612), .ZN(G323));
  OAI21_X1  g189(.A(KEYINPUT12), .B1(new_n477), .B2(new_n464), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT12), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n463), .A2(new_n616), .A3(G2104), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  INV_X1    g194(.A(G2100), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  MUX2_X1   g197(.A(G99), .B(G111), .S(G2105), .Z(new_n623));
  AOI22_X1  g198(.A1(G123), .A2(new_n473), .B1(new_n623), .B2(G2104), .ZN(new_n624));
  INV_X1    g199(.A(G135), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(new_n477), .ZN(new_n626));
  INV_X1    g201(.A(G2096), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n621), .A2(new_n622), .A3(new_n628), .ZN(G156));
  INV_X1    g204(.A(KEYINPUT14), .ZN(new_n630));
  XOR2_X1   g205(.A(KEYINPUT15), .B(G2435), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2427), .ZN(new_n633));
  INV_X1    g208(.A(G2430), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n630), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(new_n634), .B2(new_n633), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n636), .A2(new_n642), .ZN(new_n644));
  AND3_X1   g219(.A1(new_n643), .A2(G14), .A3(new_n644), .ZN(G401));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2072), .B(G2078), .Z(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  NOR3_X1   g225(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT18), .ZN(new_n652));
  INV_X1    g227(.A(new_n648), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT17), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n649), .B1(new_n655), .B2(new_n646), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(new_n647), .B2(new_n654), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n647), .A2(new_n650), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n653), .B1(new_n658), .B2(KEYINPUT17), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n652), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(new_n627), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2100), .ZN(G227));
  XOR2_X1   g237(.A(G1971), .B(G1976), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1956), .B(G2474), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1961), .B(G1966), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT80), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT79), .B(KEYINPUT20), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n665), .A2(new_n666), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n664), .A2(new_n667), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n664), .B2(new_n672), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1981), .B(G1986), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT81), .ZN(new_n679));
  XOR2_X1   g254(.A(G1991), .B(G1996), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n677), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G229));
  NOR2_X1   g258(.A1(G6), .A2(G16), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n579), .B2(G16), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT85), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT32), .B(G1981), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G23), .ZN(new_n691));
  INV_X1    g266(.A(G288), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT33), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(G16), .A2(G22), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G166), .B2(G16), .ZN(new_n697));
  INV_X1    g272(.A(G1971), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND4_X1  g274(.A1(new_n688), .A2(new_n689), .A3(new_n695), .A4(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT84), .B(KEYINPUT34), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(G24), .B(G290), .S(G16), .Z(new_n703));
  NOR2_X1   g278(.A1(new_n703), .A2(G1986), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n703), .A2(G1986), .ZN(new_n705));
  MUX2_X1   g280(.A(G95), .B(G107), .S(G2105), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G2104), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT82), .Z(new_n708));
  AOI22_X1  g283(.A1(G119), .A2(new_n473), .B1(new_n463), .B2(G131), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  MUX2_X1   g285(.A(G25), .B(new_n710), .S(G29), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT83), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT35), .B(G1991), .Z(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n712), .B(new_n714), .ZN(new_n715));
  NOR4_X1   g290(.A1(new_n702), .A2(new_n704), .A3(new_n705), .A4(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT36), .Z(new_n717));
  NOR2_X1   g292(.A1(G16), .A2(G19), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n543), .B2(G16), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT87), .B(G1341), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(G4), .A2(G16), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n606), .B2(G16), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT86), .B(G1348), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(G27), .A2(G29), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G164), .B2(G29), .ZN(new_n727));
  AOI211_X1 g302(.A(new_n721), .B(new_n725), .C1(G2078), .C2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G29), .A2(G35), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G162), .B2(G29), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT29), .Z(new_n731));
  INV_X1    g306(.A(G2090), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(KEYINPUT94), .ZN(new_n734));
  NAND3_X1  g309(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT26), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G105), .B2(new_n465), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n463), .A2(G141), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n473), .A2(G129), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT89), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G29), .ZN(new_n742));
  NOR2_X1   g317(.A1(G29), .A2(G32), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(KEYINPUT90), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(KEYINPUT90), .B2(new_n742), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT27), .B(G1996), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n690), .A2(G21), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G168), .B2(new_n690), .ZN(new_n749));
  INV_X1    g324(.A(G1966), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n728), .A2(new_n734), .A3(new_n747), .A4(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G29), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G26), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT28), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n463), .A2(G140), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT88), .Z(new_n757));
  MUX2_X1   g332(.A(G104), .B(G116), .S(G2105), .Z(new_n758));
  AOI22_X1  g333(.A1(G128), .A2(new_n473), .B1(new_n758), .B2(G2104), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n755), .B1(new_n760), .B2(G29), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2067), .ZN(new_n762));
  NOR2_X1   g337(.A1(G5), .A2(G16), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT92), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G171), .B2(G16), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n762), .B1(new_n765), .B2(G1961), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n753), .A2(G33), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n484), .A2(G127), .ZN(new_n768));
  NAND2_X1  g343(.A1(G115), .A2(G2104), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n472), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n465), .A2(G103), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT25), .ZN(new_n772));
  AOI211_X1 g347(.A(new_n770), .B(new_n772), .C1(G139), .C2(new_n463), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n767), .B1(new_n773), .B2(new_n753), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2072), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT31), .B(G11), .Z(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT30), .B(G28), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n776), .B1(new_n753), .B2(new_n777), .ZN(new_n778));
  OAI221_X1 g353(.A(new_n778), .B1(new_n753), .B2(new_n626), .C1(new_n727), .C2(G2078), .ZN(new_n779));
  OR2_X1    g354(.A1(KEYINPUT24), .A2(G34), .ZN(new_n780));
  NAND2_X1  g355(.A1(KEYINPUT24), .A2(G34), .ZN(new_n781));
  AOI21_X1  g356(.A(G29), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G160), .B2(G29), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G2084), .ZN(new_n784));
  OR3_X1    g359(.A1(new_n775), .A2(new_n779), .A3(new_n784), .ZN(new_n785));
  AOI211_X1 g360(.A(new_n766), .B(new_n785), .C1(new_n732), .C2(new_n731), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n765), .A2(G1961), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT93), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n690), .A2(G20), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT23), .ZN(new_n790));
  INV_X1    g365(.A(G299), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(new_n690), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(G1956), .Z(new_n793));
  NAND3_X1  g368(.A1(new_n786), .A2(new_n788), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n745), .A2(new_n746), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT91), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(KEYINPUT94), .B2(new_n733), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n752), .A2(new_n794), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n717), .A2(new_n798), .ZN(G150));
  INV_X1    g374(.A(G150), .ZN(G311));
  NAND2_X1  g375(.A1(new_n606), .A2(G559), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT95), .ZN(new_n802));
  INV_X1    g377(.A(G55), .ZN(new_n803));
  INV_X1    g378(.A(G93), .ZN(new_n804));
  OAI22_X1  g379(.A1(new_n803), .A2(new_n498), .B1(new_n504), .B2(new_n804), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(new_n508), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n543), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n543), .A2(new_n808), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT38), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n802), .B(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT39), .ZN(new_n814));
  AOI21_X1  g389(.A(G860), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n814), .B2(new_n813), .ZN(new_n816));
  INV_X1    g391(.A(new_n808), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G860), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT37), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n816), .A2(new_n819), .ZN(G145));
  MUX2_X1   g395(.A(G106), .B(G118), .S(G2105), .Z(new_n821));
  AOI22_X1  g396(.A1(G130), .A2(new_n473), .B1(new_n821), .B2(G2104), .ZN(new_n822));
  INV_X1    g397(.A(G142), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(new_n477), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n618), .B(new_n824), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(new_n710), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT96), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n483), .A2(new_n486), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(new_n491), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n827), .B1(new_n483), .B2(new_n486), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n760), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n826), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n741), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(new_n773), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n773), .B2(new_n740), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n833), .B(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(G162), .B(G160), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n626), .ZN(new_n839));
  AOI21_X1  g414(.A(G37), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n839), .B2(new_n837), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g417(.A(G290), .B(G288), .ZN(new_n843));
  XNOR2_X1  g418(.A(G305), .B(G166), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n843), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT42), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n606), .B1(new_n556), .B2(new_n557), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT41), .ZN(new_n849));
  INV_X1    g424(.A(new_n557), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n597), .A2(new_n850), .A3(new_n555), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n848), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(KEYINPUT97), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT97), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n848), .A2(new_n854), .A3(new_n849), .A4(new_n851), .ZN(new_n855));
  NOR2_X1   g430(.A1(G299), .A2(new_n597), .ZN(new_n856));
  INV_X1    g431(.A(new_n851), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT41), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n853), .A2(new_n855), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n811), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(G559), .B2(new_n597), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n609), .A2(new_n811), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  AND4_X1   g439(.A1(new_n848), .A2(new_n861), .A3(new_n851), .A4(new_n862), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n847), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  AOI211_X1 g442(.A(KEYINPUT42), .B(new_n865), .C1(new_n859), .C2(new_n863), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n846), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n863), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n849), .B1(new_n848), .B2(new_n851), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n871), .B1(KEYINPUT97), .B2(new_n852), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n870), .B1(new_n872), .B2(new_n855), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT42), .B1(new_n873), .B2(new_n865), .ZN(new_n874));
  INV_X1    g449(.A(new_n846), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n864), .A2(new_n847), .A3(new_n866), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n598), .B1(new_n869), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n817), .A2(G868), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(G295));
  NAND2_X1  g455(.A1(new_n869), .A2(new_n877), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(G868), .ZN(new_n882));
  INV_X1    g457(.A(new_n879), .ZN(new_n883));
  AOI21_X1  g458(.A(KEYINPUT98), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT98), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n878), .A2(new_n885), .A3(new_n879), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n884), .A2(new_n886), .ZN(G331));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n858), .A2(new_n852), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT99), .ZN(new_n890));
  AOI21_X1  g465(.A(G286), .B1(new_n561), .B2(new_n562), .ZN(new_n891));
  NOR2_X1   g466(.A1(G168), .A2(G171), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n562), .ZN(new_n894));
  OAI21_X1  g469(.A(G168), .B1(new_n894), .B2(new_n560), .ZN(new_n895));
  NAND3_X1  g470(.A1(G286), .A2(new_n536), .A3(new_n533), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(KEYINPUT99), .A3(new_n896), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n893), .A2(new_n811), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n811), .B1(new_n893), .B2(new_n897), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n889), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n898), .A2(new_n899), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n856), .A2(new_n857), .ZN(new_n903));
  AOI22_X1  g478(.A1(new_n900), .A2(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n900), .A2(new_n901), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n846), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n897), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT99), .B1(new_n895), .B2(new_n896), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n860), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n893), .A2(new_n897), .A3(new_n811), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n903), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n859), .B1(new_n898), .B2(new_n899), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n909), .A2(KEYINPUT100), .A3(new_n903), .A4(new_n910), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n913), .A2(new_n846), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G37), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT43), .B1(new_n906), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n913), .A2(new_n915), .A3(new_n914), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n875), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n921), .A2(new_n922), .A3(new_n917), .A4(new_n916), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n888), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n922), .B1(new_n906), .B2(new_n918), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n921), .A2(KEYINPUT43), .A3(new_n917), .A4(new_n916), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT44), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n924), .A2(new_n927), .ZN(G397));
  NAND2_X1  g503(.A1(new_n487), .A2(KEYINPUT96), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(new_n491), .A3(new_n828), .ZN(new_n930));
  INV_X1    g505(.A(G1384), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XOR2_X1   g507(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n466), .A2(new_n470), .A3(G40), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n740), .ZN(new_n938));
  INV_X1    g513(.A(G1996), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n940), .B(KEYINPUT104), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n760), .B(G2067), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(KEYINPUT105), .A3(new_n937), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n937), .A2(new_n939), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n944), .A2(new_n834), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT105), .B1(new_n942), .B2(new_n937), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n941), .A2(new_n943), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n710), .A2(new_n714), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n713), .B1(new_n708), .B2(new_n709), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n937), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(G290), .A2(G1986), .ZN(new_n953));
  NOR2_X1   g528(.A1(G290), .A2(G1986), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n937), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT103), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT125), .ZN(new_n958));
  INV_X1    g533(.A(G8), .ZN(new_n959));
  OR3_X1    g534(.A1(G168), .A2(KEYINPUT120), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT120), .B1(G168), .B2(new_n959), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT50), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n963), .B(new_n931), .C1(new_n829), .C2(new_n830), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT106), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT106), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n930), .A2(new_n966), .A3(new_n963), .A4(new_n931), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n969));
  INV_X1    g544(.A(G2084), .ZN(new_n970));
  AOI21_X1  g545(.A(G1384), .B1(new_n487), .B2(new_n491), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n935), .B1(new_n971), .B2(new_n963), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n968), .A2(new_n969), .A3(new_n970), .A4(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n831), .A2(G1384), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n975), .A2(KEYINPUT45), .ZN(new_n976));
  INV_X1    g551(.A(new_n971), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n935), .B1(new_n977), .B2(new_n933), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n750), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n974), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n972), .B1(new_n965), .B2(new_n967), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n969), .B1(new_n981), .B2(new_n970), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n962), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT121), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n968), .A2(new_n970), .A3(new_n973), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT113), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(new_n974), .A3(new_n979), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT121), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(new_n988), .A3(new_n962), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n984), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n962), .B1(new_n987), .B2(G8), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT122), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(G8), .B1(new_n980), .B2(new_n982), .ZN(new_n995));
  INV_X1    g570(.A(new_n962), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n997), .A2(KEYINPUT122), .A3(KEYINPUT51), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n990), .B1(new_n994), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT62), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n958), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1981), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n571), .A2(new_n577), .A3(new_n1002), .A4(new_n572), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n1003), .B(KEYINPUT109), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n578), .B1(new_n573), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n571), .A2(KEYINPUT110), .A3(new_n572), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1002), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1005), .A2(new_n1010), .A3(KEYINPUT49), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT49), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(new_n1004), .B2(new_n1009), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n930), .A2(new_n931), .A3(new_n935), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1014), .A2(G8), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1011), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n567), .A2(G1976), .A3(new_n568), .A4(new_n569), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT108), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1019), .A2(G8), .A3(new_n1014), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT52), .ZN(new_n1021));
  INV_X1    g596(.A(G1976), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(G288), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1015), .A2(new_n1019), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1016), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n930), .A2(KEYINPUT45), .A3(new_n931), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n977), .A2(new_n933), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(new_n935), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n698), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n971), .A2(new_n963), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT112), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n971), .A2(new_n1032), .A3(new_n963), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n936), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n932), .A2(KEYINPUT50), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1029), .B1(new_n1036), .B2(G2090), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(G8), .ZN(new_n1038));
  OAI211_X1 g613(.A(G303), .B(G8), .C1(KEYINPUT107), .C2(KEYINPUT55), .ZN(new_n1039));
  NAND2_X1  g614(.A1(KEYINPUT107), .A2(KEYINPUT55), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n1039), .B(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1025), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n981), .A2(new_n732), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n959), .B1(new_n1044), .B2(new_n1029), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n1041), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT45), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n978), .B1(new_n1047), .B2(new_n932), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(G2078), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1049), .B1(new_n1028), .B2(G2078), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1051), .B(new_n1052), .C1(G1961), .C2(new_n981), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1053), .A2(new_n563), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1043), .A2(new_n1046), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n999), .B2(new_n1000), .ZN(new_n1056));
  INV_X1    g631(.A(new_n990), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT51), .B1(new_n997), .B2(KEYINPUT122), .ZN(new_n1058));
  AOI211_X1 g633(.A(new_n993), .B(new_n991), .C1(new_n995), .C2(new_n996), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1060), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1001), .A2(new_n1056), .A3(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n934), .A2(new_n935), .A3(new_n1026), .A4(new_n1050), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1052), .B(new_n1063), .C1(G1961), .C2(new_n981), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(G171), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT54), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1053), .A2(new_n563), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1043), .B(new_n1046), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n981), .A2(G1348), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1014), .A2(KEYINPUT119), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n930), .A2(new_n935), .A3(new_n1071), .A4(new_n931), .ZN(new_n1072));
  AOI21_X1  g647(.A(G2067), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  NOR4_X1   g648(.A1(new_n1069), .A2(new_n1073), .A3(KEYINPUT60), .A4(new_n597), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT117), .B(G1956), .Z(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1076));
  XOR2_X1   g651(.A(KEYINPUT56), .B(G2072), .Z(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1026), .A2(new_n935), .A3(new_n1027), .A4(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  XOR2_X1   g655(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n551), .A2(new_n554), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n551), .B2(new_n554), .ZN(new_n1084));
  OAI22_X1  g659(.A1(new_n1076), .A2(new_n1080), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1087), .A2(new_n935), .A3(new_n1035), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1086), .B(new_n1079), .C1(new_n1088), .C2(new_n1075), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT61), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1074), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1093));
  OAI221_X1 g668(.A(new_n597), .B1(new_n981), .B2(G1348), .C1(new_n1093), .C2(G2067), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n606), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT60), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1085), .A2(new_n1089), .A3(KEYINPUT61), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT58), .B(G1341), .ZN(new_n1100));
  OAI22_X1  g675(.A1(new_n1099), .A2(new_n1100), .B1(new_n1028), .B2(G1996), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n543), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT59), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1101), .A2(new_n1104), .A3(new_n543), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1092), .A2(new_n1097), .A3(new_n1098), .A4(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1089), .B(new_n606), .C1(new_n1073), .C2(new_n1069), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1108), .A2(new_n1085), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1068), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT123), .B(KEYINPUT54), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1064), .A2(new_n563), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1111), .B1(new_n1054), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT124), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1115), .B(new_n1111), .C1(new_n1054), .C2(new_n1112), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1110), .A2(new_n1060), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT115), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1045), .A2(new_n1119), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n981), .A2(new_n732), .B1(new_n1028), .B2(new_n698), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT115), .B1(new_n1121), .B2(new_n959), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n1042), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT116), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1025), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1041), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT116), .B1(new_n1128), .B2(new_n1025), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1046), .A2(KEYINPUT63), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n987), .A2(G8), .A3(G168), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1127), .A2(new_n1129), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT63), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1135), .A2(new_n1046), .A3(new_n1126), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1134), .B1(new_n1136), .B2(new_n1131), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT114), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT114), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1139), .B(new_n1134), .C1(new_n1136), .C2(new_n1131), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1133), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1046), .A2(new_n1025), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1016), .A2(new_n1022), .A3(new_n692), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n1005), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n1144), .A2(KEYINPUT111), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1015), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1146), .B1(new_n1144), .B2(KEYINPUT111), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1142), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1118), .A2(new_n1141), .A3(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n957), .B1(new_n1062), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n937), .B1(new_n942), .B2(new_n740), .ZN(new_n1151));
  XOR2_X1   g726(.A(new_n1151), .B(KEYINPUT127), .Z(new_n1152));
  XNOR2_X1  g727(.A(new_n944), .B(KEYINPUT46), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1154), .B(KEYINPUT47), .Z(new_n1155));
  INV_X1    g730(.A(new_n937), .ZN(new_n1156));
  XOR2_X1   g731(.A(new_n949), .B(KEYINPUT126), .Z(new_n1157));
  NAND2_X1  g732(.A1(new_n948), .A2(new_n1157), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n760), .A2(G2067), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1156), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n954), .A2(new_n937), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT48), .ZN(new_n1162));
  AOI211_X1 g737(.A(new_n1155), .B(new_n1160), .C1(new_n952), .C2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1150), .A2(new_n1163), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g739(.A(G319), .ZN(new_n1166));
  NOR3_X1   g740(.A1(G227), .A2(G401), .A3(new_n1166), .ZN(new_n1167));
  AND3_X1   g741(.A1(new_n841), .A2(new_n682), .A3(new_n1167), .ZN(new_n1168));
  NAND3_X1  g742(.A1(new_n1168), .A2(new_n925), .A3(new_n926), .ZN(G225));
  INV_X1    g743(.A(G225), .ZN(G308));
endmodule


