

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U549 ( .A1(n757), .A2(n756), .ZN(n759) );
  XOR2_X1 U550 ( .A(KEYINPUT29), .B(n658), .Z(n516) );
  INV_X1 U551 ( .A(KEYINPUT97), .ZN(n632) );
  XNOR2_X1 U552 ( .A(n633), .B(n632), .ZN(n634) );
  INV_X1 U553 ( .A(n642), .ZN(n643) );
  XNOR2_X1 U554 ( .A(KEYINPUT31), .B(KEYINPUT101), .ZN(n602) );
  XNOR2_X1 U555 ( .A(n603), .B(n602), .ZN(n667) );
  AND2_X1 U556 ( .A1(n706), .A2(n987), .ZN(n675) );
  INV_X1 U557 ( .A(KEYINPUT103), .ZN(n680) );
  NAND2_X1 U558 ( .A1(n590), .A2(n690), .ZN(n642) );
  NOR2_X2 U559 ( .A1(G2104), .A2(n542), .ZN(n872) );
  NOR2_X1 U560 ( .A1(G2104), .A2(G2105), .ZN(n535) );
  NOR2_X1 U561 ( .A1(G651), .A2(n570), .ZN(n790) );
  INV_X1 U562 ( .A(KEYINPUT40), .ZN(n758) );
  NOR2_X1 U563 ( .A1(G543), .A2(G651), .ZN(n791) );
  NAND2_X1 U564 ( .A1(n791), .A2(G89), .ZN(n517) );
  XNOR2_X1 U565 ( .A(n517), .B(KEYINPUT4), .ZN(n519) );
  XOR2_X1 U566 ( .A(G543), .B(KEYINPUT0), .Z(n570) );
  XNOR2_X1 U567 ( .A(KEYINPUT65), .B(G651), .ZN(n521) );
  NOR2_X1 U568 ( .A1(n570), .A2(n521), .ZN(n787) );
  NAND2_X1 U569 ( .A1(G76), .A2(n787), .ZN(n518) );
  NAND2_X1 U570 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U571 ( .A(KEYINPUT5), .B(n520), .ZN(n528) );
  NAND2_X1 U572 ( .A1(n790), .A2(G51), .ZN(n524) );
  NOR2_X1 U573 ( .A1(G543), .A2(n521), .ZN(n522) );
  XOR2_X1 U574 ( .A(KEYINPUT1), .B(n522), .Z(n786) );
  NAND2_X1 U575 ( .A1(G63), .A2(n786), .ZN(n523) );
  NAND2_X1 U576 ( .A1(n524), .A2(n523), .ZN(n526) );
  XOR2_X1 U577 ( .A(KEYINPUT6), .B(KEYINPUT72), .Z(n525) );
  XNOR2_X1 U578 ( .A(n526), .B(n525), .ZN(n527) );
  NAND2_X1 U579 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U580 ( .A(KEYINPUT7), .B(n529), .ZN(G168) );
  INV_X1 U581 ( .A(G2105), .ZN(n542) );
  NAND2_X1 U582 ( .A1(n872), .A2(G125), .ZN(n533) );
  NAND2_X1 U583 ( .A1(G101), .A2(G2104), .ZN(n530) );
  OR2_X1 U584 ( .A1(n530), .A2(G2105), .ZN(n531) );
  XOR2_X1 U585 ( .A(KEYINPUT23), .B(n531), .Z(n532) );
  NAND2_X1 U586 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U587 ( .A(n534), .B(KEYINPUT64), .ZN(n539) );
  XOR2_X2 U588 ( .A(KEYINPUT17), .B(n535), .Z(n876) );
  NAND2_X1 U589 ( .A1(G137), .A2(n876), .ZN(n537) );
  AND2_X1 U590 ( .A1(G2104), .A2(G2105), .ZN(n873) );
  NAND2_X1 U591 ( .A1(G113), .A2(n873), .ZN(n536) );
  NAND2_X1 U592 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U593 ( .A1(n539), .A2(n538), .ZN(G160) );
  NAND2_X1 U594 ( .A1(n876), .A2(G138), .ZN(n546) );
  NAND2_X1 U595 ( .A1(G126), .A2(n872), .ZN(n541) );
  NAND2_X1 U596 ( .A1(G114), .A2(n873), .ZN(n540) );
  AND2_X1 U597 ( .A1(n541), .A2(n540), .ZN(n544) );
  AND2_X1 U598 ( .A1(n542), .A2(G2104), .ZN(n877) );
  NAND2_X1 U599 ( .A1(G102), .A2(n877), .ZN(n543) );
  AND2_X1 U600 ( .A1(n544), .A2(n543), .ZN(n545) );
  AND2_X1 U601 ( .A1(n546), .A2(n545), .ZN(G164) );
  NAND2_X1 U602 ( .A1(n790), .A2(G52), .ZN(n548) );
  NAND2_X1 U603 ( .A1(G64), .A2(n786), .ZN(n547) );
  NAND2_X1 U604 ( .A1(n548), .A2(n547), .ZN(n553) );
  NAND2_X1 U605 ( .A1(n791), .A2(G90), .ZN(n550) );
  NAND2_X1 U606 ( .A1(G77), .A2(n787), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U608 ( .A(KEYINPUT9), .B(n551), .Z(n552) );
  NOR2_X1 U609 ( .A1(n553), .A2(n552), .ZN(G171) );
  NAND2_X1 U610 ( .A1(n790), .A2(G50), .ZN(n560) );
  NAND2_X1 U611 ( .A1(G62), .A2(n786), .ZN(n555) );
  NAND2_X1 U612 ( .A1(G75), .A2(n787), .ZN(n554) );
  NAND2_X1 U613 ( .A1(n555), .A2(n554), .ZN(n558) );
  NAND2_X1 U614 ( .A1(n791), .A2(G88), .ZN(n556) );
  XOR2_X1 U615 ( .A(KEYINPUT80), .B(n556), .Z(n557) );
  NOR2_X1 U616 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U617 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U618 ( .A(KEYINPUT81), .B(n561), .Z(G303) );
  NAND2_X1 U619 ( .A1(G53), .A2(n790), .ZN(n563) );
  NAND2_X1 U620 ( .A1(G91), .A2(n791), .ZN(n562) );
  NAND2_X1 U621 ( .A1(n563), .A2(n562), .ZN(n566) );
  NAND2_X1 U622 ( .A1(n786), .A2(G65), .ZN(n564) );
  XOR2_X1 U623 ( .A(KEYINPUT66), .B(n564), .Z(n565) );
  NOR2_X1 U624 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U625 ( .A1(G78), .A2(n787), .ZN(n567) );
  NAND2_X1 U626 ( .A1(n568), .A2(n567), .ZN(G299) );
  XNOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .ZN(n569) );
  XNOR2_X1 U628 ( .A(n569), .B(KEYINPUT73), .ZN(G286) );
  NAND2_X1 U629 ( .A1(G87), .A2(n570), .ZN(n572) );
  NAND2_X1 U630 ( .A1(G74), .A2(G651), .ZN(n571) );
  NAND2_X1 U631 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U632 ( .A1(n786), .A2(n573), .ZN(n575) );
  NAND2_X1 U633 ( .A1(n790), .A2(G49), .ZN(n574) );
  NAND2_X1 U634 ( .A1(n575), .A2(n574), .ZN(G288) );
  NAND2_X1 U635 ( .A1(G48), .A2(n790), .ZN(n577) );
  NAND2_X1 U636 ( .A1(G86), .A2(n791), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n577), .A2(n576), .ZN(n581) );
  NAND2_X1 U638 ( .A1(n787), .A2(G73), .ZN(n578) );
  XNOR2_X1 U639 ( .A(n578), .B(KEYINPUT2), .ZN(n579) );
  XNOR2_X1 U640 ( .A(n579), .B(KEYINPUT79), .ZN(n580) );
  NOR2_X1 U641 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U642 ( .A1(G61), .A2(n786), .ZN(n582) );
  NAND2_X1 U643 ( .A1(n583), .A2(n582), .ZN(G305) );
  INV_X1 U644 ( .A(G303), .ZN(G166) );
  NAND2_X1 U645 ( .A1(G60), .A2(n786), .ZN(n585) );
  NAND2_X1 U646 ( .A1(G72), .A2(n787), .ZN(n584) );
  NAND2_X1 U647 ( .A1(n585), .A2(n584), .ZN(n589) );
  NAND2_X1 U648 ( .A1(G47), .A2(n790), .ZN(n587) );
  NAND2_X1 U649 ( .A1(G85), .A2(n791), .ZN(n586) );
  NAND2_X1 U650 ( .A1(n587), .A2(n586), .ZN(n588) );
  OR2_X1 U651 ( .A1(n589), .A2(n588), .ZN(G290) );
  AND2_X1 U652 ( .A1(G160), .A2(G40), .ZN(n590) );
  NOR2_X1 U653 ( .A1(G164), .A2(G1384), .ZN(n690) );
  NOR2_X1 U654 ( .A1(G2084), .A2(n642), .ZN(n669) );
  NAND2_X1 U655 ( .A1(G8), .A2(n642), .ZN(n713) );
  NOR2_X1 U656 ( .A1(G1966), .A2(n713), .ZN(n592) );
  INV_X1 U657 ( .A(KEYINPUT94), .ZN(n591) );
  XNOR2_X1 U658 ( .A(n592), .B(n591), .ZN(n673) );
  NAND2_X1 U659 ( .A1(n673), .A2(G8), .ZN(n593) );
  NOR2_X1 U660 ( .A1(n669), .A2(n593), .ZN(n595) );
  XOR2_X1 U661 ( .A(KEYINPUT30), .B(KEYINPUT100), .Z(n594) );
  XNOR2_X1 U662 ( .A(n595), .B(n594), .ZN(n596) );
  NOR2_X1 U663 ( .A1(G168), .A2(n596), .ZN(n601) );
  XOR2_X1 U664 ( .A(KEYINPUT25), .B(G2078), .Z(n917) );
  NOR2_X1 U665 ( .A1(n917), .A2(n642), .ZN(n598) );
  NOR2_X1 U666 ( .A1(n643), .A2(G1961), .ZN(n597) );
  NOR2_X1 U667 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U668 ( .A(KEYINPUT95), .B(n599), .ZN(n610) );
  NOR2_X1 U669 ( .A1(G171), .A2(n610), .ZN(n600) );
  NOR2_X1 U670 ( .A1(n601), .A2(n600), .ZN(n603) );
  INV_X1 U671 ( .A(G8), .ZN(n609) );
  NOR2_X1 U672 ( .A1(G1971), .A2(n713), .ZN(n605) );
  NOR2_X1 U673 ( .A1(G2090), .A2(n642), .ZN(n604) );
  NOR2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U675 ( .A(n606), .B(KEYINPUT102), .ZN(n607) );
  NAND2_X1 U676 ( .A1(n607), .A2(G303), .ZN(n608) );
  OR2_X1 U677 ( .A1(n609), .A2(n608), .ZN(n661) );
  AND2_X1 U678 ( .A1(n667), .A2(n661), .ZN(n660) );
  NAND2_X1 U679 ( .A1(n610), .A2(G171), .ZN(n659) );
  NAND2_X1 U680 ( .A1(n643), .A2(G2072), .ZN(n611) );
  XNOR2_X1 U681 ( .A(n611), .B(KEYINPUT27), .ZN(n613) );
  AND2_X1 U682 ( .A1(G1956), .A2(n642), .ZN(n612) );
  NOR2_X1 U683 ( .A1(n613), .A2(n612), .ZN(n653) );
  INV_X1 U684 ( .A(G299), .ZN(n989) );
  NOR2_X1 U685 ( .A1(n653), .A2(n989), .ZN(n615) );
  XOR2_X1 U686 ( .A(KEYINPUT96), .B(KEYINPUT28), .Z(n614) );
  XNOR2_X1 U687 ( .A(n615), .B(n614), .ZN(n657) );
  NAND2_X1 U688 ( .A1(n790), .A2(G43), .ZN(n616) );
  XNOR2_X1 U689 ( .A(KEYINPUT69), .B(n616), .ZN(n623) );
  NAND2_X1 U690 ( .A1(n791), .A2(G81), .ZN(n617) );
  XNOR2_X1 U691 ( .A(n617), .B(KEYINPUT12), .ZN(n619) );
  NAND2_X1 U692 ( .A1(G68), .A2(n787), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U694 ( .A(KEYINPUT68), .B(n620), .Z(n621) );
  XNOR2_X1 U695 ( .A(KEYINPUT13), .B(n621), .ZN(n622) );
  NOR2_X1 U696 ( .A1(n623), .A2(n622), .ZN(n627) );
  XOR2_X1 U697 ( .A(KEYINPUT67), .B(KEYINPUT14), .Z(n625) );
  NAND2_X1 U698 ( .A1(G56), .A2(n786), .ZN(n624) );
  XNOR2_X1 U699 ( .A(n625), .B(n624), .ZN(n626) );
  NAND2_X1 U700 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U701 ( .A(n628), .B(KEYINPUT70), .ZN(n996) );
  NAND2_X1 U702 ( .A1(G1996), .A2(n643), .ZN(n629) );
  XNOR2_X1 U703 ( .A(n629), .B(KEYINPUT26), .ZN(n631) );
  NAND2_X1 U704 ( .A1(G1341), .A2(n642), .ZN(n630) );
  NAND2_X1 U705 ( .A1(n631), .A2(n630), .ZN(n633) );
  NOR2_X1 U706 ( .A1(n996), .A2(n634), .ZN(n648) );
  NAND2_X1 U707 ( .A1(G66), .A2(n786), .ZN(n636) );
  NAND2_X1 U708 ( .A1(G79), .A2(n787), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U710 ( .A1(G54), .A2(n790), .ZN(n638) );
  NAND2_X1 U711 ( .A1(G92), .A2(n791), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U713 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U714 ( .A(KEYINPUT15), .B(n641), .Z(n998) );
  NAND2_X1 U715 ( .A1(G1348), .A2(n642), .ZN(n645) );
  NAND2_X1 U716 ( .A1(G2067), .A2(n643), .ZN(n644) );
  NAND2_X1 U717 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U718 ( .A(KEYINPUT98), .B(n646), .Z(n649) );
  OR2_X1 U719 ( .A1(n998), .A2(n649), .ZN(n647) );
  NAND2_X1 U720 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U721 ( .A1(n649), .A2(n998), .ZN(n650) );
  NAND2_X1 U722 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U723 ( .A(n652), .B(KEYINPUT99), .ZN(n655) );
  NAND2_X1 U724 ( .A1(n653), .A2(n989), .ZN(n654) );
  NAND2_X1 U725 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U726 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U727 ( .A1(n659), .A2(n516), .ZN(n668) );
  NAND2_X1 U728 ( .A1(n660), .A2(n668), .ZN(n665) );
  INV_X1 U729 ( .A(n661), .ZN(n663) );
  AND2_X1 U730 ( .A1(G286), .A2(G8), .ZN(n662) );
  OR2_X1 U731 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U732 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U733 ( .A(n666), .B(KEYINPUT32), .ZN(n707) );
  NAND2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n672) );
  NAND2_X1 U735 ( .A1(G8), .A2(n669), .ZN(n670) );
  XOR2_X1 U736 ( .A(KEYINPUT93), .B(n670), .Z(n671) );
  AND2_X1 U737 ( .A1(n672), .A2(n671), .ZN(n674) );
  NAND2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n706) );
  NAND2_X1 U739 ( .A1(G1976), .A2(G288), .ZN(n987) );
  NAND2_X1 U740 ( .A1(n707), .A2(n675), .ZN(n679) );
  INV_X1 U741 ( .A(n987), .ZN(n677) );
  NOR2_X1 U742 ( .A1(G1976), .A2(G288), .ZN(n685) );
  NOR2_X1 U743 ( .A1(G1971), .A2(G303), .ZN(n676) );
  NOR2_X1 U744 ( .A1(n685), .A2(n676), .ZN(n995) );
  OR2_X1 U745 ( .A1(n677), .A2(n995), .ZN(n678) );
  AND2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n681) );
  XNOR2_X1 U747 ( .A(n681), .B(n680), .ZN(n682) );
  NOR2_X1 U748 ( .A1(n682), .A2(n713), .ZN(n683) );
  NOR2_X1 U749 ( .A1(KEYINPUT33), .A2(n683), .ZN(n684) );
  XNOR2_X1 U750 ( .A(n684), .B(KEYINPUT104), .ZN(n688) );
  NAND2_X1 U751 ( .A1(n685), .A2(KEYINPUT33), .ZN(n686) );
  NOR2_X1 U752 ( .A1(n713), .A2(n686), .ZN(n687) );
  NOR2_X1 U753 ( .A1(n688), .A2(n687), .ZN(n703) );
  XOR2_X1 U754 ( .A(G1981), .B(G305), .Z(n1006) );
  NAND2_X1 U755 ( .A1(G160), .A2(G40), .ZN(n689) );
  NOR2_X1 U756 ( .A1(n690), .A2(n689), .ZN(n752) );
  NAND2_X1 U757 ( .A1(G140), .A2(n876), .ZN(n692) );
  NAND2_X1 U758 ( .A1(G104), .A2(n877), .ZN(n691) );
  NAND2_X1 U759 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U760 ( .A(KEYINPUT34), .B(n693), .ZN(n698) );
  NAND2_X1 U761 ( .A1(G128), .A2(n872), .ZN(n695) );
  NAND2_X1 U762 ( .A1(G116), .A2(n873), .ZN(n694) );
  NAND2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U764 ( .A(n696), .B(KEYINPUT35), .Z(n697) );
  NOR2_X1 U765 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U766 ( .A(KEYINPUT36), .B(n699), .Z(n700) );
  XOR2_X1 U767 ( .A(KEYINPUT86), .B(n700), .Z(n891) );
  XNOR2_X1 U768 ( .A(G2067), .B(KEYINPUT37), .ZN(n746) );
  OR2_X1 U769 ( .A1(n891), .A2(n746), .ZN(n701) );
  XNOR2_X1 U770 ( .A(n701), .B(KEYINPUT87), .ZN(n982) );
  NAND2_X1 U771 ( .A1(n752), .A2(n982), .ZN(n744) );
  AND2_X1 U772 ( .A1(n1006), .A2(n744), .ZN(n702) );
  NAND2_X1 U773 ( .A1(n703), .A2(n702), .ZN(n751) );
  NAND2_X1 U774 ( .A1(G8), .A2(G166), .ZN(n704) );
  NOR2_X1 U775 ( .A1(G2090), .A2(n704), .ZN(n705) );
  XNOR2_X1 U776 ( .A(n705), .B(KEYINPUT105), .ZN(n709) );
  NAND2_X1 U777 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U778 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U779 ( .A1(n710), .A2(n713), .ZN(n715) );
  NOR2_X1 U780 ( .A1(G1981), .A2(G305), .ZN(n711) );
  XOR2_X1 U781 ( .A(n711), .B(KEYINPUT24), .Z(n712) );
  OR2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U783 ( .A1(n715), .A2(n714), .ZN(n716) );
  AND2_X1 U784 ( .A1(n744), .A2(n716), .ZN(n749) );
  NAND2_X1 U785 ( .A1(n873), .A2(G117), .ZN(n723) );
  NAND2_X1 U786 ( .A1(G141), .A2(n876), .ZN(n718) );
  NAND2_X1 U787 ( .A1(G129), .A2(n872), .ZN(n717) );
  NAND2_X1 U788 ( .A1(n718), .A2(n717), .ZN(n721) );
  NAND2_X1 U789 ( .A1(n877), .A2(G105), .ZN(n719) );
  XOR2_X1 U790 ( .A(KEYINPUT38), .B(n719), .Z(n720) );
  NOR2_X1 U791 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U792 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U793 ( .A(KEYINPUT91), .B(n724), .Z(n861) );
  NOR2_X1 U794 ( .A1(G1996), .A2(n861), .ZN(n970) );
  NOR2_X1 U795 ( .A1(G1986), .A2(G290), .ZN(n735) );
  NAND2_X1 U796 ( .A1(G95), .A2(n877), .ZN(n725) );
  XNOR2_X1 U797 ( .A(n725), .B(KEYINPUT88), .ZN(n732) );
  NAND2_X1 U798 ( .A1(G119), .A2(n872), .ZN(n727) );
  NAND2_X1 U799 ( .A1(G107), .A2(n873), .ZN(n726) );
  NAND2_X1 U800 ( .A1(n727), .A2(n726), .ZN(n730) );
  NAND2_X1 U801 ( .A1(G131), .A2(n876), .ZN(n728) );
  XNOR2_X1 U802 ( .A(KEYINPUT89), .B(n728), .ZN(n729) );
  NOR2_X1 U803 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U804 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U805 ( .A(KEYINPUT90), .B(n733), .ZN(n860) );
  NOR2_X1 U806 ( .A1(n860), .A2(G1991), .ZN(n734) );
  XNOR2_X1 U807 ( .A(n734), .B(KEYINPUT106), .ZN(n977) );
  NOR2_X1 U808 ( .A1(n735), .A2(n977), .ZN(n736) );
  XNOR2_X1 U809 ( .A(n736), .B(KEYINPUT107), .ZN(n740) );
  NAND2_X1 U810 ( .A1(G1991), .A2(n860), .ZN(n738) );
  NAND2_X1 U811 ( .A1(G1996), .A2(n861), .ZN(n737) );
  NAND2_X1 U812 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U813 ( .A(KEYINPUT92), .B(n739), .Z(n983) );
  NAND2_X1 U814 ( .A1(n740), .A2(n983), .ZN(n741) );
  XOR2_X1 U815 ( .A(KEYINPUT108), .B(n741), .Z(n742) );
  NOR2_X1 U816 ( .A1(n970), .A2(n742), .ZN(n743) );
  XNOR2_X1 U817 ( .A(n743), .B(KEYINPUT39), .ZN(n745) );
  NAND2_X1 U818 ( .A1(n745), .A2(n744), .ZN(n747) );
  NAND2_X1 U819 ( .A1(n891), .A2(n746), .ZN(n967) );
  NAND2_X1 U820 ( .A1(n747), .A2(n967), .ZN(n748) );
  AND2_X1 U821 ( .A1(n748), .A2(n752), .ZN(n755) );
  NOR2_X1 U822 ( .A1(n749), .A2(n755), .ZN(n750) );
  NAND2_X1 U823 ( .A1(n751), .A2(n750), .ZN(n757) );
  XOR2_X1 U824 ( .A(G1986), .B(G290), .Z(n988) );
  NAND2_X1 U825 ( .A1(n988), .A2(n983), .ZN(n753) );
  NAND2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n754) );
  OR2_X1 U827 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U828 ( .A(n759), .B(n758), .ZN(G329) );
  AND2_X1 U829 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U830 ( .A1(G135), .A2(n876), .ZN(n760) );
  XNOR2_X1 U831 ( .A(n760), .B(KEYINPUT76), .ZN(n769) );
  NAND2_X1 U832 ( .A1(G123), .A2(n872), .ZN(n761) );
  XOR2_X1 U833 ( .A(KEYINPUT75), .B(n761), .Z(n762) );
  XNOR2_X1 U834 ( .A(n762), .B(KEYINPUT18), .ZN(n764) );
  NAND2_X1 U835 ( .A1(G111), .A2(n873), .ZN(n763) );
  NAND2_X1 U836 ( .A1(n764), .A2(n763), .ZN(n767) );
  NAND2_X1 U837 ( .A1(G99), .A2(n877), .ZN(n765) );
  XNOR2_X1 U838 ( .A(KEYINPUT77), .B(n765), .ZN(n766) );
  NOR2_X1 U839 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U840 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U841 ( .A(KEYINPUT78), .B(n770), .ZN(n974) );
  XNOR2_X1 U842 ( .A(n974), .B(G2096), .ZN(n771) );
  OR2_X1 U843 ( .A1(G2100), .A2(n771), .ZN(G156) );
  INV_X1 U844 ( .A(G57), .ZN(G237) );
  INV_X1 U845 ( .A(G69), .ZN(G235) );
  INV_X1 U846 ( .A(G108), .ZN(G238) );
  INV_X1 U847 ( .A(G120), .ZN(G236) );
  INV_X1 U848 ( .A(G132), .ZN(G219) );
  INV_X1 U849 ( .A(G82), .ZN(G220) );
  NAND2_X1 U850 ( .A1(G7), .A2(G661), .ZN(n772) );
  XNOR2_X1 U851 ( .A(n772), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U852 ( .A(G223), .ZN(n826) );
  NAND2_X1 U853 ( .A1(n826), .A2(G567), .ZN(n773) );
  XOR2_X1 U854 ( .A(KEYINPUT11), .B(n773), .Z(G234) );
  INV_X1 U855 ( .A(G860), .ZN(n780) );
  OR2_X1 U856 ( .A1(n780), .A2(n996), .ZN(n774) );
  XOR2_X1 U857 ( .A(KEYINPUT71), .B(n774), .Z(G153) );
  INV_X1 U858 ( .A(G171), .ZN(G301) );
  NAND2_X1 U859 ( .A1(G868), .A2(G301), .ZN(n776) );
  OR2_X1 U860 ( .A1(n998), .A2(G868), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n776), .A2(n775), .ZN(G284) );
  INV_X1 U862 ( .A(G868), .ZN(n808) );
  NOR2_X1 U863 ( .A1(G286), .A2(n808), .ZN(n777) );
  XNOR2_X1 U864 ( .A(n777), .B(KEYINPUT74), .ZN(n779) );
  NOR2_X1 U865 ( .A1(G299), .A2(G868), .ZN(n778) );
  NOR2_X1 U866 ( .A1(n779), .A2(n778), .ZN(G297) );
  NAND2_X1 U867 ( .A1(n780), .A2(G559), .ZN(n781) );
  NAND2_X1 U868 ( .A1(n781), .A2(n998), .ZN(n782) );
  XNOR2_X1 U869 ( .A(n782), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U870 ( .A1(n996), .A2(G868), .ZN(n785) );
  NAND2_X1 U871 ( .A1(G868), .A2(n998), .ZN(n783) );
  NOR2_X1 U872 ( .A1(G559), .A2(n783), .ZN(n784) );
  NOR2_X1 U873 ( .A1(n785), .A2(n784), .ZN(G282) );
  NAND2_X1 U874 ( .A1(G67), .A2(n786), .ZN(n789) );
  NAND2_X1 U875 ( .A1(G80), .A2(n787), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n789), .A2(n788), .ZN(n795) );
  NAND2_X1 U877 ( .A1(G55), .A2(n790), .ZN(n793) );
  NAND2_X1 U878 ( .A1(G93), .A2(n791), .ZN(n792) );
  NAND2_X1 U879 ( .A1(n793), .A2(n792), .ZN(n794) );
  OR2_X1 U880 ( .A1(n795), .A2(n794), .ZN(n809) );
  NAND2_X1 U881 ( .A1(n998), .A2(G559), .ZN(n806) );
  XNOR2_X1 U882 ( .A(n996), .B(n806), .ZN(n796) );
  NOR2_X1 U883 ( .A1(G860), .A2(n796), .ZN(n797) );
  XOR2_X1 U884 ( .A(n809), .B(n797), .Z(G145) );
  XNOR2_X1 U885 ( .A(KEYINPUT82), .B(KEYINPUT83), .ZN(n799) );
  XNOR2_X1 U886 ( .A(G288), .B(KEYINPUT19), .ZN(n798) );
  XNOR2_X1 U887 ( .A(n799), .B(n798), .ZN(n800) );
  XNOR2_X1 U888 ( .A(G166), .B(n800), .ZN(n802) );
  XNOR2_X1 U889 ( .A(G290), .B(n989), .ZN(n801) );
  XNOR2_X1 U890 ( .A(n802), .B(n801), .ZN(n803) );
  XOR2_X1 U891 ( .A(n809), .B(n803), .Z(n804) );
  XNOR2_X1 U892 ( .A(n804), .B(G305), .ZN(n805) );
  XNOR2_X1 U893 ( .A(n996), .B(n805), .ZN(n894) );
  XOR2_X1 U894 ( .A(n894), .B(n806), .Z(n807) );
  NAND2_X1 U895 ( .A1(G868), .A2(n807), .ZN(n811) );
  NAND2_X1 U896 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U897 ( .A1(n811), .A2(n810), .ZN(G295) );
  NAND2_X1 U898 ( .A1(G2078), .A2(G2084), .ZN(n812) );
  XOR2_X1 U899 ( .A(KEYINPUT20), .B(n812), .Z(n813) );
  NAND2_X1 U900 ( .A1(G2090), .A2(n813), .ZN(n814) );
  XNOR2_X1 U901 ( .A(KEYINPUT21), .B(n814), .ZN(n815) );
  NAND2_X1 U902 ( .A1(n815), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U903 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U904 ( .A1(G220), .A2(G219), .ZN(n816) );
  XOR2_X1 U905 ( .A(KEYINPUT22), .B(n816), .Z(n817) );
  NOR2_X1 U906 ( .A1(G218), .A2(n817), .ZN(n818) );
  NAND2_X1 U907 ( .A1(G96), .A2(n818), .ZN(n830) );
  NAND2_X1 U908 ( .A1(n830), .A2(G2106), .ZN(n823) );
  NOR2_X1 U909 ( .A1(G236), .A2(G238), .ZN(n820) );
  NOR2_X1 U910 ( .A1(G235), .A2(G237), .ZN(n819) );
  NAND2_X1 U911 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U912 ( .A(KEYINPUT84), .B(n821), .ZN(n831) );
  NAND2_X1 U913 ( .A1(n831), .A2(G567), .ZN(n822) );
  NAND2_X1 U914 ( .A1(n823), .A2(n822), .ZN(n832) );
  NAND2_X1 U915 ( .A1(G661), .A2(G483), .ZN(n824) );
  XOR2_X1 U916 ( .A(KEYINPUT85), .B(n824), .Z(n825) );
  NOR2_X1 U917 ( .A1(n832), .A2(n825), .ZN(n829) );
  NAND2_X1 U918 ( .A1(n829), .A2(G36), .ZN(G176) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n826), .ZN(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U921 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(G188) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  NOR2_X1 U926 ( .A1(n831), .A2(n830), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  INV_X1 U928 ( .A(n832), .ZN(G319) );
  XOR2_X1 U929 ( .A(G2096), .B(KEYINPUT43), .Z(n834) );
  XNOR2_X1 U930 ( .A(G2090), .B(G2678), .ZN(n833) );
  XNOR2_X1 U931 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U932 ( .A(n835), .B(KEYINPUT42), .Z(n837) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2072), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U935 ( .A(KEYINPUT110), .B(G2100), .Z(n839) );
  XNOR2_X1 U936 ( .A(G2078), .B(G2084), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n841), .B(n840), .ZN(G227) );
  XOR2_X1 U939 ( .A(G1976), .B(G1956), .Z(n843) );
  XNOR2_X1 U940 ( .A(G1996), .B(G1961), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U942 ( .A(G1981), .B(G1971), .Z(n845) );
  XNOR2_X1 U943 ( .A(G1986), .B(G1966), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U945 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U946 ( .A(KEYINPUT111), .B(G2474), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n851) );
  XOR2_X1 U948 ( .A(G1991), .B(KEYINPUT41), .Z(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(G229) );
  NAND2_X1 U950 ( .A1(G124), .A2(n872), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n852), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U952 ( .A1(G100), .A2(n877), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n853), .B(KEYINPUT112), .ZN(n854) );
  NAND2_X1 U954 ( .A1(n855), .A2(n854), .ZN(n859) );
  NAND2_X1 U955 ( .A1(G136), .A2(n876), .ZN(n857) );
  NAND2_X1 U956 ( .A1(G112), .A2(n873), .ZN(n856) );
  NAND2_X1 U957 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U958 ( .A1(n859), .A2(n858), .ZN(G162) );
  XNOR2_X1 U959 ( .A(G160), .B(n860), .ZN(n890) );
  XNOR2_X1 U960 ( .A(KEYINPUT48), .B(KEYINPUT114), .ZN(n863) );
  XNOR2_X1 U961 ( .A(n861), .B(KEYINPUT46), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(n886) );
  NAND2_X1 U963 ( .A1(G127), .A2(n872), .ZN(n865) );
  NAND2_X1 U964 ( .A1(G115), .A2(n873), .ZN(n864) );
  NAND2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n866), .B(KEYINPUT47), .ZN(n868) );
  NAND2_X1 U967 ( .A1(G139), .A2(n876), .ZN(n867) );
  NAND2_X1 U968 ( .A1(n868), .A2(n867), .ZN(n871) );
  NAND2_X1 U969 ( .A1(G103), .A2(n877), .ZN(n869) );
  XNOR2_X1 U970 ( .A(KEYINPUT113), .B(n869), .ZN(n870) );
  NOR2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n963) );
  XNOR2_X1 U972 ( .A(G162), .B(n963), .ZN(n884) );
  NAND2_X1 U973 ( .A1(G130), .A2(n872), .ZN(n875) );
  NAND2_X1 U974 ( .A1(G118), .A2(n873), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n882) );
  NAND2_X1 U976 ( .A1(G142), .A2(n876), .ZN(n879) );
  NAND2_X1 U977 ( .A1(G106), .A2(n877), .ZN(n878) );
  NAND2_X1 U978 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U979 ( .A(KEYINPUT45), .B(n880), .Z(n881) );
  NOR2_X1 U980 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U982 ( .A(n886), .B(n885), .Z(n888) );
  XNOR2_X1 U983 ( .A(G164), .B(n974), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U985 ( .A(n890), .B(n889), .ZN(n892) );
  XNOR2_X1 U986 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U987 ( .A1(G37), .A2(n893), .ZN(G395) );
  XNOR2_X1 U988 ( .A(n998), .B(G286), .ZN(n895) );
  XNOR2_X1 U989 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U990 ( .A(G301), .B(n896), .Z(n897) );
  NOR2_X1 U991 ( .A1(G37), .A2(n897), .ZN(n898) );
  XOR2_X1 U992 ( .A(KEYINPUT115), .B(n898), .Z(G397) );
  XOR2_X1 U993 ( .A(KEYINPUT109), .B(G2427), .Z(n900) );
  XNOR2_X1 U994 ( .A(G2435), .B(G2438), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n907) );
  XOR2_X1 U996 ( .A(G2443), .B(G2430), .Z(n902) );
  XNOR2_X1 U997 ( .A(G2454), .B(G2446), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U999 ( .A(n903), .B(G2451), .Z(n905) );
  XNOR2_X1 U1000 ( .A(G1341), .B(G1348), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n908) );
  NAND2_X1 U1003 ( .A1(n908), .A2(G14), .ZN(n914) );
  NAND2_X1 U1004 ( .A1(G319), .A2(n914), .ZN(n911) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1009 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(n914), .ZN(G401) );
  XNOR2_X1 U1012 ( .A(G2067), .B(G26), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(G1996), .B(G32), .ZN(n915) );
  NOR2_X1 U1014 ( .A1(n916), .A2(n915), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(n917), .B(G27), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(G33), .B(G2072), .ZN(n918) );
  NOR2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1019 ( .A(KEYINPUT117), .B(n922), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n923), .A2(G28), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(G25), .B(G1991), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1023 ( .A(KEYINPUT53), .B(n926), .Z(n929) );
  XOR2_X1 U1024 ( .A(G34), .B(KEYINPUT54), .Z(n927) );
  XNOR2_X1 U1025 ( .A(G2084), .B(n927), .ZN(n928) );
  NAND2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(G35), .B(G2090), .ZN(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(n932), .B(KEYINPUT118), .ZN(n933) );
  NOR2_X1 U1030 ( .A1(G29), .A2(n933), .ZN(n934) );
  XNOR2_X1 U1031 ( .A(KEYINPUT55), .B(n934), .ZN(n1018) );
  XOR2_X1 U1032 ( .A(G4), .B(KEYINPUT123), .Z(n936) );
  XNOR2_X1 U1033 ( .A(G1348), .B(KEYINPUT59), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(n936), .B(n935), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(G1956), .B(G20), .ZN(n938) );
  XNOR2_X1 U1036 ( .A(G1981), .B(G6), .ZN(n937) );
  NOR2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(KEYINPUT122), .B(G1341), .ZN(n941) );
  XNOR2_X1 U1040 ( .A(G19), .B(n941), .ZN(n942) );
  NOR2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1042 ( .A(KEYINPUT60), .B(n944), .ZN(n955) );
  XOR2_X1 U1043 ( .A(G1971), .B(G22), .Z(n945) );
  XNOR2_X1 U1044 ( .A(KEYINPUT125), .B(n945), .ZN(n947) );
  XNOR2_X1 U1045 ( .A(G23), .B(G1976), .ZN(n946) );
  NOR2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1047 ( .A(KEYINPUT126), .B(n948), .Z(n950) );
  XNOR2_X1 U1048 ( .A(G1986), .B(G24), .ZN(n949) );
  NOR2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1050 ( .A(KEYINPUT58), .B(n951), .Z(n953) );
  XNOR2_X1 U1051 ( .A(G1961), .B(G5), .ZN(n952) );
  NOR2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1053 ( .A1(n955), .A2(n954), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(KEYINPUT124), .B(G1966), .ZN(n956) );
  XNOR2_X1 U1055 ( .A(G21), .B(n956), .ZN(n957) );
  NOR2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1057 ( .A(n959), .B(KEYINPUT61), .ZN(n961) );
  XNOR2_X1 U1058 ( .A(G16), .B(KEYINPUT121), .ZN(n960) );
  NAND2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1060 ( .A1(G11), .A2(n962), .ZN(n1016) );
  XOR2_X1 U1061 ( .A(G2072), .B(n963), .Z(n965) );
  XOR2_X1 U1062 ( .A(G164), .B(G2078), .Z(n964) );
  NOR2_X1 U1063 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1064 ( .A(n966), .B(KEYINPUT50), .ZN(n968) );
  NAND2_X1 U1065 ( .A1(n968), .A2(n967), .ZN(n973) );
  XOR2_X1 U1066 ( .A(G2090), .B(G162), .Z(n969) );
  NOR2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(n971), .B(KEYINPUT51), .ZN(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(G160), .B(G2084), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(n978), .B(KEYINPUT116), .ZN(n979) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(n985), .B(KEYINPUT52), .ZN(n986) );
  NAND2_X1 U1078 ( .A1(n986), .A2(G29), .ZN(n1014) );
  XNOR2_X1 U1079 ( .A(KEYINPUT56), .B(G16), .ZN(n1012) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(n989), .B(G1956), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(G1971), .A2(G303), .ZN(n990) );
  NAND2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n1005) );
  XOR2_X1 U1086 ( .A(n996), .B(G1341), .Z(n1003) );
  XNOR2_X1 U1087 ( .A(G171), .B(G1961), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(n997), .B(KEYINPUT119), .ZN(n1000) );
  XOR2_X1 U1089 ( .A(G1348), .B(n998), .Z(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(KEYINPUT120), .B(n1001), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(G1966), .B(G168), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(n1008), .B(KEYINPUT57), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1100 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1101 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1102 ( .A(n1019), .B(KEYINPUT62), .ZN(n1020) );
  XNOR2_X1 U1103 ( .A(KEYINPUT127), .B(n1020), .ZN(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

