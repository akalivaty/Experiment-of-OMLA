//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0' ..
//Module:
 module locked_c2670( 
    G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
    G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
    G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
    G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
    G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
    G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
    G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136,
    G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180,
    G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194,
    G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206,
    G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241,
    G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253,
    G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269,
    G270, G271, G272, G273, G274, G275, G276, G277, G278, G279, G452, G483,
    G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384,
    G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066,
    G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106,
    G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  , KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0);
input KEYINPUT0;
input KEYINPUT1;
input KEYINPUT2;
input KEYINPUT3;
input KEYINPUT4;
input KEYINPUT5;
input KEYINPUT6;
input KEYINPUT7;
input KEYINPUT8;
input KEYINPUT9;
input KEYINPUT10;
input KEYINPUT11;
input KEYINPUT12;
input KEYINPUT13;
input KEYINPUT14;
input KEYINPUT15;
input KEYINPUT16;
input KEYINPUT17;
input KEYINPUT18;
input KEYINPUT19;
input KEYINPUT20;
input KEYINPUT21;
input KEYINPUT22;
input KEYINPUT23;
input KEYINPUT24;
input KEYINPUT25;
input KEYINPUT26;
input KEYINPUT27;
input KEYINPUT28;
input KEYINPUT29;
input KEYINPUT30;
input KEYINPUT31;
input KEYINPUT32;
input KEYINPUT33;
input KEYINPUT34;
input KEYINPUT35;
input KEYINPUT36;
input KEYINPUT37;
input KEYINPUT38;
input KEYINPUT39;
input KEYINPUT40;
input KEYINPUT41;
input KEYINPUT42;
input KEYINPUT43;
input KEYINPUT44;
input KEYINPUT45;
input KEYINPUT46;
input KEYINPUT47;
input KEYINPUT48;
input KEYINPUT49;
input KEYINPUT50;
input KEYINPUT51;
input KEYINPUT52;
input KEYINPUT53;
input KEYINPUT54;
input KEYINPUT55;
input KEYINPUT56;
input KEYINPUT57;
input KEYINPUT58;
input KEYINPUT59;
input KEYINPUT60;
input KEYINPUT61;
input KEYINPUT62;
input KEYINPUT63;
//Header:
   input  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20,
    G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36,
    G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74,
    G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90,
    G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105,
    G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
    G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135,
    G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179,
    G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193,
    G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205,
    G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240,
    G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252,
    G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268,
    G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279, G452,
    G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348,
    G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996,
    G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105,
    G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474,
    G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n321_, new_n322_, new_n323_, new_n324_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n341_, new_n342_, new_n343_,
    new_n344_, new_n345_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n361_, new_n362_, new_n363_, new_n364_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n374_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n381_, new_n382_, new_n383_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n405_, new_n406_, new_n409_,
    new_n411_, new_n412_, new_n413_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n736_, new_n737_,
    new_n738_;
wire RLL_wire_A_0;
wire RLL_wire_A_1;
wire RLL_wire_A_2;
wire RLL_wire_A_3;
wire RLL_wire_A_4;
wire RLL_wire_A_5;
wire RLL_wire_A_6;
wire RLL_wire_A_7;
wire RLL_wire_A_8;
wire RLL_wire_A_9;
wire RLL_wire_A_10;
wire RLL_wire_A_11;
wire RLL_wire_A_12;
wire RLL_wire_A_13;
wire RLL_wire_A_14;
wire RLL_wire_A_15;
wire RLL_wire_A_16;
wire RLL_wire_A_17;
wire RLL_wire_A_18;
wire RLL_wire_A_19;
wire RLL_wire_A_20;
wire RLL_wire_A_21;
wire RLL_wire_A_22;
wire RLL_wire_A_23;
wire RLL_wire_A_24;
wire RLL_wire_A_25;
wire RLL_wire_A_26;
wire RLL_wire_A_27;
wire RLL_wire_A_28;
wire RLL_wire_A_29;
wire RLL_wire_A_30;
wire RLL_wire_A_31;
wire RLL_wire_A_32;
wire RLL_wire_A_33;
wire RLL_wire_A_34;
wire RLL_wire_A_35;
wire RLL_wire_A_36;
wire RLL_wire_A_37;
wire RLL_wire_A_38;
wire RLL_wire_A_39;
wire RLL_wire_A_40;
wire RLL_wire_A_41;
wire RLL_wire_A_42;
wire RLL_wire_A_43;
wire RLL_wire_A_44;
wire RLL_wire_A_45;
wire RLL_wire_A_46;
wire RLL_wire_A_47;
wire RLL_wire_A_48;
wire RLL_wire_A_49;
wire RLL_wire_A_50;
wire RLL_wire_A_51;
wire RLL_wire_A_52;
wire RLL_wire_A_53;
wire RLL_wire_A_54;
wire RLL_wire_A_55;
wire RLL_wire_A_56;
wire RLL_wire_A_57;
wire RLL_wire_A_58;
wire RLL_wire_A_59;
wire RLL_wire_A_60;
wire RLL_wire_A_61;
wire RLL_wire_A_62;
wire RLL_wire_A_63;

//Body:
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  INV_X1    g010(.A(G82), .ZN(RLL_wire_A_0));
  XOR2_X1 RLL_XOR_0 (.A(RLL_wire_A_0), .B(KEYINPUT0), .Z(G220) );
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(RLL_wire_A_1));
  XOR2_X1 RLL_XOR_1 (.A(RLL_wire_A_1), .B(KEYINPUT1), .Z(G223) );
  NAND3_X1  g021(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g022(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g023(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n321_));
  INV_X1    g024(.A(new_n321_), .ZN(new_n322_));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(RLL_wire_A_2));
  XNOR2_X1 RLL_XNOR_2 (.A(RLL_wire_A_2), .B(KEYINPUT2), .ZN(new_n323_) );
  INV_X1    g026(.A(new_n323_), .ZN(new_n324_));
  NOR2_X1   g027(.A1(new_n322_), .A2(new_n324_), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  AOI22_X1  g029(.A1(G567), .A2(new_n322_), .B1(new_n324_), .B2(G2106), .ZN(G319));
  INV_X1    g030(.A(G2105), .ZN(new_n328_));
  NAND3_X1  g031(.A1(new_n328_), .A2(G101), .A3(G2104), .ZN(new_n329_));
  INV_X1    g032(.A(G2104), .ZN(RLL_wire_A_3));
  XOR2_X1 RLL_XOR_3 (.A(RLL_wire_A_3), .B(KEYINPUT3), .Z(new_n330_) );
  NAND3_X1  g033(.A1(new_n330_), .A2(new_n328_), .A3(G137), .ZN(new_n331_));
  NAND3_X1  g034(.A1(G113), .A2(G2104), .A3(G2105), .ZN(new_n332_));
  NAND3_X1  g035(.A1(new_n330_), .A2(G125), .A3(G2105), .ZN(new_n333_));
  AND4_X1   g036(.A1(new_n329_), .A2(new_n331_), .A3(new_n332_), .A4(new_n333_), .ZN(G160));
  NAND3_X1  g037(.A1(new_n330_), .A2(new_n328_), .A3(G136), .ZN(new_n335_));
  NAND3_X1  g038(.A1(new_n328_), .A2(G100), .A3(G2104), .ZN(new_n336_));
  NAND3_X1  g039(.A1(new_n330_), .A2(G124), .A3(G2105), .ZN(new_n337_));
  NAND3_X1  g040(.A1(G112), .A2(G2104), .A3(G2105), .ZN(new_n338_));
  NAND4_X1  g041(.A1(new_n335_), .A2(new_n336_), .A3(new_n337_), .A4(new_n338_), .ZN(new_n339_));
  INV_X1    g042(.A(new_n339_), .ZN(G162));
  NAND3_X1  g043(.A1(new_n330_), .A2(new_n328_), .A3(G138), .ZN(RLL_wire_A_4));
  XNOR2_X1 RLL_XNOR_4 (.A(RLL_wire_A_4), .B(KEYINPUT4), .ZN(new_n341_) );
  NAND3_X1  g044(.A1(new_n328_), .A2(G102), .A3(G2104), .ZN(new_n342_));
  NAND3_X1  g045(.A1(new_n330_), .A2(G126), .A3(G2105), .ZN(new_n343_));
  NAND3_X1  g046(.A1(G114), .A2(G2104), .A3(G2105), .ZN(new_n344_));
  NAND4_X1  g047(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .A4(new_n344_), .ZN(new_n345_));
  INV_X1    g048(.A(new_n345_), .ZN(G164));
  INV_X1    g049(.A(G543), .ZN(RLL_wire_A_5));
  XOR2_X1 RLL_XOR_5 (.A(RLL_wire_A_5), .B(KEYINPUT5), .Z(new_n347_) );
  INV_X1    g050(.A(G651), .ZN(RLL_wire_A_6));
  XOR2_X1 RLL_XOR_6 (.A(RLL_wire_A_6), .B(KEYINPUT6), .Z(new_n348_) );
  NAND3_X1  g051(.A1(new_n347_), .A2(new_n348_), .A3(G88), .ZN(new_n349_));
  NAND3_X1  g052(.A1(new_n348_), .A2(G50), .A3(G543), .ZN(new_n350_));
  NAND3_X1  g053(.A1(new_n347_), .A2(G62), .A3(G651), .ZN(new_n351_));
  NAND3_X1  g054(.A1(G75), .A2(G543), .A3(G651), .ZN(new_n352_));
  NAND4_X1  g055(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .A4(new_n352_), .ZN(G303));
  INV_X1    g056(.A(G303), .ZN(G166));
  NAND3_X1  g057(.A1(new_n347_), .A2(new_n348_), .A3(G89), .ZN(new_n355_));
  NAND3_X1  g058(.A1(new_n348_), .A2(G51), .A3(G543), .ZN(new_n356_));
  NAND3_X1  g059(.A1(new_n347_), .A2(G63), .A3(G651), .ZN(new_n357_));
  NAND3_X1  g060(.A1(G76), .A2(G543), .A3(G651), .ZN(RLL_wire_A_7));
  XNOR2_X1 RLL_XNOR_7 (.A(RLL_wire_A_7), .B(KEYINPUT7), .ZN(new_n358_) );
  NAND4_X1  g061(.A1(new_n355_), .A2(new_n356_), .A3(new_n357_), .A4(new_n358_), .ZN(G286));
  INV_X1    g062(.A(G286), .ZN(G168));
  NAND3_X1  g063(.A1(new_n347_), .A2(new_n348_), .A3(G90), .ZN(new_n361_));
  NAND3_X1  g064(.A1(new_n348_), .A2(G52), .A3(G543), .ZN(new_n362_));
  NAND3_X1  g065(.A1(new_n347_), .A2(G64), .A3(G651), .ZN(new_n363_));
  NAND3_X1  g066(.A1(G77), .A2(G543), .A3(G651), .ZN(new_n364_));
  NAND4_X1  g067(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .A4(new_n364_), .ZN(G301));
  INV_X1    g068(.A(G301), .ZN(G171));
  NAND3_X1  g069(.A1(new_n347_), .A2(new_n348_), .A3(G81), .ZN(new_n367_));
  NAND3_X1  g070(.A1(new_n347_), .A2(G56), .A3(G651), .ZN(new_n368_));
  NAND3_X1  g071(.A1(G68), .A2(G543), .A3(G651), .ZN(new_n369_));
  AND3_X1   g072(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  NAND3_X1  g073(.A1(new_n348_), .A2(G43), .A3(G543), .ZN(new_n371_));
  NAND3_X1  g074(.A1(new_n370_), .A2(G860), .A3(new_n371_), .ZN(G153));
  NAND4_X1  g075(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g076(.A1(G1), .A2(G3), .ZN(RLL_wire_A_8));
  XNOR2_X1 RLL_XNOR_8 (.A(RLL_wire_A_8), .B(KEYINPUT8), .ZN(new_n374_) );
  NAND4_X1  g077(.A1(G319), .A2(G483), .A3(G661), .A4(new_n374_), .ZN(G188));
  NAND3_X1  g078(.A1(new_n347_), .A2(new_n348_), .A3(G91), .ZN(new_n376_));
  NAND3_X1  g079(.A1(new_n348_), .A2(G53), .A3(G543), .ZN(RLL_wire_A_9));
  XNOR2_X1 RLL_XNOR_9 (.A(RLL_wire_A_9), .B(KEYINPUT9), .ZN(new_n377_) );
  NAND3_X1  g080(.A1(new_n347_), .A2(G65), .A3(G651), .ZN(new_n378_));
  NAND3_X1  g081(.A1(G78), .A2(G543), .A3(G651), .ZN(new_n379_));
  NAND4_X1  g082(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .A4(new_n379_), .ZN(G299));
  OAI21_X1  g083(.A(G651), .B1(new_n347_), .B2(G74), .ZN(new_n381_));
  NAND3_X1  g084(.A1(new_n347_), .A2(new_n348_), .A3(G87), .ZN(new_n382_));
  NAND3_X1  g085(.A1(new_n348_), .A2(G49), .A3(G543), .ZN(new_n383_));
  NAND3_X1  g086(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(G288));
  NAND3_X1  g087(.A1(new_n347_), .A2(new_n348_), .A3(G86), .ZN(new_n385_));
  NAND3_X1  g088(.A1(new_n348_), .A2(G48), .A3(G543), .ZN(new_n386_));
  NAND3_X1  g089(.A1(new_n347_), .A2(G61), .A3(G651), .ZN(new_n387_));
  NAND3_X1  g090(.A1(G73), .A2(G543), .A3(G651), .ZN(new_n388_));
  NAND4_X1  g091(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .A4(new_n388_), .ZN(G305));
  NAND3_X1  g092(.A1(new_n347_), .A2(new_n348_), .A3(G85), .ZN(new_n390_));
  NAND3_X1  g093(.A1(new_n348_), .A2(G47), .A3(G543), .ZN(new_n391_));
  NAND3_X1  g094(.A1(new_n347_), .A2(G60), .A3(G651), .ZN(new_n392_));
  NAND3_X1  g095(.A1(G72), .A2(G543), .A3(G651), .ZN(new_n393_));
  NAND4_X1  g096(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .A4(new_n393_), .ZN(G290));
  NAND2_X1  g097(.A1(G301), .A2(G868), .ZN(new_n395_));
  NAND3_X1  g098(.A1(new_n347_), .A2(new_n348_), .A3(G92), .ZN(RLL_wire_A_10));
  XOR2_X1 RLL_XOR_10 (.A(RLL_wire_A_10), .B(KEYINPUT10), .Z(new_n396_) );
  NAND3_X1  g099(.A1(new_n347_), .A2(G66), .A3(G651), .ZN(new_n397_));
  NAND3_X1  g100(.A1(G79), .A2(G543), .A3(G651), .ZN(new_n398_));
  AND3_X1   g101(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  NAND3_X1  g102(.A1(new_n348_), .A2(G54), .A3(G543), .ZN(new_n400_));
  NAND2_X1  g103(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g104(.A(new_n401_), .ZN(new_n402_));
  OAI21_X1  g105(.A(new_n395_), .B1(new_n402_), .B2(G868), .ZN(G284));
  OAI21_X1  g106(.A(new_n395_), .B1(new_n402_), .B2(G868), .ZN(G321));
  INV_X1    g107(.A(G868), .ZN(new_n405_));
  NAND2_X1  g108(.A1(G299), .A2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g109(.A(new_n406_), .B1(G168), .B2(new_n405_), .ZN(G297));
  OAI21_X1  g110(.A(new_n406_), .B1(G168), .B2(new_n405_), .ZN(G280));
  INV_X1    g111(.A(G559), .ZN(new_n409_));
  OAI21_X1  g112(.A(new_n402_), .B1(new_n409_), .B2(G860), .ZN(G148));
  NAND2_X1  g113(.A1(new_n370_), .A2(new_n371_), .ZN(new_n411_));
  NAND2_X1  g114(.A1(new_n411_), .A2(new_n405_), .ZN(new_n412_));
  NOR2_X1   g115(.A1(new_n401_), .A2(G559), .ZN(new_n413_));
  OAI21_X1  g116(.A(new_n412_), .B1(new_n413_), .B2(new_n405_), .ZN(RLL_wire_A_11));
  XNOR2_X1 RLL_XNOR_11 (.A(RLL_wire_A_11), .B(KEYINPUT11), .ZN(G282) );
  OAI21_X1  g117(.A(new_n412_), .B1(new_n413_), .B2(new_n405_), .ZN(G323));
  NAND3_X1  g118(.A1(new_n330_), .A2(new_n328_), .A3(G135), .ZN(new_n416_));
  NAND3_X1  g119(.A1(new_n328_), .A2(G99), .A3(G2104), .ZN(new_n417_));
  NAND3_X1  g120(.A1(new_n330_), .A2(G123), .A3(G2105), .ZN(new_n418_));
  NAND3_X1  g121(.A1(G111), .A2(G2104), .A3(G2105), .ZN(new_n419_));
  NAND4_X1  g122(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .A4(new_n419_), .ZN(new_n420_));
  XOR2_X1   g123(.A(new_n420_), .B(G2096), .Z(new_n421_));
  NOR2_X1   g124(.A1(new_n330_), .A2(G2105), .ZN(new_n422_));
  NAND2_X1  g125(.A1(new_n328_), .A2(G2104), .ZN(new_n423_));
  NOR2_X1   g126(.A1(new_n422_), .A2(new_n423_), .ZN(RLL_wire_A_12));
  XOR2_X1 RLL_XOR_12 (.A(RLL_wire_A_12), .B(KEYINPUT12), .Z(new_n424_) );
  XNOR2_X1  g127(.A(new_n424_), .B(G2100), .ZN(RLL_wire_A_13));
  XNOR2_X1 RLL_XNOR_13 (.A(RLL_wire_A_13), .B(KEYINPUT13), .ZN(new_n425_) );
  NAND2_X1  g128(.A1(new_n421_), .A2(new_n425_), .ZN(G156));
  XNOR2_X1  g129(.A(G2435), .B(G2438), .ZN(new_n427_));
  INV_X1    g130(.A(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g131(.A(G2443), .B(G2446), .ZN(new_n429_));
  INV_X1    g132(.A(new_n429_), .ZN(RLL_wire_A_14));
  XNOR2_X1 RLL_XNOR_14 (.A(RLL_wire_A_14), .B(KEYINPUT14), .ZN(new_n430_) );
  XNOR2_X1  g133(.A(G2427), .B(G2430), .ZN(RLL_wire_A_15));
  XOR2_X1 RLL_XOR_15 (.A(RLL_wire_A_15), .B(KEYINPUT15), .Z(new_n431_) );
  INV_X1    g134(.A(new_n431_), .ZN(new_n432_));
  NAND3_X1  g135(.A1(new_n428_), .A2(new_n430_), .A3(new_n432_), .ZN(new_n433_));
  NAND3_X1  g136(.A1(new_n432_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n434_));
  NAND3_X1  g137(.A1(new_n430_), .A2(new_n427_), .A3(new_n431_), .ZN(new_n435_));
  NAND3_X1  g138(.A1(new_n428_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n436_));
  NAND4_X1  g139(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .A4(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g140(.A(G2451), .B(G2454), .ZN(RLL_wire_A_16));
  XNOR2_X1 RLL_XNOR_16 (.A(RLL_wire_A_16), .B(KEYINPUT16), .ZN(new_n438_) );
  XNOR2_X1  g141(.A(G1341), .B(G1348), .ZN(new_n439_));
  XNOR2_X1  g142(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  XOR2_X1   g143(.A(new_n437_), .B(new_n440_), .Z(new_n441_));
  NAND2_X1  g144(.A1(new_n441_), .A2(G14), .ZN(new_n442_));
  INV_X1    g145(.A(new_n442_), .ZN(G401));
  XNOR2_X1  g146(.A(G2072), .B(G2078), .ZN(new_n444_));
  INV_X1    g147(.A(new_n444_), .ZN(RLL_wire_A_17));
  XNOR2_X1 RLL_XNOR_17 (.A(RLL_wire_A_17), .B(KEYINPUT17), .ZN(new_n445_) );
  XNOR2_X1  g148(.A(G2084), .B(G2090), .ZN(new_n446_));
  INV_X1    g149(.A(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g150(.A(G2067), .B(G2678), .ZN(new_n448_));
  INV_X1    g151(.A(new_n448_), .ZN(new_n449_));
  NAND3_X1  g152(.A1(new_n445_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n450_));
  NAND3_X1  g153(.A1(new_n449_), .A2(new_n444_), .A3(new_n446_), .ZN(new_n451_));
  NAND3_X1  g154(.A1(new_n447_), .A2(new_n444_), .A3(new_n448_), .ZN(RLL_wire_A_18));
  XOR2_X1 RLL_XOR_18 (.A(RLL_wire_A_18), .B(KEYINPUT18), .Z(new_n452_) );
  NAND3_X1  g155(.A1(new_n445_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n453_));
  NAND4_X1  g156(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .A4(new_n453_), .ZN(new_n454_));
  XOR2_X1   g157(.A(G2096), .B(G2100), .Z(new_n455_));
  XNOR2_X1  g158(.A(new_n454_), .B(new_n455_), .ZN(G227));
  XNOR2_X1  g159(.A(G1961), .B(G1966), .ZN(new_n457_));
  INV_X1    g160(.A(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g161(.A(G1971), .B(G1976), .ZN(RLL_wire_A_19));
  XNOR2_X1 RLL_XNOR_19 (.A(RLL_wire_A_19), .B(KEYINPUT19), .ZN(new_n459_) );
  INV_X1    g162(.A(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g163(.A(G1956), .B(G2474), .ZN(new_n461_));
  INV_X1    g164(.A(new_n461_), .ZN(new_n462_));
  NAND3_X1  g165(.A1(new_n458_), .A2(new_n460_), .A3(new_n462_), .ZN(RLL_wire_A_20));
  XNOR2_X1 RLL_XNOR_20 (.A(RLL_wire_A_20), .B(KEYINPUT20), .ZN(new_n463_) );
  NAND3_X1  g166(.A1(new_n462_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n464_));
  NAND3_X1  g167(.A1(new_n460_), .A2(new_n457_), .A3(new_n461_), .ZN(new_n465_));
  NAND3_X1  g168(.A1(new_n458_), .A2(new_n459_), .A3(new_n461_), .ZN(new_n466_));
  NAND4_X1  g169(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .A4(new_n466_), .ZN(new_n467_));
  XOR2_X1   g170(.A(G1981), .B(G1986), .Z(RLL_wire_A_21));
  XOR2_X1 RLL_XOR_21 (.A(RLL_wire_A_21), .B(KEYINPUT21), .Z(new_n468_) );
  XNOR2_X1  g171(.A(G1991), .B(G1996), .ZN(new_n469_));
  XNOR2_X1  g172(.A(new_n468_), .B(new_n469_), .ZN(RLL_wire_A_22));
  XNOR2_X1 RLL_XNOR_22 (.A(RLL_wire_A_22), .B(KEYINPUT22), .ZN(new_n470_) );
  XNOR2_X1  g173(.A(new_n467_), .B(new_n470_), .ZN(G229));
  INV_X1    g174(.A(G19), .ZN(new_n472_));
  NOR2_X1   g175(.A1(new_n472_), .A2(G16), .ZN(new_n473_));
  AOI21_X1  g176(.A(new_n473_), .B1(new_n411_), .B2(G16), .ZN(new_n474_));
  XNOR2_X1  g177(.A(new_n474_), .B(G1341), .ZN(new_n475_));
  INV_X1    g178(.A(G4), .ZN(new_n476_));
  NOR2_X1   g179(.A1(new_n476_), .A2(G16), .ZN(new_n477_));
  AOI21_X1  g180(.A(new_n477_), .B1(new_n401_), .B2(G16), .ZN(new_n478_));
  XNOR2_X1  g181(.A(new_n478_), .B(G1348), .ZN(new_n479_));
  INV_X1    g182(.A(G20), .ZN(new_n480_));
  NOR2_X1   g183(.A1(new_n480_), .A2(G16), .ZN(RLL_wire_A_23));
  XNOR2_X1 RLL_XNOR_23 (.A(RLL_wire_A_23), .B(KEYINPUT23), .ZN(new_n481_) );
  AOI21_X1  g184(.A(new_n481_), .B1(G299), .B2(G16), .ZN(new_n482_));
  XNOR2_X1  g185(.A(new_n482_), .B(G1956), .ZN(new_n483_));
  NAND3_X1  g186(.A1(new_n475_), .A2(new_n479_), .A3(new_n483_), .ZN(new_n484_));
  MUX2_X1   g187(.A(G5), .B(G301), .S(G16), .Z(new_n485_));
  XNOR2_X1  g188(.A(new_n485_), .B(G1961), .ZN(new_n486_));
  INV_X1    g189(.A(G21), .ZN(new_n487_));
  NOR2_X1   g190(.A1(new_n487_), .A2(G16), .ZN(new_n488_));
  AOI21_X1  g191(.A(new_n488_), .B1(G286), .B2(G16), .ZN(new_n489_));
  XOR2_X1   g192(.A(new_n489_), .B(G1966), .Z(new_n490_));
  NOR3_X1   g193(.A1(new_n484_), .A2(new_n486_), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g194(.A(G34), .ZN(RLL_wire_A_24));
  XOR2_X1 RLL_XOR_24 (.A(RLL_wire_A_24), .B(KEYINPUT24), .Z(new_n492_) );
  NOR2_X1   g195(.A1(new_n492_), .A2(G29), .ZN(new_n493_));
  NAND4_X1  g196(.A1(new_n331_), .A2(new_n329_), .A3(new_n333_), .A4(new_n332_), .ZN(new_n494_));
  AOI21_X1  g197(.A(new_n493_), .B1(new_n494_), .B2(G29), .ZN(new_n495_));
  XNOR2_X1  g198(.A(new_n495_), .B(G2084), .ZN(new_n496_));
  INV_X1    g199(.A(G33), .ZN(new_n497_));
  NOR2_X1   g200(.A1(new_n497_), .A2(G29), .ZN(new_n498_));
  NAND3_X1  g201(.A1(new_n330_), .A2(new_n328_), .A3(G139), .ZN(new_n499_));
  NAND3_X1  g202(.A1(new_n328_), .A2(G103), .A3(G2104), .ZN(RLL_wire_A_25));
  XOR2_X1 RLL_XOR_25 (.A(RLL_wire_A_25), .B(KEYINPUT25), .Z(new_n500_) );
  NAND3_X1  g203(.A1(new_n330_), .A2(G127), .A3(G2105), .ZN(new_n501_));
  NAND3_X1  g204(.A1(G115), .A2(G2104), .A3(G2105), .ZN(new_n502_));
  NAND4_X1  g205(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .A4(new_n502_), .ZN(new_n503_));
  AOI21_X1  g206(.A(new_n498_), .B1(new_n503_), .B2(G29), .ZN(new_n504_));
  XNOR2_X1  g207(.A(new_n504_), .B(G2072), .ZN(new_n505_));
  INV_X1    g208(.A(G32), .ZN(new_n506_));
  NOR2_X1   g209(.A1(new_n506_), .A2(G29), .ZN(new_n507_));
  NAND3_X1  g210(.A1(new_n330_), .A2(new_n328_), .A3(G141), .ZN(new_n508_));
  NAND3_X1  g211(.A1(new_n328_), .A2(G105), .A3(G2104), .ZN(new_n509_));
  NAND3_X1  g212(.A1(new_n330_), .A2(G129), .A3(G2105), .ZN(new_n510_));
  NAND3_X1  g213(.A1(G117), .A2(G2104), .A3(G2105), .ZN(RLL_wire_A_26));
  XOR2_X1 RLL_XOR_26 (.A(RLL_wire_A_26), .B(KEYINPUT26), .Z(new_n511_) );
  NAND4_X1  g214(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .A4(new_n511_), .ZN(new_n512_));
  AOI21_X1  g215(.A(new_n507_), .B1(new_n512_), .B2(G29), .ZN(new_n513_));
  XNOR2_X1  g216(.A(new_n513_), .B(G1996), .ZN(RLL_wire_A_27));
  XOR2_X1 RLL_XOR_27 (.A(RLL_wire_A_27), .B(KEYINPUT27), .Z(new_n514_) );
  INV_X1    g217(.A(G26), .ZN(new_n515_));
  NOR2_X1   g218(.A1(new_n515_), .A2(G29), .ZN(RLL_wire_A_28));
  XNOR2_X1 RLL_XNOR_28 (.A(RLL_wire_A_28), .B(KEYINPUT28), .ZN(new_n516_) );
  NAND3_X1  g219(.A1(new_n330_), .A2(new_n328_), .A3(G140), .ZN(new_n517_));
  NAND3_X1  g220(.A1(new_n328_), .A2(G104), .A3(G2104), .ZN(new_n518_));
  NAND3_X1  g221(.A1(new_n330_), .A2(G128), .A3(G2105), .ZN(new_n519_));
  NAND3_X1  g222(.A1(G116), .A2(G2104), .A3(G2105), .ZN(new_n520_));
  NAND4_X1  g223(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .A4(new_n520_), .ZN(new_n521_));
  AOI21_X1  g224(.A(new_n516_), .B1(new_n521_), .B2(G29), .ZN(new_n522_));
  XNOR2_X1  g225(.A(new_n522_), .B(G2067), .ZN(new_n523_));
  NAND4_X1  g226(.A1(new_n496_), .A2(new_n505_), .A3(new_n514_), .A4(new_n523_), .ZN(new_n524_));
  MUX2_X1   g227(.A(G35), .B(new_n339_), .S(G29), .Z(RLL_wire_A_29));
  XNOR2_X1 RLL_XNOR_29 (.A(RLL_wire_A_29), .B(KEYINPUT29), .ZN(new_n525_) );
  XNOR2_X1  g228(.A(new_n525_), .B(G2090), .ZN(new_n526_));
  MUX2_X1   g229(.A(G27), .B(new_n345_), .S(G29), .Z(new_n527_));
  XNOR2_X1  g230(.A(new_n527_), .B(G2078), .ZN(new_n528_));
  INV_X1    g231(.A(G28), .ZN(RLL_wire_A_30));
  XOR2_X1 RLL_XOR_30 (.A(RLL_wire_A_30), .B(KEYINPUT30), .Z(new_n529_) );
  NOR2_X1   g232(.A1(new_n529_), .A2(G29), .ZN(new_n530_));
  AOI21_X1  g233(.A(new_n530_), .B1(new_n420_), .B2(G29), .ZN(new_n531_));
  NOR4_X1   g234(.A1(new_n524_), .A2(new_n526_), .A3(new_n528_), .A4(new_n531_), .ZN(new_n532_));
  NAND2_X1  g235(.A1(new_n405_), .A2(G11), .ZN(new_n533_));
  NAND2_X1  g236(.A1(G11), .A2(G868), .ZN(new_n534_));
  NAND2_X1  g237(.A1(new_n533_), .A2(new_n534_), .ZN(RLL_wire_A_31));
  XNOR2_X1 RLL_XNOR_31 (.A(RLL_wire_A_31), .B(KEYINPUT31), .ZN(new_n535_) );
  INV_X1    g238(.A(G6), .ZN(new_n536_));
  NOR2_X1   g239(.A1(new_n536_), .A2(G16), .ZN(new_n537_));
  AOI21_X1  g240(.A(new_n537_), .B1(G305), .B2(G16), .ZN(RLL_wire_A_32));
  XNOR2_X1 RLL_XNOR_32 (.A(RLL_wire_A_32), .B(KEYINPUT32), .ZN(new_n538_) );
  XNOR2_X1  g241(.A(new_n538_), .B(G1981), .ZN(new_n539_));
  INV_X1    g242(.A(G22), .ZN(new_n540_));
  NOR2_X1   g243(.A1(new_n540_), .A2(G16), .ZN(new_n541_));
  AOI21_X1  g244(.A(new_n541_), .B1(G303), .B2(G16), .ZN(new_n542_));
  XNOR2_X1  g245(.A(new_n542_), .B(G1971), .ZN(new_n543_));
  INV_X1    g246(.A(G23), .ZN(new_n544_));
  NOR2_X1   g247(.A1(new_n544_), .A2(G16), .ZN(new_n545_));
  AOI21_X1  g248(.A(new_n545_), .B1(G288), .B2(G16), .ZN(new_n546_));
  XNOR2_X1  g249(.A(new_n546_), .B(G1976), .ZN(RLL_wire_A_33));
  XOR2_X1 RLL_XOR_33 (.A(RLL_wire_A_33), .B(KEYINPUT33), .Z(new_n547_) );
  NAND3_X1  g250(.A1(new_n539_), .A2(new_n543_), .A3(new_n547_), .ZN(RLL_wire_A_34));
  XNOR2_X1 RLL_XNOR_34 (.A(RLL_wire_A_34), .B(KEYINPUT34), .ZN(new_n548_) );
  MUX2_X1   g251(.A(G24), .B(G290), .S(G16), .Z(new_n549_));
  XNOR2_X1  g252(.A(new_n549_), .B(G1986), .ZN(new_n550_));
  INV_X1    g253(.A(G25), .ZN(new_n551_));
  NOR2_X1   g254(.A1(new_n551_), .A2(G29), .ZN(new_n552_));
  NAND3_X1  g255(.A1(new_n330_), .A2(new_n328_), .A3(G131), .ZN(new_n553_));
  NAND3_X1  g256(.A1(new_n328_), .A2(G95), .A3(G2104), .ZN(new_n554_));
  NAND3_X1  g257(.A1(new_n330_), .A2(G119), .A3(G2105), .ZN(new_n555_));
  NAND3_X1  g258(.A1(G107), .A2(G2104), .A3(G2105), .ZN(new_n556_));
  NAND4_X1  g259(.A1(new_n553_), .A2(new_n554_), .A3(new_n555_), .A4(new_n556_), .ZN(new_n557_));
  AOI21_X1  g260(.A(new_n552_), .B1(new_n557_), .B2(G29), .ZN(new_n558_));
  INV_X1    g261(.A(G1991), .ZN(RLL_wire_A_35));
  XNOR2_X1 RLL_XNOR_35 (.A(RLL_wire_A_35), .B(KEYINPUT35), .ZN(new_n559_) );
  XNOR2_X1  g262(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  NOR3_X1   g263(.A1(new_n548_), .A2(new_n550_), .A3(new_n560_), .ZN(RLL_wire_A_36));
  XOR2_X1 RLL_XOR_36 (.A(RLL_wire_A_36), .B(KEYINPUT36), .Z(new_n561_) );
  NAND4_X1  g264(.A1(new_n491_), .A2(new_n532_), .A3(new_n535_), .A4(new_n561_), .ZN(G150));
  INV_X1    g265(.A(G150), .ZN(G311));
  NAND3_X1  g266(.A1(new_n347_), .A2(new_n348_), .A3(G93), .ZN(new_n564_));
  NAND3_X1  g267(.A1(new_n348_), .A2(G55), .A3(G543), .ZN(new_n565_));
  NAND3_X1  g268(.A1(new_n347_), .A2(G67), .A3(G651), .ZN(new_n566_));
  NAND3_X1  g269(.A1(G80), .A2(G543), .A3(G651), .ZN(new_n567_));
  NAND4_X1  g270(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .A4(new_n567_), .ZN(new_n568_));
  NAND2_X1  g271(.A1(new_n568_), .A2(G860), .ZN(RLL_wire_A_37));
  XOR2_X1 RLL_XOR_37 (.A(RLL_wire_A_37), .B(KEYINPUT37), .Z(new_n569_) );
  XNOR2_X1  g272(.A(new_n411_), .B(new_n401_), .ZN(new_n570_));
  XNOR2_X1  g273(.A(new_n570_), .B(new_n413_), .ZN(RLL_wire_A_38));
  XNOR2_X1 RLL_XNOR_38 (.A(RLL_wire_A_38), .B(KEYINPUT38), .ZN(new_n571_) );
  XNOR2_X1  g274(.A(new_n571_), .B(new_n568_), .ZN(RLL_wire_A_39));
  XNOR2_X1 RLL_XNOR_39 (.A(RLL_wire_A_39), .B(KEYINPUT39), .ZN(new_n572_) );
  OAI21_X1  g275(.A(new_n569_), .B1(new_n572_), .B2(G860), .ZN(G145));
  XNOR2_X1  g276(.A(new_n512_), .B(new_n521_), .ZN(new_n574_));
  INV_X1    g277(.A(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g278(.A(new_n345_), .B(new_n503_), .ZN(new_n576_));
  INV_X1    g279(.A(new_n576_), .ZN(new_n577_));
  NAND3_X1  g280(.A1(new_n330_), .A2(new_n328_), .A3(G142), .ZN(new_n578_));
  NAND3_X1  g281(.A1(new_n328_), .A2(G106), .A3(G2104), .ZN(new_n579_));
  NAND3_X1  g282(.A1(new_n330_), .A2(G130), .A3(G2105), .ZN(new_n580_));
  NAND3_X1  g283(.A1(G118), .A2(G2104), .A3(G2105), .ZN(new_n581_));
  NAND4_X1  g284(.A1(new_n578_), .A2(new_n579_), .A3(new_n580_), .A4(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g285(.A(new_n557_), .B(new_n582_), .ZN(new_n583_));
  INV_X1    g286(.A(new_n583_), .ZN(new_n584_));
  NAND3_X1  g287(.A1(new_n575_), .A2(new_n577_), .A3(new_n584_), .ZN(new_n585_));
  NAND3_X1  g288(.A1(new_n584_), .A2(new_n574_), .A3(new_n576_), .ZN(new_n586_));
  NAND3_X1  g289(.A1(new_n577_), .A2(new_n574_), .A3(new_n583_), .ZN(new_n587_));
  NAND3_X1  g290(.A1(new_n575_), .A2(new_n576_), .A3(new_n583_), .ZN(new_n588_));
  NAND4_X1  g291(.A1(new_n585_), .A2(new_n586_), .A3(new_n587_), .A4(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g292(.A(G160), .B(new_n339_), .ZN(new_n590_));
  XOR2_X1   g293(.A(new_n420_), .B(new_n424_), .Z(new_n591_));
  XNOR2_X1  g294(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g295(.A(new_n589_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g296(.A(G37), .ZN(new_n594_));
  NAND2_X1  g297(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g298(.A(new_n595_), .ZN(RLL_wire_A_40));
  XOR2_X1 RLL_XOR_40 (.A(RLL_wire_A_40), .B(KEYINPUT40), .Z(G395) );
  NAND2_X1  g299(.A1(new_n568_), .A2(new_n405_), .ZN(new_n597_));
  XNOR2_X1  g300(.A(new_n411_), .B(new_n568_), .ZN(new_n598_));
  INV_X1    g301(.A(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g302(.A(new_n401_), .B(G299), .ZN(new_n600_));
  INV_X1    g303(.A(new_n600_), .ZN(RLL_wire_A_41));
  XNOR2_X1 RLL_XNOR_41 (.A(RLL_wire_A_41), .B(KEYINPUT41), .ZN(new_n601_) );
  INV_X1    g304(.A(new_n413_), .ZN(new_n602_));
  NAND3_X1  g305(.A1(new_n599_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  NAND3_X1  g306(.A1(new_n601_), .A2(new_n413_), .A3(new_n598_), .ZN(new_n604_));
  NAND3_X1  g307(.A1(new_n599_), .A2(new_n413_), .A3(new_n600_), .ZN(new_n605_));
  NAND3_X1  g308(.A1(new_n598_), .A2(new_n600_), .A3(new_n602_), .ZN(new_n606_));
  NAND4_X1  g309(.A1(new_n603_), .A2(new_n604_), .A3(new_n605_), .A4(new_n606_), .ZN(RLL_wire_A_42));
  XNOR2_X1 RLL_XNOR_42 (.A(RLL_wire_A_42), .B(KEYINPUT42), .ZN(new_n607_) );
  XOR2_X1   g310(.A(G305), .B(G290), .Z(new_n608_));
  XOR2_X1   g311(.A(G303), .B(G288), .Z(new_n609_));
  XNOR2_X1  g312(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XOR2_X1   g313(.A(new_n607_), .B(new_n610_), .Z(new_n611_));
  OAI21_X1  g314(.A(new_n597_), .B1(new_n611_), .B2(new_n405_), .ZN(G295));
  OAI21_X1  g315(.A(new_n597_), .B1(new_n611_), .B2(new_n405_), .ZN(G331));
  XNOR2_X1  g316(.A(G286), .B(G301), .ZN(new_n614_));
  INV_X1    g317(.A(new_n614_), .ZN(new_n615_));
  NAND3_X1  g318(.A1(new_n599_), .A2(new_n601_), .A3(new_n615_), .ZN(new_n616_));
  NAND3_X1  g319(.A1(new_n599_), .A2(new_n600_), .A3(new_n614_), .ZN(new_n617_));
  NAND3_X1  g320(.A1(new_n601_), .A2(new_n598_), .A3(new_n614_), .ZN(new_n618_));
  NAND3_X1  g321(.A1(new_n598_), .A2(new_n600_), .A3(new_n615_), .ZN(new_n619_));
  NAND4_X1  g322(.A1(new_n616_), .A2(new_n617_), .A3(new_n618_), .A4(new_n619_), .ZN(new_n620_));
  OR2_X1    g323(.A1(new_n620_), .A2(new_n610_), .ZN(new_n621_));
  NAND2_X1  g324(.A1(new_n620_), .A2(new_n610_), .ZN(new_n622_));
  NAND3_X1  g325(.A1(new_n621_), .A2(new_n594_), .A3(new_n622_), .ZN(RLL_wire_A_43));
  XNOR2_X1 RLL_XNOR_43 (.A(RLL_wire_A_43), .B(KEYINPUT43), .ZN(new_n623_) );
  INV_X1    g326(.A(new_n623_), .ZN(RLL_wire_A_44));
  XNOR2_X1 RLL_XNOR_44 (.A(RLL_wire_A_44), .B(KEYINPUT44), .ZN(G397) );
  INV_X1    g327(.A(G1384), .ZN(new_n625_));
  AND2_X1   g328(.A1(new_n345_), .A2(new_n625_), .ZN(RLL_wire_A_45));
  XOR2_X1 RLL_XOR_45 (.A(RLL_wire_A_45), .B(KEYINPUT45), .Z(new_n626_) );
  INV_X1    g329(.A(G40), .ZN(new_n627_));
  NOR3_X1   g330(.A1(new_n626_), .A2(new_n627_), .A3(new_n494_), .ZN(new_n628_));
  NAND4_X1  g331(.A1(G160), .A2(G40), .A3(new_n625_), .A4(new_n345_), .ZN(new_n629_));
  NAND3_X1  g332(.A1(new_n628_), .A2(new_n521_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g333(.A(G2067), .ZN(new_n631_));
  NAND3_X1  g334(.A1(new_n628_), .A2(new_n631_), .A3(new_n629_), .ZN(new_n632_));
  XNOR2_X1  g335(.A(new_n630_), .B(new_n632_), .ZN(new_n633_));
  NAND3_X1  g336(.A1(new_n628_), .A2(new_n512_), .A3(new_n629_), .ZN(new_n634_));
  INV_X1    g337(.A(G1996), .ZN(new_n635_));
  NAND3_X1  g338(.A1(new_n628_), .A2(new_n635_), .A3(new_n629_), .ZN(new_n636_));
  INV_X1    g339(.A(new_n636_), .ZN(RLL_wire_A_46));
  XOR2_X1 RLL_XOR_46 (.A(RLL_wire_A_46), .B(KEYINPUT46), .Z(new_n637_) );
  NAND3_X1  g340(.A1(new_n633_), .A2(new_n634_), .A3(new_n637_), .ZN(RLL_wire_A_47));
  XNOR2_X1 RLL_XNOR_47 (.A(RLL_wire_A_47), .B(KEYINPUT47), .ZN(new_n638_) );
  NAND3_X1  g341(.A1(new_n628_), .A2(new_n557_), .A3(new_n629_), .ZN(new_n639_));
  NAND3_X1  g342(.A1(new_n628_), .A2(new_n559_), .A3(new_n629_), .ZN(new_n640_));
  XNOR2_X1  g343(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g344(.A(new_n634_), .B(new_n636_), .ZN(new_n642_));
  INV_X1    g345(.A(G1986), .ZN(new_n643_));
  NAND3_X1  g346(.A1(new_n628_), .A2(G290), .A3(new_n629_), .ZN(new_n644_));
  AND4_X1   g347(.A1(new_n643_), .A2(new_n644_), .A3(new_n628_), .A4(new_n629_), .ZN(RLL_wire_A_48));
  XOR2_X1 RLL_XOR_48 (.A(RLL_wire_A_48), .B(KEYINPUT48), .Z(new_n645_) );
  NAND4_X1  g348(.A1(new_n633_), .A2(new_n641_), .A3(new_n642_), .A4(new_n645_), .ZN(new_n646_));
  INV_X1    g349(.A(new_n640_), .ZN(new_n647_));
  NAND4_X1  g350(.A1(new_n633_), .A2(new_n642_), .A3(new_n639_), .A4(new_n647_), .ZN(new_n648_));
  NAND4_X1  g351(.A1(new_n630_), .A2(new_n631_), .A3(new_n628_), .A4(new_n629_), .ZN(new_n649_));
  AND4_X1   g352(.A1(new_n638_), .A2(new_n646_), .A3(new_n648_), .A4(new_n649_), .ZN(new_n650_));
  INV_X1    g353(.A(G1981), .ZN(RLL_wire_A_49));
  XNOR2_X1 RLL_XNOR_49 (.A(RLL_wire_A_49), .B(KEYINPUT49), .ZN(new_n651_) );
  AND4_X1   g354(.A1(G8), .A2(new_n629_), .A3(new_n651_), .A4(G305), .ZN(new_n652_));
  OAI211_X1 g355(.A(new_n629_), .B(G8), .C1(new_n651_), .C2(G305), .ZN(new_n653_));
  NOR2_X1   g356(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g357(.A1(new_n494_), .A2(new_n627_), .ZN(new_n655_));
  AOI21_X1  g358(.A(G1966), .B1(new_n626_), .B2(new_n655_), .ZN(new_n656_));
  AND2_X1   g359(.A1(new_n333_), .A2(new_n332_), .ZN(new_n657_));
  NAND4_X1  g360(.A1(new_n657_), .A2(G40), .A3(new_n329_), .A4(new_n331_), .ZN(new_n658_));
  NAND2_X1  g361(.A1(new_n345_), .A2(new_n625_), .ZN(RLL_wire_A_50));
  XNOR2_X1 RLL_XNOR_50 (.A(RLL_wire_A_50), .B(KEYINPUT50), .ZN(new_n659_) );
  NOR3_X1   g362(.A1(new_n658_), .A2(new_n659_), .A3(G2084), .ZN(new_n660_));
  OAI21_X1  g363(.A(G8), .B1(new_n656_), .B2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g364(.A1(G286), .A2(G8), .ZN(new_n662_));
  NAND2_X1  g365(.A1(new_n661_), .A2(new_n662_), .ZN(RLL_wire_A_51));
  XNOR2_X1 RLL_XNOR_51 (.A(RLL_wire_A_51), .B(KEYINPUT51), .ZN(new_n663_) );
  INV_X1    g366(.A(new_n662_), .ZN(new_n664_));
  OAI211_X1 g367(.A(G8), .B(new_n664_), .C1(new_n656_), .C2(new_n660_), .ZN(new_n665_));
  AOI21_X1  g368(.A(new_n654_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g369(.A(G1976), .ZN(new_n667_));
  AND4_X1   g370(.A1(G8), .A2(new_n629_), .A3(new_n667_), .A4(G288), .ZN(new_n668_));
  OAI211_X1 g371(.A(new_n629_), .B(G8), .C1(new_n667_), .C2(G288), .ZN(RLL_wire_A_52));
  XOR2_X1 RLL_XOR_52 (.A(RLL_wire_A_52), .B(KEYINPUT52), .Z(new_n669_) );
  NOR2_X1   g372(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g373(.A(new_n670_), .ZN(new_n671_));
  INV_X1    g374(.A(G2078), .ZN(new_n672_));
  NAND3_X1  g375(.A1(new_n626_), .A2(new_n672_), .A3(new_n655_), .ZN(RLL_wire_A_53));
  XNOR2_X1 RLL_XNOR_53 (.A(RLL_wire_A_53), .B(KEYINPUT53), .ZN(new_n673_) );
  INV_X1    g376(.A(G1961), .ZN(new_n674_));
  OAI21_X1  g377(.A(new_n674_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n675_));
  NAND2_X1  g378(.A1(new_n673_), .A2(new_n675_), .ZN(RLL_wire_A_54));
  XOR2_X1 RLL_XOR_54 (.A(RLL_wire_A_54), .B(KEYINPUT54), .Z(new_n676_) );
  XNOR2_X1  g379(.A(new_n676_), .B(G301), .ZN(new_n677_));
  AOI21_X1  g380(.A(G1971), .B1(new_n626_), .B2(new_n655_), .ZN(new_n678_));
  NOR3_X1   g381(.A1(new_n658_), .A2(new_n659_), .A3(G2090), .ZN(new_n679_));
  OAI21_X1  g382(.A(G8), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g383(.A1(G303), .A2(G8), .ZN(RLL_wire_A_55));
  XOR2_X1 RLL_XOR_55 (.A(RLL_wire_A_55), .B(KEYINPUT55), .Z(new_n681_) );
  NAND2_X1  g384(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g385(.A(new_n681_), .ZN(new_n683_));
  OAI211_X1 g386(.A(G8), .B(new_n683_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n684_));
  NAND2_X1  g387(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  NAND4_X1  g388(.A1(new_n666_), .A2(new_n671_), .A3(new_n677_), .A4(new_n685_), .ZN(new_n686_));
  INV_X1    g389(.A(G1348), .ZN(new_n687_));
  OAI21_X1  g390(.A(new_n687_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n688_));
  NAND4_X1  g391(.A1(new_n655_), .A2(new_n625_), .A3(new_n631_), .A4(new_n345_), .ZN(new_n689_));
  AOI21_X1  g392(.A(new_n401_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g393(.A(G2072), .ZN(RLL_wire_A_56));
  XOR2_X1 RLL_XOR_56 (.A(RLL_wire_A_56), .B(KEYINPUT56), .Z(new_n691_) );
  NAND3_X1  g394(.A1(new_n626_), .A2(new_n691_), .A3(new_n655_), .ZN(new_n692_));
  INV_X1    g395(.A(G1956), .ZN(new_n693_));
  OAI21_X1  g396(.A(new_n693_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n694_));
  INV_X1    g397(.A(G299), .ZN(RLL_wire_A_57));
  XOR2_X1 RLL_XOR_57 (.A(RLL_wire_A_57), .B(KEYINPUT57), .Z(new_n695_) );
  AND3_X1   g398(.A1(new_n692_), .A2(new_n694_), .A3(new_n695_), .ZN(new_n696_));
  AOI21_X1  g399(.A(new_n695_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n697_));
  OAI21_X1  g400(.A(new_n690_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g401(.A1(new_n692_), .A2(new_n694_), .ZN(new_n699_));
  NAND2_X1  g402(.A1(new_n699_), .A2(new_n695_), .ZN(new_n700_));
  INV_X1    g403(.A(G1341), .ZN(RLL_wire_A_58));
  XNOR2_X1 RLL_XNOR_58 (.A(RLL_wire_A_58), .B(KEYINPUT58), .ZN(new_n701_) );
  NAND2_X1  g404(.A1(new_n629_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g405(.A1(new_n626_), .A2(new_n635_), .A3(new_n655_), .ZN(new_n703_));
  AOI21_X1  g406(.A(new_n411_), .B1(new_n702_), .B2(new_n703_), .ZN(RLL_wire_A_59));
  XOR2_X1 RLL_XOR_59 (.A(RLL_wire_A_59), .B(KEYINPUT59), .Z(new_n704_) );
  AND3_X1   g407(.A1(new_n688_), .A2(new_n689_), .A3(new_n402_), .ZN(RLL_wire_A_60));
  XNOR2_X1 RLL_XNOR_60 (.A(RLL_wire_A_60), .B(KEYINPUT60), .ZN(new_n705_) );
  AOI21_X1  g408(.A(new_n402_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n706_));
  OAI21_X1  g409(.A(new_n704_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g410(.A1(new_n696_), .A2(new_n697_), .ZN(RLL_wire_A_61));
  XOR2_X1 RLL_XOR_61 (.A(RLL_wire_A_61), .B(KEYINPUT61), .Z(new_n708_) );
  OAI211_X1 g411(.A(new_n698_), .B(new_n700_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n709_));
  INV_X1    g412(.A(new_n709_), .ZN(new_n710_));
  NOR2_X1   g413(.A1(new_n686_), .A2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g414(.A(G301), .B1(new_n673_), .B2(new_n675_), .ZN(new_n712_));
  OAI21_X1  g415(.A(new_n712_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n713_));
  NOR2_X1   g416(.A1(new_n713_), .A2(new_n654_), .ZN(new_n714_));
  NAND2_X1  g417(.A1(new_n663_), .A2(new_n665_), .ZN(RLL_wire_A_62));
  XOR2_X1 RLL_XOR_62 (.A(RLL_wire_A_62), .B(KEYINPUT62), .Z(new_n715_) );
  NAND3_X1  g418(.A1(new_n714_), .A2(new_n685_), .A3(new_n715_), .ZN(new_n716_));
  OAI211_X1 g419(.A(G8), .B(new_n662_), .C1(new_n656_), .C2(new_n660_), .ZN(new_n717_));
  NOR2_X1   g420(.A1(new_n670_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g421(.A(new_n654_), .ZN(new_n719_));
  NAND3_X1  g422(.A1(new_n685_), .A2(new_n718_), .A3(new_n719_), .ZN(RLL_wire_A_63));
  XOR2_X1 RLL_XOR_63 (.A(RLL_wire_A_63), .B(KEYINPUT63), .Z(new_n720_) );
  INV_X1    g423(.A(G8), .ZN(new_n721_));
  INV_X1    g424(.A(new_n629_), .ZN(new_n722_));
  OR4_X1    g425(.A1(new_n721_), .A2(new_n722_), .A3(G1981), .A4(G305), .ZN(new_n723_));
  NOR2_X1   g426(.A1(new_n680_), .A2(new_n683_), .ZN(new_n724_));
  NAND3_X1  g427(.A1(new_n719_), .A2(new_n671_), .A3(new_n724_), .ZN(new_n725_));
  NAND4_X1  g428(.A1(new_n716_), .A2(new_n720_), .A3(new_n723_), .A4(new_n725_), .ZN(new_n726_));
  AND2_X1   g429(.A1(new_n629_), .A2(G288), .ZN(new_n727_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n667_), .ZN(new_n728_));
  NOR4_X1   g431(.A1(new_n654_), .A2(new_n721_), .A3(new_n727_), .A4(new_n728_), .ZN(new_n729_));
  NOR3_X1   g432(.A1(new_n711_), .A2(new_n726_), .A3(new_n729_), .ZN(new_n730_));
  NAND3_X1  g433(.A1(new_n628_), .A2(new_n643_), .A3(new_n629_), .ZN(new_n731_));
  XNOR2_X1  g434(.A(new_n644_), .B(new_n731_), .ZN(new_n732_));
  NAND4_X1  g435(.A1(new_n633_), .A2(new_n641_), .A3(new_n642_), .A4(new_n732_), .ZN(new_n733_));
  OAI21_X1  g436(.A(new_n650_), .B1(new_n730_), .B2(new_n733_), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g437(.A(G227), .B1(new_n593_), .B2(new_n594_), .ZN(new_n736_));
  OR2_X1    g438(.A1(G401), .A2(G229), .ZN(new_n737_));
  INV_X1    g439(.A(new_n737_), .ZN(new_n738_));
  NAND4_X1  g440(.A1(new_n736_), .A2(new_n623_), .A3(G319), .A4(new_n738_), .ZN(G225));
  INV_X1    g441(.A(G225), .ZN(G308));

endmodule
