//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n815, new_n816, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n203), .B1(new_n205), .B2(KEYINPUT26), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(KEYINPUT26), .B2(new_n205), .ZN(new_n207));
  XOR2_X1   g006(.A(KEYINPUT27), .B(G183gat), .Z(new_n208));
  OAI21_X1  g007(.A(KEYINPUT28), .B1(new_n208), .B2(G190gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT68), .ZN(new_n211));
  INV_X1    g010(.A(G183gat), .ZN(new_n212));
  OR3_X1    g011(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT27), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT27), .B1(new_n211), .B2(new_n212), .ZN(new_n214));
  NOR2_X1   g013(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n207), .A2(new_n209), .A3(new_n210), .A4(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G226gat), .ZN(new_n218));
  INV_X1    g017(.A(G233gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G190gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n212), .A2(new_n221), .A3(KEYINPUT64), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(G183gat), .B2(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  AND3_X1   g024(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AND3_X1   g027(.A1(new_n225), .A2(new_n228), .A3(KEYINPUT65), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT65), .B1(new_n225), .B2(new_n228), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n202), .B1(new_n205), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT67), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT66), .B(KEYINPUT23), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n234), .B1(new_n235), .B2(new_n204), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n232), .A2(KEYINPUT66), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n232), .A2(KEYINPUT66), .ZN(new_n238));
  OAI211_X1 g037(.A(KEYINPUT67), .B(new_n205), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n233), .B1(new_n236), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT25), .B1(new_n231), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT25), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n212), .A2(new_n221), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n242), .B1(new_n228), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n217), .B(new_n220), .C1(new_n241), .C2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G197gat), .B(G204gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT22), .ZN(new_n249));
  INV_X1    g048(.A(G211gat), .ZN(new_n250));
  INV_X1    g049(.A(G218gat), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G211gat), .B(G218gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n217), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n236), .A2(new_n239), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n222), .A2(new_n224), .ZN(new_n259));
  INV_X1    g058(.A(new_n227), .ZN(new_n260));
  NAND3_X1  g059(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n258), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n233), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n225), .A2(new_n228), .A3(KEYINPUT65), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n257), .A2(new_n263), .A3(new_n264), .A4(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(new_n242), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n256), .B1(new_n267), .B2(new_n245), .ZN(new_n268));
  INV_X1    g067(.A(new_n220), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT29), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n247), .B(new_n255), .C1(new_n268), .C2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT74), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n266), .A2(new_n242), .B1(new_n240), .B2(new_n244), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n270), .B(new_n269), .C1(new_n275), .C2(new_n256), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n276), .A2(KEYINPUT74), .A3(new_n255), .A4(new_n247), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n247), .B1(new_n268), .B2(new_n271), .ZN(new_n279));
  INV_X1    g078(.A(new_n254), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n253), .B(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT75), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n279), .A2(KEYINPUT75), .A3(new_n281), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n278), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G8gat), .B(G36gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(G92gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT76), .B(G64gat), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n288), .B(new_n289), .Z(new_n290));
  NAND2_X1  g089(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n290), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n278), .A2(new_n292), .A3(new_n284), .A4(new_n285), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(KEYINPUT30), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n286), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT30), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(new_n296), .A3(new_n292), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT2), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT77), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT77), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT2), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G141gat), .B(G148gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n302), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT78), .B(G155gat), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n303), .B1(new_n310), .B2(G162gat), .ZN(new_n311));
  INV_X1    g110(.A(G148gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G141gat), .ZN(new_n313));
  INV_X1    g112(.A(G141gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G148gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n316), .B1(new_n301), .B2(new_n300), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n309), .B1(new_n311), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT79), .ZN(new_n319));
  XNOR2_X1  g118(.A(G127gat), .B(G134gat), .ZN(new_n320));
  INV_X1    g119(.A(G113gat), .ZN(new_n321));
  INV_X1    g120(.A(G120gat), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT1), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT69), .B(G120gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G113gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n323), .B1(new_n321), .B2(new_n322), .ZN(new_n328));
  INV_X1    g127(.A(new_n320), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n302), .A2(new_n308), .ZN(new_n332));
  INV_X1    g131(.A(G155gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT78), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT78), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G155gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n336), .A3(G162gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT2), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT79), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(new_n340), .A3(new_n309), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n319), .A2(new_n331), .A3(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n327), .A2(new_n330), .ZN(new_n343));
  INV_X1    g142(.A(new_n318), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT5), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n309), .B(new_n351), .C1(new_n311), .C2(new_n317), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n339), .A2(KEYINPUT80), .A3(new_n351), .A4(new_n309), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n319), .A2(KEYINPUT3), .A3(new_n341), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(new_n357), .A3(new_n331), .ZN(new_n358));
  OR3_X1    g157(.A1(new_n331), .A2(new_n318), .A3(KEYINPUT4), .ZN(new_n359));
  OAI21_X1  g158(.A(KEYINPUT4), .B1(new_n331), .B2(new_n318), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n358), .A2(new_n361), .A3(new_n347), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT81), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n350), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n350), .B1(new_n362), .B2(new_n363), .ZN(new_n366));
  XNOR2_X1  g165(.A(G1gat), .B(G29gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(G85gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT0), .B(G57gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n365), .A2(new_n366), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT6), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n371), .B1(new_n365), .B2(new_n366), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT6), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n373), .B1(new_n376), .B2(new_n372), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n298), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G78gat), .B(G106gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(G22gat), .B(G50gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n351), .B1(new_n255), .B2(KEYINPUT29), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n318), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT29), .B1(new_n354), .B2(new_n355), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n385), .B1(new_n386), .B2(new_n281), .ZN(new_n387));
  INV_X1    g186(.A(G228gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n388), .A2(new_n219), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT83), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n387), .A2(KEYINPUT83), .A3(new_n390), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n384), .A2(new_n319), .A3(new_n341), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n389), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n386), .A2(new_n281), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n383), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n383), .ZN(new_n402));
  AOI211_X1 g201(.A(new_n402), .B(new_n399), .C1(new_n393), .C2(new_n394), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n382), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n387), .A2(KEYINPUT83), .A3(new_n390), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT83), .B1(new_n387), .B2(new_n390), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n400), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n402), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n395), .A2(new_n383), .A3(new_n400), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n409), .A3(new_n381), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT34), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n343), .B1(new_n275), .B2(new_n256), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n331), .B(new_n217), .C1(new_n241), .C2(new_n246), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G227gat), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n416), .A2(new_n219), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n412), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  AOI211_X1 g218(.A(KEYINPUT34), .B(new_n417), .C1(new_n413), .C2(new_n414), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n413), .A2(new_n417), .A3(new_n414), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT32), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT33), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  XOR2_X1   g224(.A(G15gat), .B(G43gat), .Z(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT70), .ZN(new_n427));
  XOR2_X1   g226(.A(G71gat), .B(G99gat), .Z(new_n428));
  XNOR2_X1  g227(.A(new_n427), .B(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n423), .A2(new_n425), .A3(new_n430), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n422), .B(KEYINPUT32), .C1(new_n424), .C2(new_n429), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n421), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT72), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT72), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n421), .A2(new_n431), .A3(new_n435), .A4(new_n432), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n431), .A2(new_n432), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT71), .ZN(new_n439));
  INV_X1    g238(.A(new_n421), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT71), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n431), .A2(new_n441), .A3(new_n432), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n439), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n411), .A2(new_n437), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT35), .B1(new_n378), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT35), .B1(new_n404), .B2(new_n410), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n434), .A2(new_n436), .B1(new_n440), .B2(new_n438), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n362), .A2(new_n363), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n448), .A2(KEYINPUT5), .A3(new_n349), .ZN(new_n449));
  XOR2_X1   g248(.A(new_n370), .B(KEYINPUT85), .Z(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n364), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n374), .A2(new_n375), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n373), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n298), .A2(new_n446), .A3(new_n447), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n445), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT73), .ZN(new_n456));
  AND4_X1   g255(.A1(new_n456), .A2(new_n437), .A3(KEYINPUT36), .A4(new_n443), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n437), .A2(new_n443), .A3(KEYINPUT36), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n456), .B1(new_n447), .B2(KEYINPUT36), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT84), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n408), .A2(new_n409), .A3(new_n381), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n381), .B1(new_n408), .B2(new_n409), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n404), .A2(KEYINPUT84), .A3(new_n410), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n378), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT40), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n347), .B1(new_n358), .B2(new_n361), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT39), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n450), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT39), .B1(new_n346), .B2(new_n348), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n468), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n475), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n477), .A2(KEYINPUT40), .A3(new_n472), .A4(new_n471), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n476), .A2(new_n478), .A3(new_n451), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n294), .A2(new_n479), .A3(new_n297), .ZN(new_n480));
  XNOR2_X1  g279(.A(KEYINPUT86), .B(KEYINPUT38), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT37), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n278), .A2(new_n483), .A3(new_n284), .A4(new_n285), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n484), .A2(new_n290), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n286), .A2(KEYINPUT37), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n282), .A2(new_n272), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n481), .B1(new_n488), .B2(KEYINPUT37), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n484), .A2(new_n290), .A3(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n373), .A2(new_n490), .A3(new_n452), .A4(new_n293), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n480), .B(new_n411), .C1(new_n487), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n467), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n455), .B1(new_n460), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G229gat), .A2(G233gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(G15gat), .B(G22gat), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n496), .A2(KEYINPUT91), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n497), .A2(G1gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(G1gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT16), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n498), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(G8gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(G29gat), .A2(G36gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(KEYINPUT14), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT89), .ZN(new_n507));
  INV_X1    g306(.A(G29gat), .ZN(new_n508));
  INV_X1    g307(.A(G36gat), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G43gat), .B(G50gat), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(KEYINPUT15), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(KEYINPUT15), .B2(new_n511), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g313(.A(KEYINPUT15), .B(new_n511), .C1(new_n506), .C2(new_n510), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT90), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT90), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n514), .A2(new_n518), .A3(new_n515), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n504), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT17), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n517), .A2(new_n522), .A3(new_n519), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n516), .A2(KEYINPUT17), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n504), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n495), .B(new_n521), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT18), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n523), .A2(new_n524), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n520), .B1(new_n530), .B2(new_n504), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(KEYINPUT18), .A3(new_n495), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n519), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(new_n526), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(new_n495), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G169gat), .B(G197gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(new_n314), .ZN(new_n539));
  XOR2_X1   g338(.A(KEYINPUT87), .B(KEYINPUT11), .Z(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT88), .B(G113gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT12), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n529), .A2(new_n532), .A3(new_n537), .A4(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n527), .A2(new_n528), .B1(new_n534), .B2(new_n536), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n544), .B1(new_n547), .B2(new_n532), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n494), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT93), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT93), .B1(new_n494), .B2(new_n549), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G64gat), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n555), .A2(G57gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT95), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n555), .A2(G57gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT95), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n557), .B1(new_n560), .B2(new_n556), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT96), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G71gat), .B(G78gat), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n565), .B(KEYINPUT94), .Z(new_n566));
  NAND2_X1  g365(.A1(new_n561), .A2(new_n562), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n563), .A2(new_n564), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n566), .B1(new_n558), .B2(new_n556), .ZN(new_n569));
  INV_X1    g368(.A(new_n564), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT98), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n526), .B1(new_n573), .B2(KEYINPUT21), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT21), .B1(new_n568), .B2(new_n571), .ZN(new_n577));
  XNOR2_X1  g376(.A(G183gat), .B(G211gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT99), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n579), .B(KEYINPUT97), .Z(new_n580));
  XNOR2_X1  g379(.A(new_n577), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582));
  INV_X1    g381(.A(G127gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(new_n333), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n581), .B(new_n585), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n576), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n576), .A2(new_n586), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(KEYINPUT41), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT100), .ZN(new_n593));
  XOR2_X1   g392(.A(G134gat), .B(G162gat), .Z(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n595), .A2(KEYINPUT105), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(KEYINPUT105), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G99gat), .B(G106gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT103), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT104), .ZN(new_n601));
  NAND2_X1  g400(.A1(G85gat), .A2(G92gat), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT7), .B1(new_n602), .B2(KEYINPUT101), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(KEYINPUT101), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT102), .B1(G99gat), .B2(G106gat), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT8), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(KEYINPUT102), .A2(G99gat), .A3(G106gat), .ZN(new_n609));
  INV_X1    g408(.A(G85gat), .ZN(new_n610));
  INV_X1    g409(.A(G92gat), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n608), .A2(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n601), .A2(new_n605), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT104), .ZN(new_n614));
  INV_X1    g413(.A(new_n600), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n614), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n617), .A2(new_n605), .A3(new_n601), .A4(new_n612), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n530), .A2(new_n620), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n533), .A2(new_n619), .B1(KEYINPUT41), .B2(new_n591), .ZN(new_n622));
  XNOR2_X1  g421(.A(G190gat), .B(G218gat), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n621), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n624), .B1(new_n621), .B2(new_n622), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n598), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n627), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n629), .A2(new_n596), .A3(new_n625), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n619), .A2(new_n572), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n616), .A2(new_n618), .A3(new_n571), .A4(new_n568), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n573), .A2(KEYINPUT10), .A3(new_n619), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G230gat), .A2(G233gat), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(G176gat), .B(G204gat), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT106), .ZN(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n642), .B(new_n643), .Z(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n640), .B(new_n645), .C1(new_n639), .C2(new_n634), .ZN(new_n646));
  INV_X1    g445(.A(new_n639), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n636), .B2(new_n637), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n634), .A2(new_n639), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n644), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n589), .A2(new_n631), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n554), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n377), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g458(.A1(new_n655), .A2(new_n298), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n503), .A2(KEYINPUT42), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(KEYINPUT108), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT107), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT16), .B(G8gat), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n665), .B(new_n666), .Z(new_n667));
  AOI21_X1  g466(.A(new_n662), .B1(new_n660), .B2(new_n667), .ZN(G1325gat));
  AND3_X1   g467(.A1(new_n656), .A2(G15gat), .A3(new_n460), .ZN(new_n669));
  AOI21_X1  g468(.A(G15gat), .B1(new_n656), .B2(new_n447), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(G1326gat));
  INV_X1    g470(.A(new_n466), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n655), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT43), .B(G22gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  NOR3_X1   g474(.A1(new_n589), .A2(new_n631), .A3(new_n651), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n554), .A2(new_n508), .A3(new_n657), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT45), .ZN(new_n678));
  INV_X1    g477(.A(new_n631), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n494), .A2(KEYINPUT109), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n494), .A2(KEYINPUT109), .A3(KEYINPUT44), .A4(new_n679), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n546), .A2(new_n548), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n684), .A2(new_n589), .A3(new_n651), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(KEYINPUT110), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT110), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n682), .A2(new_n688), .A3(new_n683), .A4(new_n685), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n377), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n678), .B1(new_n508), .B2(new_n690), .ZN(G1328gat));
  INV_X1    g490(.A(new_n298), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n554), .A2(new_n509), .A3(new_n692), .A4(new_n676), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(KEYINPUT46), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(KEYINPUT46), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n298), .B1(new_n687), .B2(new_n689), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n694), .B(new_n695), .C1(new_n509), .C2(new_n696), .ZN(G1329gat));
  NAND2_X1  g496(.A1(new_n459), .A2(new_n458), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(KEYINPUT73), .B2(new_n458), .ZN(new_n699));
  OAI21_X1  g498(.A(G43gat), .B1(new_n686), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n554), .A2(new_n676), .ZN(new_n701));
  INV_X1    g500(.A(new_n447), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n702), .A2(G43gat), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n700), .B(KEYINPUT47), .C1(new_n701), .C2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n701), .A2(new_n703), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n687), .A2(new_n689), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n460), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n705), .B1(new_n707), .B2(G43gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n704), .B1(new_n708), .B2(new_n709), .ZN(G1330gat));
  INV_X1    g509(.A(KEYINPUT48), .ZN(new_n711));
  INV_X1    g510(.A(G50gat), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n712), .B1(new_n706), .B2(new_n466), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT112), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(new_n554), .B2(new_n676), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n714), .B(new_n676), .C1(new_n552), .C2(new_n553), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n716), .A2(new_n712), .A3(new_n466), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n711), .B1(new_n713), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G50gat), .B1(new_n686), .B2(new_n411), .ZN(new_n720));
  OAI211_X1 g519(.A(KEYINPUT48), .B(new_n720), .C1(new_n715), .C2(new_n717), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(G1331gat));
  NAND2_X1  g521(.A1(new_n684), .A2(new_n651), .ZN(new_n723));
  INV_X1    g522(.A(new_n589), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n723), .A2(new_n724), .A3(new_n679), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n494), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(new_n377), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT113), .B(G57gat), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1332gat));
  NOR2_X1   g528(.A1(new_n726), .A2(new_n298), .ZN(new_n730));
  NOR2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  AND2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n730), .B2(new_n731), .ZN(G1333gat));
  INV_X1    g533(.A(G71gat), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n726), .A2(new_n735), .A3(new_n699), .ZN(new_n736));
  INV_X1    g535(.A(new_n726), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n447), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n736), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n466), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G78gat), .ZN(G1335gat));
  NAND4_X1  g541(.A1(new_n494), .A2(new_n684), .A3(new_n724), .A4(new_n679), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n743), .A2(KEYINPUT51), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(KEYINPUT51), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n744), .A2(new_n651), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(new_n610), .A3(new_n657), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n682), .A2(new_n683), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n723), .A2(new_n589), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n749), .A2(new_n657), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n748), .B1(new_n751), .B2(new_n610), .ZN(G1336gat));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n682), .A2(new_n692), .A3(new_n683), .A4(new_n750), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G92gat), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n753), .B1(new_n755), .B2(KEYINPUT114), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n692), .A2(new_n611), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n746), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n756), .B(new_n758), .ZN(G1337gat));
  OR3_X1    g558(.A1(new_n746), .A2(G99gat), .A3(new_n702), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n749), .A2(new_n460), .A3(new_n750), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(G99gat), .B1(new_n761), .B2(new_n762), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n760), .B1(new_n763), .B2(new_n764), .ZN(G1338gat));
  NOR2_X1   g564(.A1(new_n411), .A2(G106gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n747), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n411), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n749), .A2(new_n768), .A3(new_n750), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G106gat), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n767), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n749), .A2(new_n466), .A3(new_n750), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n747), .A2(new_n766), .B1(new_n773), .B2(G106gat), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n772), .B1(new_n774), .B2(new_n771), .ZN(G1339gat));
  NAND2_X1  g574(.A1(new_n654), .A2(new_n684), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n636), .A2(new_n637), .A3(new_n647), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n640), .A2(KEYINPUT54), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n645), .B1(new_n648), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n778), .A2(KEYINPUT55), .A3(new_n780), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n646), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n531), .A2(new_n495), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n534), .A2(new_n536), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n543), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n545), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n679), .B1(new_n785), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n724), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n651), .A2(new_n545), .A3(new_n788), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n631), .ZN(new_n793));
  INV_X1    g592(.A(new_n785), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(new_n794), .B2(new_n549), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n776), .B1(new_n791), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n684), .A2(new_n785), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n790), .B(new_n724), .C1(new_n799), .C2(new_n793), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n800), .A2(KEYINPUT116), .A3(new_n776), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n798), .A2(new_n657), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n444), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(new_n692), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n806), .A2(new_n321), .A3(new_n549), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n803), .A2(new_n447), .A3(new_n298), .A4(new_n672), .ZN(new_n808));
  OAI21_X1  g607(.A(G113gat), .B1(new_n808), .B2(new_n684), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(G1340gat));
  NOR2_X1   g609(.A1(new_n652), .A2(new_n325), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n806), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(G120gat), .B1(new_n808), .B2(new_n652), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(G1341gat));
  NOR3_X1   g613(.A1(new_n808), .A2(new_n583), .A3(new_n724), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n806), .A2(new_n589), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n815), .B1(new_n816), .B2(new_n583), .ZN(G1342gat));
  OAI21_X1  g616(.A(G134gat), .B1(new_n808), .B2(new_n631), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI211_X1 g619(.A(KEYINPUT117), .B(G134gat), .C1(new_n808), .C2(new_n631), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n692), .A2(new_n631), .A3(G134gat), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OR3_X1    g622(.A1(new_n805), .A2(KEYINPUT56), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT56), .B1(new_n805), .B2(new_n823), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n820), .A2(new_n821), .A3(new_n824), .A4(new_n825), .ZN(G1343gat));
  AND2_X1   g625(.A1(new_n798), .A2(new_n801), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n828), .A3(new_n657), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n460), .A2(new_n411), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n831), .B1(new_n802), .B2(KEYINPUT119), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n684), .A2(G141gat), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n829), .A2(new_n832), .A3(new_n298), .A4(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n798), .A2(new_n835), .A3(new_n768), .A4(new_n801), .ZN(new_n836));
  INV_X1    g635(.A(new_n796), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT57), .B1(new_n837), .B2(new_n672), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n699), .A2(new_n657), .A3(new_n298), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT118), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n836), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(G141gat), .B1(new_n841), .B2(new_n684), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n834), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT58), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n834), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(G1344gat));
  NAND2_X1  g646(.A1(new_n829), .A2(new_n832), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n692), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n312), .A3(new_n651), .ZN(new_n850));
  XNOR2_X1  g649(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n851));
  AOI211_X1 g650(.A(KEYINPUT57), .B(new_n672), .C1(new_n800), .C2(new_n776), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n798), .A2(new_n768), .A3(new_n801), .ZN(new_n853));
  AOI211_X1 g652(.A(new_n652), .B(new_n852), .C1(new_n853), .C2(KEYINPUT57), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n840), .B(KEYINPUT121), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n851), .B1(new_n856), .B2(G148gat), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n652), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n858), .A2(KEYINPUT59), .A3(new_n312), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n850), .B1(new_n857), .B2(new_n859), .ZN(G1345gat));
  INV_X1    g659(.A(new_n310), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n841), .A2(new_n861), .A3(new_n724), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n849), .A2(new_n589), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(new_n861), .ZN(G1346gat));
  OAI21_X1  g663(.A(G162gat), .B1(new_n841), .B2(new_n631), .ZN(new_n865));
  INV_X1    g664(.A(G162gat), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n679), .A2(new_n866), .A3(new_n298), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n865), .B1(new_n848), .B2(new_n867), .ZN(G1347gat));
  NOR2_X1   g667(.A1(new_n657), .A2(new_n298), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n798), .A2(new_n801), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n804), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n684), .A2(G169gat), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT122), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n869), .B(KEYINPUT123), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n875), .A2(new_n447), .A3(new_n672), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n827), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(G169gat), .B1(new_n877), .B2(new_n684), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n874), .A2(new_n878), .ZN(G1348gat));
  INV_X1    g678(.A(G176gat), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n877), .A2(new_n880), .A3(new_n652), .ZN(new_n881));
  INV_X1    g680(.A(new_n871), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n651), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n881), .B1(new_n883), .B2(new_n880), .ZN(G1349gat));
  OAI21_X1  g683(.A(G183gat), .B1(new_n877), .B2(new_n724), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n724), .A2(new_n208), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n885), .B(KEYINPUT124), .C1(new_n871), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT60), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n871), .A2(new_n886), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT60), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n889), .A2(KEYINPUT124), .A3(new_n890), .A4(new_n885), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n888), .A2(new_n891), .ZN(G1350gat));
  NAND3_X1  g691(.A1(new_n882), .A2(new_n221), .A3(new_n679), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n827), .A2(new_n679), .A3(new_n876), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n894), .A2(new_n895), .A3(G190gat), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n894), .B2(G190gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n893), .B1(new_n896), .B2(new_n897), .ZN(G1351gat));
  NAND2_X1  g697(.A1(new_n853), .A2(KEYINPUT57), .ZN(new_n899));
  INV_X1    g698(.A(new_n852), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n875), .A2(new_n699), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(G197gat), .B1(new_n902), .B2(new_n684), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n798), .A2(new_n801), .A3(new_n830), .A4(new_n869), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n684), .A2(G197gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(G1352gat));
  INV_X1    g705(.A(G204gat), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n907), .B1(new_n854), .B2(new_n901), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n651), .A2(new_n907), .ZN(new_n909));
  OR3_X1    g708(.A1(new_n904), .A2(KEYINPUT62), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT62), .B1(new_n904), .B2(new_n909), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(KEYINPUT125), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n899), .A2(new_n651), .A3(new_n900), .A4(new_n901), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(G204gat), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT125), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n915), .A2(new_n916), .A3(new_n911), .A4(new_n910), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n913), .A2(new_n917), .ZN(G1353gat));
  NAND4_X1  g717(.A1(new_n899), .A2(new_n589), .A3(new_n900), .A4(new_n901), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n919), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT63), .B1(new_n919), .B2(G211gat), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n589), .A2(new_n250), .ZN(new_n922));
  OAI22_X1  g721(.A1(new_n920), .A2(new_n921), .B1(new_n904), .B2(new_n922), .ZN(G1354gat));
  NOR2_X1   g722(.A1(new_n902), .A2(KEYINPUT127), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n679), .A2(G218gat), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n902), .A2(KEYINPUT127), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n251), .B1(new_n904), .B2(new_n631), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT126), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n928), .A2(KEYINPUT126), .ZN(new_n930));
  AOI22_X1  g729(.A1(new_n926), .A2(new_n927), .B1(new_n929), .B2(new_n930), .ZN(G1355gat));
endmodule


