

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n545, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739;

  INV_X1 U372 ( .A(n531), .ZN(n350) );
  INV_X1 U373 ( .A(KEYINPUT48), .ZN(n352) );
  XNOR2_X1 U374 ( .A(n548), .B(n547), .ZN(n614) );
  XNOR2_X1 U375 ( .A(n543), .B(n355), .ZN(n354) );
  INV_X1 U376 ( .A(KEYINPUT34), .ZN(n355) );
  OR2_X1 U377 ( .A1(n564), .A2(n577), .ZN(n536) );
  BUF_X1 U378 ( .A(n663), .Z(n353) );
  XNOR2_X1 U379 ( .A(n489), .B(n484), .ZN(n663) );
  OR2_X1 U380 ( .A1(n643), .A2(G902), .ZN(n390) );
  AND2_X1 U381 ( .A1(n598), .A2(n467), .ZN(n375) );
  XNOR2_X1 U382 ( .A(n726), .B(G146), .ZN(n406) );
  BUF_X1 U383 ( .A(n424), .Z(n728) );
  NOR2_X2 U384 ( .A1(G953), .A2(G237), .ZN(n446) );
  INV_X1 U385 ( .A(G953), .ZN(n424) );
  INV_X2 U386 ( .A(G125), .ZN(n358) );
  AND2_X2 U387 ( .A1(n351), .A2(n350), .ZN(n727) );
  XNOR2_X1 U388 ( .A(n522), .B(n352), .ZN(n351) );
  AND2_X4 U389 ( .A1(n660), .A2(n597), .ZN(n647) );
  NAND2_X1 U390 ( .A1(n354), .A2(n545), .ZN(n548) );
  INV_X2 U391 ( .A(n669), .ZN(n486) );
  NOR2_X1 U392 ( .A1(n735), .A2(n739), .ZN(n519) );
  XNOR2_X1 U393 ( .A(G107), .B(G104), .ZN(n417) );
  XNOR2_X2 U394 ( .A(n486), .B(KEYINPUT6), .ZN(n577) );
  NOR2_X1 U395 ( .A1(n586), .A2(n589), .ZN(n588) );
  XNOR2_X1 U396 ( .A(n585), .B(n584), .ZN(n589) );
  AND2_X1 U397 ( .A1(n515), .A2(n473), .ZN(n713) );
  XNOR2_X1 U398 ( .A(KEYINPUT71), .B(KEYINPUT4), .ZN(n429) );
  OR2_X1 U399 ( .A1(n490), .A2(n489), .ZN(n517) );
  NOR2_X4 U400 ( .A1(n517), .A2(n493), .ZN(n714) );
  NOR2_X1 U401 ( .A1(n524), .A2(n492), .ZN(n483) );
  XNOR2_X2 U402 ( .A(n472), .B(KEYINPUT108), .ZN(n737) );
  XNOR2_X2 U403 ( .A(n358), .B(G146), .ZN(n430) );
  XNOR2_X1 U404 ( .A(n413), .B(n412), .ZN(n414) );
  AND2_X1 U405 ( .A1(n569), .A2(n478), .ZN(n415) );
  INV_X1 U406 ( .A(KEYINPUT30), .ZN(n412) );
  OR2_X1 U407 ( .A1(n669), .A2(n676), .ZN(n413) );
  INV_X1 U408 ( .A(KEYINPUT44), .ZN(n562) );
  NOR2_X1 U409 ( .A1(n728), .A2(G952), .ZN(n654) );
  XNOR2_X1 U410 ( .A(n588), .B(n587), .ZN(n660) );
  XNOR2_X1 U411 ( .A(n511), .B(KEYINPUT109), .ZN(n512) );
  INV_X1 U412 ( .A(KEYINPUT40), .ZN(n511) );
  XNOR2_X1 U413 ( .A(n483), .B(n482), .ZN(n485) );
  INV_X1 U414 ( .A(KEYINPUT36), .ZN(n482) );
  INV_X1 U415 ( .A(KEYINPUT107), .ZN(n439) );
  XOR2_X1 U416 ( .A(n405), .B(n420), .Z(n356) );
  AND2_X1 U417 ( .A1(n581), .A2(n605), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n609), .B(KEYINPUT85), .ZN(n503) );
  XNOR2_X1 U419 ( .A(KEYINPUT23), .B(KEYINPUT81), .ZN(n360) );
  BUF_X1 U420 ( .A(n533), .Z(n664) );
  XNOR2_X1 U421 ( .A(KEYINPUT10), .B(n430), .ZN(n359) );
  NOR2_X1 U422 ( .A1(n533), .A2(n489), .ZN(n569) );
  NOR2_X1 U423 ( .A1(n507), .A2(n529), .ZN(n440) );
  INV_X1 U424 ( .A(KEYINPUT80), .ZN(n587) );
  NOR2_X1 U425 ( .A1(n507), .A2(n677), .ZN(n510) );
  OR2_X2 U426 ( .A1(n485), .A2(n353), .ZN(n609) );
  XNOR2_X1 U427 ( .A(n513), .B(n512), .ZN(n735) );
  BUF_X1 U428 ( .A(n737), .Z(n738) );
  INV_X1 U429 ( .A(KEYINPUT82), .ZN(n476) );
  INV_X1 U430 ( .A(n359), .ZN(n442) );
  XNOR2_X1 U431 ( .A(n442), .B(n360), .ZN(n367) );
  NAND2_X1 U432 ( .A1(G234), .A2(n424), .ZN(n361) );
  XOR2_X1 U433 ( .A(KEYINPUT8), .B(n361), .Z(n462) );
  NAND2_X1 U434 ( .A1(G221), .A2(n462), .ZN(n365) );
  XOR2_X1 U435 ( .A(KEYINPUT24), .B(G140), .Z(n363) );
  XNOR2_X1 U436 ( .A(G137), .B(G128), .ZN(n362) );
  XOR2_X1 U437 ( .A(n363), .B(n362), .Z(n364) );
  XNOR2_X1 U438 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U439 ( .A(n367), .B(n366), .ZN(n369) );
  XNOR2_X1 U440 ( .A(G119), .B(G110), .ZN(n418) );
  XNOR2_X1 U441 ( .A(n418), .B(KEYINPUT84), .ZN(n368) );
  XNOR2_X1 U442 ( .A(n369), .B(n368), .ZN(n598) );
  INV_X1 U443 ( .A(G902), .ZN(n467) );
  XOR2_X1 U444 ( .A(KEYINPUT25), .B(KEYINPUT93), .Z(n373) );
  XNOR2_X1 U445 ( .A(KEYINPUT15), .B(G902), .ZN(n434) );
  NAND2_X1 U446 ( .A1(n434), .A2(G234), .ZN(n370) );
  XNOR2_X1 U447 ( .A(n370), .B(KEYINPUT20), .ZN(n371) );
  XNOR2_X1 U448 ( .A(KEYINPUT92), .B(n371), .ZN(n376) );
  NAND2_X1 U449 ( .A1(G217), .A2(n376), .ZN(n372) );
  XOR2_X1 U450 ( .A(n373), .B(n372), .Z(n374) );
  XNOR2_X1 U451 ( .A(n375), .B(n374), .ZN(n477) );
  AND2_X1 U452 ( .A1(n376), .A2(G221), .ZN(n378) );
  INV_X1 U453 ( .A(KEYINPUT21), .ZN(n377) );
  XNOR2_X1 U454 ( .A(n378), .B(n377), .ZN(n661) );
  OR2_X2 U455 ( .A1(n477), .A2(n661), .ZN(n533) );
  XNOR2_X2 U456 ( .A(G143), .B(G128), .ZN(n423) );
  INV_X1 U457 ( .A(G134), .ZN(n379) );
  XNOR2_X1 U458 ( .A(n423), .B(n379), .ZN(n460) );
  INV_X1 U459 ( .A(n460), .ZN(n382) );
  XNOR2_X1 U460 ( .A(KEYINPUT72), .B(G137), .ZN(n380) );
  XNOR2_X1 U461 ( .A(n429), .B(n380), .ZN(n381) );
  XNOR2_X2 U462 ( .A(n382), .B(n381), .ZN(n726) );
  XNOR2_X1 U463 ( .A(G140), .B(G131), .ZN(n441) );
  XNOR2_X1 U464 ( .A(n417), .B(n441), .ZN(n386) );
  XNOR2_X1 U465 ( .A(G110), .B(G101), .ZN(n384) );
  NAND2_X1 U466 ( .A1(n728), .A2(G227), .ZN(n383) );
  XNOR2_X1 U467 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U468 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U469 ( .A(n406), .B(n387), .ZN(n643) );
  INV_X1 U470 ( .A(KEYINPUT74), .ZN(n388) );
  XNOR2_X1 U471 ( .A(n388), .B(G469), .ZN(n389) );
  XNOR2_X2 U472 ( .A(n390), .B(n389), .ZN(n489) );
  NAND2_X1 U473 ( .A1(G237), .A2(G234), .ZN(n391) );
  XNOR2_X1 U474 ( .A(n391), .B(KEYINPUT14), .ZN(n394) );
  NAND2_X1 U475 ( .A1(n394), .A2(G952), .ZN(n392) );
  XOR2_X1 U476 ( .A(KEYINPUT91), .B(n392), .Z(n691) );
  INV_X1 U477 ( .A(n691), .ZN(n393) );
  NAND2_X1 U478 ( .A1(n393), .A2(n728), .ZN(n539) );
  NAND2_X1 U479 ( .A1(G902), .A2(n394), .ZN(n537) );
  NOR2_X1 U480 ( .A1(G900), .A2(n537), .ZN(n395) );
  NAND2_X1 U481 ( .A1(G953), .A2(n395), .ZN(n396) );
  XOR2_X1 U482 ( .A(KEYINPUT105), .B(n396), .Z(n397) );
  NAND2_X1 U483 ( .A1(n539), .A2(n397), .ZN(n478) );
  NAND2_X1 U484 ( .A1(n446), .A2(G210), .ZN(n399) );
  XNOR2_X1 U485 ( .A(G119), .B(G131), .ZN(n398) );
  XNOR2_X1 U486 ( .A(n399), .B(n398), .ZN(n401) );
  XNOR2_X1 U487 ( .A(KEYINPUT79), .B(KEYINPUT5), .ZN(n400) );
  XNOR2_X1 U488 ( .A(n401), .B(n400), .ZN(n405) );
  XNOR2_X1 U489 ( .A(G116), .B(G113), .ZN(n402) );
  XNOR2_X1 U490 ( .A(n402), .B(KEYINPUT3), .ZN(n404) );
  XNOR2_X1 U491 ( .A(G101), .B(KEYINPUT75), .ZN(n403) );
  XNOR2_X1 U492 ( .A(n404), .B(n403), .ZN(n420) );
  XNOR2_X1 U493 ( .A(n406), .B(n356), .ZN(n616) );
  OR2_X2 U494 ( .A1(n616), .A2(G902), .ZN(n410) );
  XNOR2_X1 U495 ( .A(KEYINPUT95), .B(G472), .ZN(n408) );
  INV_X1 U496 ( .A(KEYINPUT77), .ZN(n407) );
  XNOR2_X1 U497 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X2 U498 ( .A(n410), .B(n409), .ZN(n669) );
  INV_X1 U499 ( .A(G237), .ZN(n411) );
  NAND2_X1 U500 ( .A1(n467), .A2(n411), .ZN(n435) );
  AND2_X1 U501 ( .A1(n435), .A2(G214), .ZN(n676) );
  NAND2_X1 U502 ( .A1(n415), .A2(n414), .ZN(n507) );
  XNOR2_X1 U503 ( .A(KEYINPUT16), .B(G122), .ZN(n416) );
  XNOR2_X1 U504 ( .A(n417), .B(n416), .ZN(n419) );
  XNOR2_X1 U505 ( .A(n419), .B(n418), .ZN(n421) );
  XNOR2_X1 U506 ( .A(n421), .B(n420), .ZN(n630) );
  XNOR2_X1 U507 ( .A(KEYINPUT18), .B(KEYINPUT88), .ZN(n422) );
  XNOR2_X1 U508 ( .A(n423), .B(n422), .ZN(n428) );
  XNOR2_X1 U509 ( .A(KEYINPUT89), .B(KEYINPUT17), .ZN(n426) );
  NAND2_X1 U510 ( .A1(n424), .A2(G224), .ZN(n425) );
  XNOR2_X1 U511 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U512 ( .A(n428), .B(n427), .ZN(n432) );
  XNOR2_X1 U513 ( .A(n429), .B(n430), .ZN(n431) );
  XNOR2_X1 U514 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U515 ( .A(n630), .B(n433), .ZN(n651) );
  INV_X1 U516 ( .A(n434), .ZN(n593) );
  OR2_X1 U517 ( .A1(n651), .A2(n593), .ZN(n438) );
  NAND2_X1 U518 ( .A1(n435), .A2(G210), .ZN(n436) );
  XNOR2_X1 U519 ( .A(n436), .B(KEYINPUT90), .ZN(n437) );
  XNOR2_X2 U520 ( .A(n438), .B(n437), .ZN(n529) );
  XNOR2_X1 U521 ( .A(n440), .B(n439), .ZN(n471) );
  XNOR2_X1 U522 ( .A(n442), .B(n441), .ZN(n725) );
  XOR2_X1 U523 ( .A(KEYINPUT99), .B(KEYINPUT12), .Z(n444) );
  XNOR2_X1 U524 ( .A(G122), .B(G143), .ZN(n443) );
  XNOR2_X1 U525 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U526 ( .A(n725), .B(n445), .ZN(n453) );
  XOR2_X1 U527 ( .A(KEYINPUT98), .B(KEYINPUT11), .Z(n448) );
  NAND2_X1 U528 ( .A1(n446), .A2(G214), .ZN(n447) );
  XNOR2_X1 U529 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U530 ( .A(n449), .B(KEYINPUT97), .Z(n451) );
  XNOR2_X1 U531 ( .A(G113), .B(G104), .ZN(n450) );
  XOR2_X1 U532 ( .A(n451), .B(n450), .Z(n452) );
  XNOR2_X1 U533 ( .A(n453), .B(n452), .ZN(n636) );
  NAND2_X1 U534 ( .A1(n636), .A2(n467), .ZN(n457) );
  XOR2_X1 U535 ( .A(KEYINPUT13), .B(KEYINPUT101), .Z(n455) );
  XNOR2_X1 U536 ( .A(KEYINPUT100), .B(G475), .ZN(n454) );
  XOR2_X1 U537 ( .A(n455), .B(n454), .Z(n456) );
  XNOR2_X1 U538 ( .A(n457), .B(n456), .ZN(n515) );
  XOR2_X1 U539 ( .A(KEYINPUT7), .B(G122), .Z(n459) );
  XNOR2_X1 U540 ( .A(G116), .B(G107), .ZN(n458) );
  XNOR2_X1 U541 ( .A(n459), .B(n458), .ZN(n461) );
  XNOR2_X1 U542 ( .A(n461), .B(n460), .ZN(n466) );
  NAND2_X1 U543 ( .A1(G217), .A2(n462), .ZN(n464) );
  XOR2_X1 U544 ( .A(KEYINPUT9), .B(KEYINPUT102), .Z(n463) );
  XNOR2_X1 U545 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U546 ( .A(n466), .B(n465), .ZN(n634) );
  NAND2_X1 U547 ( .A1(n634), .A2(n467), .ZN(n470) );
  XNOR2_X1 U548 ( .A(G478), .B(KEYINPUT104), .ZN(n468) );
  XOR2_X1 U549 ( .A(n468), .B(KEYINPUT103), .Z(n469) );
  XNOR2_X1 U550 ( .A(n470), .B(n469), .ZN(n514) );
  AND2_X1 U551 ( .A1(n515), .A2(n514), .ZN(n545) );
  NAND2_X1 U552 ( .A1(n471), .A2(n545), .ZN(n472) );
  INV_X1 U553 ( .A(n514), .ZN(n473) );
  OR2_X1 U554 ( .A1(n515), .A2(n473), .ZN(n718) );
  INV_X1 U555 ( .A(n718), .ZN(n708) );
  NOR2_X1 U556 ( .A1(n713), .A2(n708), .ZN(n682) );
  NAND2_X1 U557 ( .A1(n682), .A2(KEYINPUT47), .ZN(n474) );
  NAND2_X1 U558 ( .A1(n737), .A2(n474), .ZN(n475) );
  XNOR2_X1 U559 ( .A(n476), .B(n475), .ZN(n505) );
  BUF_X2 U560 ( .A(n477), .Z(n554) );
  INV_X1 U561 ( .A(n478), .ZN(n479) );
  NOR2_X1 U562 ( .A1(n661), .A2(n479), .ZN(n480) );
  AND2_X1 U563 ( .A1(n554), .A2(n480), .ZN(n487) );
  NAND2_X1 U564 ( .A1(n487), .A2(n713), .ZN(n481) );
  OR2_X2 U565 ( .A1(n481), .A2(n577), .ZN(n524) );
  OR2_X1 U566 ( .A1(n529), .A2(n676), .ZN(n492) );
  XNOR2_X1 U567 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n484) );
  NAND2_X1 U568 ( .A1(n487), .A2(n486), .ZN(n488) );
  XNOR2_X1 U569 ( .A(n488), .B(KEYINPUT28), .ZN(n490) );
  XNOR2_X1 U570 ( .A(KEYINPUT68), .B(KEYINPUT19), .ZN(n491) );
  XNOR2_X1 U571 ( .A(n492), .B(n491), .ZN(n541) );
  INV_X1 U572 ( .A(n541), .ZN(n493) );
  INV_X1 U573 ( .A(KEYINPUT70), .ZN(n495) );
  NOR2_X1 U574 ( .A1(n495), .A2(KEYINPUT47), .ZN(n494) );
  NAND2_X1 U575 ( .A1(n714), .A2(n494), .ZN(n497) );
  NAND2_X1 U576 ( .A1(n495), .A2(KEYINPUT47), .ZN(n496) );
  NAND2_X1 U577 ( .A1(n497), .A2(n496), .ZN(n498) );
  XNOR2_X1 U578 ( .A(KEYINPUT83), .B(n682), .ZN(n573) );
  NAND2_X1 U579 ( .A1(n498), .A2(n573), .ZN(n501) );
  INV_X1 U580 ( .A(n714), .ZN(n499) );
  NAND2_X1 U581 ( .A1(n499), .A2(KEYINPUT47), .ZN(n500) );
  NAND2_X1 U582 ( .A1(n501), .A2(n500), .ZN(n502) );
  NOR2_X1 U583 ( .A1(n503), .A2(n502), .ZN(n504) );
  NAND2_X1 U584 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U585 ( .A(n506), .B(KEYINPUT73), .ZN(n521) );
  INV_X1 U586 ( .A(KEYINPUT38), .ZN(n508) );
  XNOR2_X1 U587 ( .A(n529), .B(n508), .ZN(n677) );
  XNOR2_X1 U588 ( .A(KEYINPUT76), .B(KEYINPUT39), .ZN(n509) );
  XNOR2_X1 U589 ( .A(n510), .B(n509), .ZN(n523) );
  INV_X1 U590 ( .A(n713), .ZN(n716) );
  NOR2_X1 U591 ( .A1(n523), .A2(n716), .ZN(n513) );
  OR2_X1 U592 ( .A1(n515), .A2(n514), .ZN(n680) );
  OR2_X1 U593 ( .A1(n677), .A2(n676), .ZN(n681) );
  NOR2_X1 U594 ( .A1(n680), .A2(n681), .ZN(n516) );
  XNOR2_X1 U595 ( .A(n516), .B(KEYINPUT41), .ZN(n693) );
  NOR2_X1 U596 ( .A1(n693), .A2(n517), .ZN(n518) );
  XNOR2_X1 U597 ( .A(n518), .B(KEYINPUT42), .ZN(n739) );
  XNOR2_X1 U598 ( .A(n519), .B(KEYINPUT46), .ZN(n520) );
  NAND2_X1 U599 ( .A1(n521), .A2(n520), .ZN(n522) );
  OR2_X1 U600 ( .A1(n523), .A2(n718), .ZN(n722) );
  INV_X1 U601 ( .A(n524), .ZN(n526) );
  INV_X1 U602 ( .A(n353), .ZN(n576) );
  NOR2_X1 U603 ( .A1(n576), .A2(n676), .ZN(n525) );
  NAND2_X1 U604 ( .A1(n526), .A2(n525), .ZN(n528) );
  XNOR2_X1 U605 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n527) );
  XNOR2_X1 U606 ( .A(n528), .B(n527), .ZN(n530) );
  NAND2_X1 U607 ( .A1(n530), .A2(n529), .ZN(n606) );
  NAND2_X1 U608 ( .A1(n722), .A2(n606), .ZN(n531) );
  NAND2_X1 U609 ( .A1(n727), .A2(KEYINPUT2), .ZN(n586) );
  NOR2_X1 U610 ( .A1(n664), .A2(n663), .ZN(n535) );
  INV_X1 U611 ( .A(KEYINPUT78), .ZN(n534) );
  XNOR2_X1 U612 ( .A(n535), .B(n534), .ZN(n564) );
  XNOR2_X2 U613 ( .A(n536), .B(KEYINPUT33), .ZN(n675) );
  OR2_X1 U614 ( .A1(G898), .A2(n728), .ZN(n629) );
  OR2_X1 U615 ( .A1(n537), .A2(n629), .ZN(n538) );
  NAND2_X1 U616 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U617 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U618 ( .A(n542), .B(KEYINPUT0), .ZN(n565) );
  INV_X1 U619 ( .A(n565), .ZN(n570) );
  NAND2_X1 U620 ( .A1(n675), .A2(n570), .ZN(n543) );
  INV_X1 U621 ( .A(KEYINPUT35), .ZN(n547) );
  INV_X1 U622 ( .A(n680), .ZN(n550) );
  INV_X1 U623 ( .A(n661), .ZN(n549) );
  NAND2_X1 U624 ( .A1(n550), .A2(n549), .ZN(n551) );
  OR2_X1 U625 ( .A1(n565), .A2(n551), .ZN(n553) );
  XNOR2_X1 U626 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n552) );
  XNOR2_X2 U627 ( .A(n553), .B(n552), .ZN(n575) );
  NAND2_X1 U628 ( .A1(n554), .A2(n576), .ZN(n556) );
  INV_X1 U629 ( .A(n577), .ZN(n555) );
  NOR2_X1 U630 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U631 ( .A1(n575), .A2(n557), .ZN(n558) );
  XNOR2_X1 U632 ( .A(n558), .B(KEYINPUT32), .ZN(n608) );
  NAND2_X1 U633 ( .A1(n554), .A2(n669), .ZN(n559) );
  NOR2_X1 U634 ( .A1(n559), .A2(n576), .ZN(n560) );
  NAND2_X1 U635 ( .A1(n575), .A2(n560), .ZN(n604) );
  AND2_X1 U636 ( .A1(n608), .A2(n604), .ZN(n561) );
  NAND2_X1 U637 ( .A1(n614), .A2(n561), .ZN(n563) );
  XNOR2_X1 U638 ( .A(n563), .B(n562), .ZN(n582) );
  OR2_X1 U639 ( .A1(n565), .A2(n669), .ZN(n566) );
  OR2_X1 U640 ( .A1(n564), .A2(n566), .ZN(n568) );
  XOR2_X1 U641 ( .A(KEYINPUT96), .B(KEYINPUT31), .Z(n567) );
  XNOR2_X1 U642 ( .A(n568), .B(n567), .ZN(n719) );
  NAND2_X1 U643 ( .A1(n569), .A2(n570), .ZN(n571) );
  XNOR2_X1 U644 ( .A(n571), .B(KEYINPUT94), .ZN(n572) );
  OR2_X1 U645 ( .A1(n572), .A2(n486), .ZN(n703) );
  NAND2_X1 U646 ( .A1(n719), .A2(n703), .ZN(n574) );
  NAND2_X1 U647 ( .A1(n574), .A2(n573), .ZN(n581) );
  INV_X1 U648 ( .A(n575), .ZN(n580) );
  NOR2_X1 U649 ( .A1(n554), .A2(n576), .ZN(n578) );
  NAND2_X1 U650 ( .A1(n578), .A2(n577), .ZN(n579) );
  OR2_X1 U651 ( .A1(n580), .A2(n579), .ZN(n605) );
  NAND2_X1 U652 ( .A1(n582), .A2(n357), .ZN(n585) );
  INV_X1 U653 ( .A(KEYINPUT64), .ZN(n583) );
  XNOR2_X1 U654 ( .A(n583), .B(KEYINPUT45), .ZN(n584) );
  INV_X1 U655 ( .A(n589), .ZN(n622) );
  NAND2_X1 U656 ( .A1(n727), .A2(n622), .ZN(n658) );
  INV_X1 U657 ( .A(KEYINPUT67), .ZN(n590) );
  NAND2_X1 U658 ( .A1(n590), .A2(KEYINPUT2), .ZN(n591) );
  NAND2_X1 U659 ( .A1(n658), .A2(n591), .ZN(n592) );
  NAND2_X1 U660 ( .A1(n592), .A2(n593), .ZN(n596) );
  NAND2_X1 U661 ( .A1(n593), .A2(KEYINPUT2), .ZN(n594) );
  NAND2_X1 U662 ( .A1(n594), .A2(KEYINPUT67), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U664 ( .A1(n647), .A2(G217), .ZN(n600) );
  INV_X1 U665 ( .A(n598), .ZN(n599) );
  XNOR2_X1 U666 ( .A(n600), .B(n599), .ZN(n601) );
  NOR2_X2 U667 ( .A1(n601), .A2(n654), .ZN(n603) );
  INV_X1 U668 ( .A(KEYINPUT123), .ZN(n602) );
  XNOR2_X1 U669 ( .A(n603), .B(n602), .ZN(G66) );
  XNOR2_X1 U670 ( .A(n604), .B(G110), .ZN(G12) );
  XNOR2_X1 U671 ( .A(n605), .B(G101), .ZN(G3) );
  XNOR2_X1 U672 ( .A(n606), .B(G140), .ZN(G42) );
  XNOR2_X1 U673 ( .A(G119), .B(KEYINPUT126), .ZN(n607) );
  XNOR2_X1 U674 ( .A(n608), .B(n607), .ZN(G21) );
  INV_X1 U675 ( .A(n609), .ZN(n613) );
  XOR2_X1 U676 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n611) );
  XNOR2_X1 U677 ( .A(G125), .B(KEYINPUT37), .ZN(n610) );
  XNOR2_X1 U678 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U679 ( .A(n613), .B(n612), .ZN(G27) );
  XNOR2_X1 U680 ( .A(n614), .B(G122), .ZN(G24) );
  NAND2_X1 U681 ( .A1(n647), .A2(G472), .ZN(n618) );
  XNOR2_X1 U682 ( .A(KEYINPUT110), .B(KEYINPUT62), .ZN(n615) );
  XNOR2_X1 U683 ( .A(n616), .B(n615), .ZN(n617) );
  XNOR2_X1 U684 ( .A(n618), .B(n617), .ZN(n619) );
  NOR2_X2 U685 ( .A1(n619), .A2(n654), .ZN(n621) );
  XNOR2_X1 U686 ( .A(KEYINPUT111), .B(KEYINPUT63), .ZN(n620) );
  XNOR2_X1 U687 ( .A(n621), .B(n620), .ZN(G57) );
  NAND2_X1 U688 ( .A1(n622), .A2(n728), .ZN(n623) );
  XNOR2_X1 U689 ( .A(n623), .B(KEYINPUT125), .ZN(n628) );
  NAND2_X1 U690 ( .A1(G953), .A2(G224), .ZN(n624) );
  XNOR2_X1 U691 ( .A(KEYINPUT61), .B(n624), .ZN(n625) );
  NAND2_X1 U692 ( .A1(n625), .A2(G898), .ZN(n626) );
  XOR2_X1 U693 ( .A(KEYINPUT124), .B(n626), .Z(n627) );
  NOR2_X1 U694 ( .A1(n628), .A2(n627), .ZN(n632) );
  NAND2_X1 U695 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U696 ( .A(n632), .B(n631), .ZN(G69) );
  NAND2_X1 U697 ( .A1(n647), .A2(G478), .ZN(n633) );
  XOR2_X1 U698 ( .A(n634), .B(n633), .Z(n635) );
  NOR2_X1 U699 ( .A1(n635), .A2(n654), .ZN(G63) );
  NAND2_X1 U700 ( .A1(n647), .A2(G475), .ZN(n638) );
  XNOR2_X1 U701 ( .A(n636), .B(KEYINPUT59), .ZN(n637) );
  XNOR2_X1 U702 ( .A(n638), .B(n637), .ZN(n639) );
  NOR2_X2 U703 ( .A1(n639), .A2(n654), .ZN(n641) );
  XOR2_X1 U704 ( .A(KEYINPUT69), .B(KEYINPUT60), .Z(n640) );
  XNOR2_X1 U705 ( .A(n641), .B(n640), .ZN(G60) );
  NAND2_X1 U706 ( .A1(n647), .A2(G469), .ZN(n645) );
  XOR2_X1 U707 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n642) );
  XNOR2_X1 U708 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U709 ( .A(n645), .B(n644), .ZN(n646) );
  NOR2_X1 U710 ( .A1(n646), .A2(n654), .ZN(G54) );
  NAND2_X1 U711 ( .A1(n647), .A2(G210), .ZN(n653) );
  XNOR2_X1 U712 ( .A(KEYINPUT87), .B(KEYINPUT54), .ZN(n649) );
  XNOR2_X1 U713 ( .A(KEYINPUT55), .B(KEYINPUT86), .ZN(n648) );
  XNOR2_X1 U714 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U715 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U716 ( .A(n653), .B(n652), .ZN(n655) );
  NOR2_X2 U717 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U718 ( .A(n656), .B(KEYINPUT56), .ZN(G51) );
  INV_X1 U719 ( .A(KEYINPUT2), .ZN(n657) );
  NAND2_X1 U720 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U721 ( .A1(n660), .A2(n659), .ZN(n699) );
  AND2_X1 U722 ( .A1(n554), .A2(n661), .ZN(n662) );
  XNOR2_X1 U723 ( .A(KEYINPUT49), .B(n662), .ZN(n668) );
  NAND2_X1 U724 ( .A1(n664), .A2(n353), .ZN(n665) );
  XNOR2_X1 U725 ( .A(n665), .B(KEYINPUT120), .ZN(n666) );
  XNOR2_X1 U726 ( .A(KEYINPUT50), .B(n666), .ZN(n667) );
  NAND2_X1 U727 ( .A1(n668), .A2(n667), .ZN(n670) );
  NAND2_X1 U728 ( .A1(n670), .A2(n669), .ZN(n672) );
  NAND2_X1 U729 ( .A1(n564), .A2(n486), .ZN(n671) );
  NAND2_X1 U730 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U731 ( .A(KEYINPUT51), .B(n673), .Z(n674) );
  NOR2_X1 U732 ( .A1(n693), .A2(n674), .ZN(n688) );
  INV_X1 U733 ( .A(n675), .ZN(n686) );
  AND2_X1 U734 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U735 ( .A(KEYINPUT121), .B(n678), .Z(n679) );
  NOR2_X1 U736 ( .A1(n680), .A2(n679), .ZN(n684) );
  NOR2_X1 U737 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U738 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U739 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U740 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U741 ( .A(n689), .B(KEYINPUT52), .Z(n690) );
  XOR2_X1 U742 ( .A(KEYINPUT122), .B(n690), .Z(n692) );
  NOR2_X1 U743 ( .A1(n692), .A2(n691), .ZN(n697) );
  INV_X1 U744 ( .A(n693), .ZN(n694) );
  NAND2_X1 U745 ( .A1(n694), .A2(n675), .ZN(n695) );
  NAND2_X1 U746 ( .A1(n695), .A2(n728), .ZN(n696) );
  NOR2_X1 U747 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U748 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U749 ( .A(KEYINPUT53), .B(n700), .Z(G75) );
  NOR2_X1 U750 ( .A1(n703), .A2(n716), .ZN(n701) );
  XOR2_X1 U751 ( .A(KEYINPUT112), .B(n701), .Z(n702) );
  XNOR2_X1 U752 ( .A(G104), .B(n702), .ZN(G6) );
  NOR2_X1 U753 ( .A1(n703), .A2(n718), .ZN(n707) );
  XOR2_X1 U754 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n705) );
  XNOR2_X1 U755 ( .A(G107), .B(KEYINPUT113), .ZN(n704) );
  XNOR2_X1 U756 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U757 ( .A(n707), .B(n706), .ZN(G9) );
  XOR2_X1 U758 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n710) );
  NAND2_X1 U759 ( .A1(n714), .A2(n708), .ZN(n709) );
  XNOR2_X1 U760 ( .A(n710), .B(n709), .ZN(n712) );
  XOR2_X1 U761 ( .A(G128), .B(KEYINPUT114), .Z(n711) );
  XNOR2_X1 U762 ( .A(n712), .B(n711), .ZN(G30) );
  NAND2_X1 U763 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U764 ( .A(n715), .B(G146), .ZN(G48) );
  NOR2_X1 U765 ( .A1(n719), .A2(n716), .ZN(n717) );
  XOR2_X1 U766 ( .A(G113), .B(n717), .Z(G15) );
  NOR2_X1 U767 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U768 ( .A(KEYINPUT116), .B(n720), .Z(n721) );
  XNOR2_X1 U769 ( .A(G116), .B(n721), .ZN(G18) );
  INV_X1 U770 ( .A(n722), .ZN(n723) );
  XNOR2_X1 U771 ( .A(G134), .B(n723), .ZN(n724) );
  XNOR2_X1 U772 ( .A(n724), .B(KEYINPUT119), .ZN(G36) );
  XOR2_X1 U773 ( .A(n726), .B(n725), .Z(n730) );
  XNOR2_X1 U774 ( .A(n727), .B(n730), .ZN(n729) );
  NAND2_X1 U775 ( .A1(n729), .A2(n728), .ZN(n734) );
  XOR2_X1 U776 ( .A(n730), .B(G227), .Z(n731) );
  NAND2_X1 U777 ( .A1(n731), .A2(G900), .ZN(n732) );
  NAND2_X1 U778 ( .A1(n732), .A2(G953), .ZN(n733) );
  NAND2_X1 U779 ( .A1(n734), .A2(n733), .ZN(G72) );
  XNOR2_X1 U780 ( .A(G131), .B(KEYINPUT127), .ZN(n736) );
  XNOR2_X1 U781 ( .A(n736), .B(n735), .ZN(G33) );
  XNOR2_X1 U782 ( .A(n738), .B(G143), .ZN(G45) );
  XOR2_X1 U783 ( .A(G137), .B(n739), .Z(G39) );
endmodule

