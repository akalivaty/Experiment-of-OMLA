//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(KEYINPUT24), .ZN(new_n204));
  INV_X1    g003(.A(G169gat), .ZN(new_n205));
  INV_X1    g004(.A(G176gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G183gat), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n211), .A2(KEYINPUT24), .A3(new_n203), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n205), .A2(new_n206), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n208), .A2(new_n212), .A3(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(new_n214), .B2(new_n213), .ZN(new_n217));
  XOR2_X1   g016(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n213), .B(KEYINPUT65), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n216), .B(KEYINPUT25), .C1(new_n214), .C2(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g021(.A(KEYINPUT27), .B(G183gat), .Z(new_n223));
  OR2_X1    g022(.A1(new_n223), .A2(G190gat), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n224), .A2(KEYINPUT28), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n224), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n207), .B1(KEYINPUT26), .B2(new_n213), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(new_n220), .B2(KEYINPUT26), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n225), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n222), .A2(new_n230), .ZN(new_n231));
  OAI211_X1 g030(.A(KEYINPUT72), .B(new_n202), .C1(new_n231), .C2(KEYINPUT29), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT72), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n219), .A2(new_n221), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT29), .B1(new_n234), .B2(new_n229), .ZN(new_n235));
  INV_X1    g034(.A(new_n202), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n233), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT70), .B1(new_n222), .B2(new_n230), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n234), .A2(new_n239), .A3(new_n229), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n236), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n232), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G197gat), .B(G204gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT22), .ZN(new_n244));
  INV_X1    g043(.A(G211gat), .ZN(new_n245));
  INV_X1    g044(.A(G218gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(G211gat), .B(G218gat), .Z(new_n249));
  XOR2_X1   g048(.A(new_n248), .B(new_n249), .Z(new_n250));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n248), .A2(KEYINPUT69), .A3(new_n249), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n242), .A2(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(KEYINPUT71), .B(KEYINPUT29), .Z(new_n257));
  NAND4_X1  g056(.A1(new_n238), .A2(new_n257), .A3(new_n202), .A4(new_n240), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n231), .A2(new_n236), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n255), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G8gat), .B(G36gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(KEYINPUT73), .ZN(new_n264));
  XNOR2_X1  g063(.A(G64gat), .B(G92gat), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n264), .B(new_n265), .Z(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n266), .B1(new_n256), .B2(new_n261), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n268), .B1(KEYINPUT30), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT74), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n260), .B1(new_n255), .B2(new_n242), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT74), .B1(new_n273), .B2(new_n266), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT30), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n272), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G1gat), .B(G29gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT0), .ZN(new_n279));
  XNOR2_X1  g078(.A(G57gat), .B(G85gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT80), .ZN(new_n283));
  XOR2_X1   g082(.A(KEYINPUT78), .B(G155gat), .Z(new_n284));
  INV_X1    g083(.A(G162gat), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT2), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G155gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n285), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n287), .A2(new_n285), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G148gat), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n292), .A2(G141gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(KEYINPUT77), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT76), .B(G141gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(new_n292), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n286), .B(new_n291), .C1(new_n294), .C2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT75), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n290), .B1(new_n299), .B2(new_n288), .ZN(new_n300));
  XNOR2_X1  g099(.A(G141gat), .B(G148gat), .ZN(new_n301));
  OAI221_X1 g100(.A(new_n300), .B1(new_n299), .B2(new_n288), .C1(KEYINPUT2), .C2(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT3), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n298), .A2(new_n302), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT3), .ZN(new_n307));
  XNOR2_X1  g106(.A(G113gat), .B(G120gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT66), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n311));
  XNOR2_X1  g110(.A(G127gat), .B(G134gat), .ZN(new_n312));
  INV_X1    g111(.A(G120gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(KEYINPUT66), .A3(G113gat), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n310), .A2(new_n311), .A3(new_n312), .A4(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n312), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n316), .B1(KEYINPUT1), .B2(new_n308), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n305), .A2(new_n307), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT4), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(new_n306), .B2(new_n318), .ZN(new_n321));
  NAND2_X1  g120(.A1(G225gat), .A2(G233gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n318), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n303), .A2(KEYINPUT4), .A3(new_n323), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n319), .A2(new_n321), .A3(new_n322), .A4(new_n324), .ZN(new_n325));
  XOR2_X1   g124(.A(KEYINPUT79), .B(KEYINPUT5), .Z(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  OR2_X1    g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n306), .B(new_n318), .ZN(new_n329));
  INV_X1    g128(.A(new_n322), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n326), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n283), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT80), .B1(new_n325), .B2(new_n331), .ZN(new_n334));
  OAI211_X1 g133(.A(KEYINPUT6), .B(new_n282), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n333), .A2(new_n334), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT6), .B1(new_n337), .B2(new_n281), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n282), .B1(new_n333), .B2(new_n334), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n336), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT81), .B1(new_n277), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n337), .A2(new_n281), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT6), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(new_n343), .A3(new_n339), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n335), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT81), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n345), .A2(new_n346), .A3(new_n276), .A4(new_n270), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT83), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n348), .B1(new_n254), .B2(KEYINPUT29), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT29), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n252), .A2(KEYINPUT83), .A3(new_n350), .A4(new_n253), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n304), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(new_n306), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT84), .ZN(new_n354));
  INV_X1    g153(.A(new_n257), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n355), .B1(new_n303), .B2(new_n304), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n354), .B1(new_n356), .B2(new_n255), .ZN(new_n357));
  NAND2_X1  g156(.A1(G228gat), .A2(G233gat), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n356), .A2(new_n255), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT84), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n353), .A2(new_n357), .A3(new_n359), .A4(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n358), .B(KEYINPUT82), .ZN(new_n363));
  OR2_X1    g162(.A1(new_n250), .A2(new_n355), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n303), .B1(new_n364), .B2(new_n304), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G78gat), .B(G106gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT31), .B(G50gat), .ZN(new_n369));
  XOR2_X1   g168(.A(new_n368), .B(new_n369), .Z(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT85), .ZN(new_n373));
  INV_X1    g172(.A(G22gat), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n367), .A2(new_n371), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n370), .B1(new_n362), .B2(new_n366), .ZN(new_n377));
  OAI21_X1  g176(.A(G22gat), .B1(new_n377), .B2(KEYINPUT85), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G15gat), .B(G43gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(G71gat), .B(G99gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G227gat), .ZN(new_n385));
  INV_X1    g184(.A(G233gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n231), .A2(new_n323), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n318), .B1(new_n222), .B2(new_n230), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT32), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n384), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT67), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n389), .A2(new_n390), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n387), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT33), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n395), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n391), .A2(KEYINPUT67), .A3(KEYINPUT33), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n394), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n383), .A2(new_n398), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n391), .A2(new_n392), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n388), .A3(new_n390), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(KEYINPUT34), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n401), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n397), .A2(new_n395), .A3(new_n398), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT67), .B1(new_n391), .B2(KEYINPUT33), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n393), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n406), .B1(new_n411), .B2(new_n403), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n376), .B1(new_n375), .B2(new_n378), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n380), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n341), .A2(new_n347), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT35), .ZN(new_n417));
  INV_X1    g216(.A(new_n277), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT87), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n339), .A2(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(KEYINPUT87), .B(new_n282), .C1(new_n333), .C2(new_n334), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n338), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n335), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT35), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n418), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n415), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n417), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n407), .B1(new_n401), .B2(new_n404), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n411), .A2(new_n403), .A3(new_n406), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT68), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT36), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n413), .A2(KEYINPUT68), .A3(KEYINPUT36), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n374), .B1(new_n372), .B2(new_n373), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n377), .A2(KEYINPUT85), .A3(G22gat), .ZN(new_n436));
  OAI22_X1  g235(.A1(new_n435), .A2(new_n436), .B1(new_n371), .B2(new_n367), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n379), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT39), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n319), .A2(new_n321), .A3(new_n324), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT86), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n441), .A3(new_n330), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n441), .B1(new_n440), .B2(new_n330), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n439), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n444), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n329), .A2(new_n330), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n447), .A2(new_n439), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n442), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n445), .A2(new_n449), .A3(new_n281), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT40), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n445), .A2(new_n449), .A3(KEYINPUT40), .A4(new_n281), .ZN(new_n453));
  AND4_X1   g252(.A1(new_n420), .A2(new_n452), .A3(new_n421), .A4(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n438), .B1(new_n454), .B2(new_n277), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n272), .A2(new_n274), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT37), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n267), .B1(new_n262), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n258), .A2(new_n255), .A3(new_n259), .ZN(new_n459));
  OAI211_X1 g258(.A(KEYINPUT37), .B(new_n459), .C1(new_n242), .C2(new_n255), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT88), .ZN(new_n461));
  OR2_X1    g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT38), .B1(new_n460), .B2(new_n461), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n458), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n456), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n266), .B1(new_n273), .B2(KEYINPUT37), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n262), .A2(new_n457), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT38), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n465), .A2(new_n335), .A3(new_n422), .A4(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n434), .B1(new_n455), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n341), .A2(new_n347), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n438), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n427), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(G113gat), .B(G141gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(G197gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT11), .B(G169gat), .ZN(new_n477));
  XOR2_X1   g276(.A(new_n476), .B(new_n477), .Z(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(KEYINPUT12), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT93), .ZN(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G22gat), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT16), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n483), .A2(G1gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(G8gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n482), .A2(G1gat), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n485), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n486), .B1(new_n490), .B2(KEYINPUT91), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT91), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n485), .B(new_n492), .C1(G1gat), .C2(new_n482), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT92), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT92), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n491), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n489), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(G43gat), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT15), .B1(new_n499), .B2(G50gat), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(new_n499), .B2(G50gat), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n501), .B1(G29gat), .B2(G36gat), .ZN(new_n502));
  NOR3_X1   g301(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT90), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT15), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT89), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(new_n499), .B2(G50gat), .ZN(new_n510));
  INV_X1    g309(.A(G50gat), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(G43gat), .B2(new_n511), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n509), .A2(new_n499), .A3(G50gat), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n502), .A2(new_n507), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n506), .ZN(new_n516));
  INV_X1    g315(.A(G29gat), .ZN(new_n517));
  INV_X1    g316(.A(G36gat), .ZN(new_n518));
  OAI22_X1  g317(.A1(new_n516), .A2(new_n503), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n501), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n481), .B1(new_n498), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n497), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n496), .B1(new_n491), .B2(new_n493), .ZN(new_n525));
  OAI22_X1  g324(.A1(new_n524), .A2(new_n525), .B1(new_n488), .B2(new_n487), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(KEYINPUT93), .A3(new_n521), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n521), .B(KEYINPUT17), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n523), .A2(new_n527), .B1(new_n528), .B2(new_n498), .ZN(new_n529));
  NAND2_X1  g328(.A1(G229gat), .A2(G233gat), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT18), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n480), .B1(new_n531), .B2(KEYINPUT95), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n523), .A2(new_n527), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n528), .A2(new_n498), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(new_n530), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT18), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT94), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n533), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n527), .A3(KEYINPUT94), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n498), .A2(new_n522), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n530), .B(KEYINPUT13), .Z(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n529), .A2(KEYINPUT18), .A3(new_n530), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n532), .A2(new_n537), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT95), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n479), .B1(new_n537), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n543), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n533), .A2(new_n538), .B1(new_n522), .B2(new_n498), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n549), .B1(new_n550), .B2(new_n540), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n537), .A2(new_n545), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n548), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n546), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(G57gat), .B(G64gat), .Z(new_n555));
  INV_X1    g354(.A(G71gat), .ZN(new_n556));
  INV_X1    g355(.A(G78gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G71gat), .A2(G78gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n555), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G57gat), .B(G64gat), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n559), .B(new_n558), .C1(new_n564), .C2(new_n561), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n565), .A3(KEYINPUT96), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT96), .B1(new_n563), .B2(new_n565), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(KEYINPUT97), .B(KEYINPUT21), .Z(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(G127gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT96), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n555), .A2(new_n560), .A3(new_n562), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n560), .B1(new_n555), .B2(new_n562), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n566), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n526), .B1(KEYINPUT21), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n575), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(G155gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(G183gat), .B(G211gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n582), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G99gat), .B(G106gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT101), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(KEYINPUT101), .A2(G99gat), .A3(G106gat), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(KEYINPUT8), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(G85gat), .A2(G92gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT102), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT102), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n593), .A2(new_n598), .A3(new_n595), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G85gat), .A2(G92gat), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT100), .ZN(new_n602));
  OR3_X1    g401(.A1(new_n601), .A2(new_n602), .A3(KEYINPUT7), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(KEYINPUT7), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT99), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n602), .B1(new_n601), .B2(KEYINPUT7), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT99), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n601), .A2(new_n607), .A3(KEYINPUT7), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n603), .A2(new_n605), .A3(new_n606), .A4(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n588), .B1(new_n600), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT8), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n611), .B1(new_n589), .B2(new_n590), .ZN(new_n612));
  AOI211_X1 g411(.A(KEYINPUT102), .B(new_n594), .C1(new_n612), .C2(new_n592), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n598), .B1(new_n593), .B2(new_n595), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n588), .B(new_n609), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n528), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n521), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT41), .ZN(new_n621));
  NAND2_X1  g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n621), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT98), .ZN(new_n627));
  XOR2_X1   g426(.A(G134gat), .B(G162gat), .Z(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n625), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n587), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT106), .ZN(new_n634));
  NAND2_X1  g433(.A1(G230gat), .A2(G233gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n609), .B1(new_n613), .B2(new_n614), .ZN(new_n637));
  INV_X1    g436(.A(new_n588), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n577), .A2(new_n578), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n639), .A2(KEYINPUT103), .A3(new_n640), .A4(new_n615), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n639), .A2(new_n640), .A3(new_n615), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT103), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n580), .B1(new_n615), .B2(new_n639), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT10), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT104), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n646), .A2(new_n650), .A3(new_n647), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n618), .A2(new_n647), .A3(new_n569), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n636), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n569), .B1(new_n610), .B2(new_n616), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n656), .A2(new_n643), .A3(new_n642), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n657), .A2(new_n641), .A3(new_n636), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n634), .B1(new_n655), .B2(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(G120gat), .B(G148gat), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT105), .ZN(new_n662));
  XNOR2_X1  g461(.A(G176gat), .B(G204gat), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n662), .B(new_n663), .Z(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n634), .B(new_n664), .C1(new_n655), .C2(new_n659), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n474), .A2(new_n554), .A3(new_n633), .A4(new_n668), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n340), .A2(KEYINPUT107), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n340), .A2(KEYINPUT107), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n673), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g473(.A1(new_n669), .A2(new_n418), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT16), .B(G8gat), .Z(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(new_n486), .B2(new_n675), .ZN(new_n678));
  MUX2_X1   g477(.A(new_n677), .B(new_n678), .S(KEYINPUT42), .Z(G1325gat));
  AND2_X1   g478(.A1(new_n432), .A2(new_n433), .ZN(new_n680));
  OAI21_X1  g479(.A(G15gat), .B1(new_n669), .B2(new_n680), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n413), .A2(G15gat), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n681), .B1(new_n669), .B2(new_n682), .ZN(G1326gat));
  NAND3_X1  g482(.A1(new_n474), .A2(new_n438), .A3(new_n554), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n633), .A2(new_n668), .ZN(new_n685));
  OR3_X1    g484(.A1(new_n684), .A2(KEYINPUT108), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT108), .B1(new_n684), .B2(new_n685), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n688), .B(new_n690), .ZN(G1327gat));
  INV_X1    g490(.A(new_n668), .ZN(new_n692));
  INV_X1    g491(.A(new_n587), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n554), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n417), .A2(new_n426), .B1(new_n470), .B2(new_n472), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n632), .B(new_n700), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n701), .A2(KEYINPUT44), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n632), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT44), .B1(new_n699), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n698), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G29gat), .B1(new_n707), .B2(new_n672), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT45), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n699), .A2(new_n704), .A3(new_n698), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n672), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n517), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n709), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n710), .A2(KEYINPUT45), .A3(new_n517), .A4(new_n712), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n708), .A2(new_n714), .A3(new_n715), .ZN(G1328gat));
  OAI21_X1  g515(.A(G36gat), .B1(new_n707), .B2(new_n418), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n277), .A2(new_n518), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT46), .B1(new_n711), .B2(new_n718), .ZN(new_n719));
  OR3_X1    g518(.A1(new_n711), .A2(KEYINPUT46), .A3(new_n718), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n717), .A2(new_n719), .A3(new_n720), .ZN(G1329gat));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n722), .B1(new_n474), .B2(new_n632), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n699), .A2(new_n702), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n434), .B(new_n697), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(G43gat), .ZN(new_n726));
  INV_X1    g525(.A(new_n413), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n710), .A2(new_n499), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1330gat));
  AOI21_X1  g530(.A(new_n511), .B1(new_n706), .B2(new_n438), .ZN(new_n732));
  NOR4_X1   g531(.A1(new_n684), .A2(G50gat), .A3(new_n704), .A4(new_n695), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT48), .ZN(new_n734));
  OR3_X1    g533(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n732), .B2(new_n733), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(G1331gat));
  NOR4_X1   g536(.A1(new_n668), .A2(new_n587), .A3(new_n554), .A4(new_n632), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n474), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n672), .ZN(new_n740));
  XOR2_X1   g539(.A(KEYINPUT110), .B(G57gat), .Z(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1332gat));
  AND2_X1   g541(.A1(new_n474), .A2(new_n738), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n418), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT111), .ZN(new_n746));
  OR2_X1    g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1333gat));
  NAND3_X1  g547(.A1(new_n743), .A2(new_n556), .A3(new_n727), .ZN(new_n749));
  OAI21_X1  g548(.A(G71gat), .B1(new_n739), .B2(new_n680), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g550(.A(new_n751), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g551(.A1(new_n380), .A2(new_n414), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n739), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(new_n557), .ZN(G1335gat));
  NOR3_X1   g554(.A1(new_n693), .A2(new_n554), .A3(new_n668), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n723), .B2(new_n724), .ZN(new_n757));
  INV_X1    g556(.A(G85gat), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n757), .A2(new_n758), .A3(new_n672), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n454), .A2(new_n277), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n753), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n456), .A2(new_n468), .A3(new_n464), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n423), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n680), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n753), .B1(new_n341), .B2(new_n347), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI22_X1  g565(.A1(new_n416), .A2(KEYINPUT35), .B1(new_n425), .B2(new_n415), .ZN(new_n767));
  OAI211_X1 g566(.A(KEYINPUT112), .B(new_n632), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n693), .A2(new_n554), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT112), .B1(new_n474), .B2(new_n632), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT51), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n699), .B2(new_n704), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n774), .A2(new_n775), .A3(new_n769), .A4(new_n768), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n772), .A2(new_n692), .A3(new_n776), .A4(new_n712), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n759), .B1(new_n777), .B2(new_n758), .ZN(G1336gat));
  NOR2_X1   g577(.A1(new_n418), .A2(G92gat), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n772), .A2(new_n692), .A3(new_n776), .A4(new_n779), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n277), .B(new_n756), .C1(new_n723), .C2(new_n724), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G92gat), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n784), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n780), .B(new_n782), .C1(new_n785), .C2(new_n784), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(G1337gat));
  INV_X1    g588(.A(G99gat), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n757), .A2(new_n790), .A3(new_n680), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n772), .A2(new_n727), .A3(new_n776), .A4(new_n692), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n791), .B1(new_n792), .B2(new_n790), .ZN(G1338gat));
  NOR2_X1   g592(.A1(new_n753), .A2(G106gat), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n772), .A2(new_n692), .A3(new_n776), .A4(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(G106gat), .B1(new_n757), .B2(new_n753), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XOR2_X1   g596(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n798), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n795), .A2(new_n800), .A3(new_n796), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(G1339gat));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n653), .A2(new_n635), .ZN(new_n804));
  AOI211_X1 g603(.A(KEYINPUT104), .B(KEYINPUT10), .C1(new_n657), .C2(new_n641), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n650), .B1(new_n646), .B2(new_n647), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT54), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n655), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n654), .B1(new_n805), .B2(new_n806), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(new_n811), .A3(new_n635), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n665), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n803), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n655), .A2(new_n659), .A3(new_n665), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n653), .B1(new_n649), .B2(new_n651), .ZN(new_n817));
  OAI211_X1 g616(.A(KEYINPUT54), .B(new_n807), .C1(new_n817), .C2(new_n636), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n818), .A2(KEYINPUT55), .A3(new_n665), .A4(new_n812), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n814), .A2(new_n554), .A3(new_n816), .A4(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n552), .A2(new_n551), .ZN(new_n821));
  OAI22_X1  g620(.A1(new_n542), .A2(new_n543), .B1(new_n530), .B2(new_n529), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n821), .A2(new_n479), .B1(new_n478), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n666), .A2(new_n823), .A3(new_n667), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n701), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n814), .A2(new_n823), .A3(new_n816), .A4(new_n819), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n701), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n587), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n633), .A2(new_n696), .A3(new_n668), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT115), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n753), .A2(new_n727), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n672), .A2(new_n833), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n832), .A2(KEYINPUT116), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT116), .B1(new_n832), .B2(new_n834), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n835), .A2(new_n836), .A3(new_n277), .ZN(new_n837));
  AOI21_X1  g636(.A(G113gat), .B1(new_n837), .B2(new_n554), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n832), .A2(new_n834), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n839), .A2(new_n277), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n554), .A2(G113gat), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(G1340gat));
  AOI21_X1  g641(.A(G120gat), .B1(new_n837), .B2(new_n692), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n668), .A2(new_n313), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n843), .B1(new_n840), .B2(new_n844), .ZN(G1341gat));
  NAND3_X1  g644(.A1(new_n837), .A2(new_n574), .A3(new_n693), .ZN(new_n846));
  INV_X1    g645(.A(new_n840), .ZN(new_n847));
  OAI21_X1  g646(.A(G127gat), .B1(new_n847), .B2(new_n587), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(G1342gat));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n277), .A2(new_n704), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(G134gat), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n835), .A2(new_n836), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT56), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(G134gat), .B1(new_n839), .B2(new_n852), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n855), .B2(new_n856), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n850), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n855), .A2(new_n856), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n862), .A2(new_n857), .A3(KEYINPUT117), .A4(new_n859), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(G1343gat));
  NOR2_X1   g663(.A1(new_n672), .A2(new_n434), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n418), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n753), .B1(new_n829), .B2(new_n831), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n867), .A2(KEYINPUT57), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n820), .A2(KEYINPUT118), .A3(new_n824), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n632), .B1(new_n825), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n828), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n831), .B1(new_n872), .B2(new_n693), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n438), .A2(KEYINPUT57), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n866), .B1(new_n868), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n554), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n296), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n867), .A2(new_n865), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n696), .A2(G141gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n880), .A2(new_n418), .A3(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(KEYINPUT58), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n878), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n295), .B1(new_n876), .B2(new_n554), .ZN(new_n887));
  INV_X1    g686(.A(new_n882), .ZN(new_n888));
  OAI211_X1 g687(.A(KEYINPUT58), .B(new_n884), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n886), .A2(new_n889), .ZN(G1344gat));
  NOR2_X1   g689(.A1(new_n827), .A2(new_n704), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n891), .B1(new_n871), .B2(new_n869), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n587), .B1(new_n892), .B2(KEYINPUT120), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n894));
  AOI211_X1 g693(.A(new_n894), .B(new_n891), .C1(new_n871), .C2(new_n869), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n830), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT57), .B1(new_n896), .B2(new_n438), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n832), .A2(new_n874), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n865), .A2(new_n418), .A3(new_n692), .ZN(new_n900));
  OAI211_X1 g699(.A(KEYINPUT59), .B(G148gat), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n879), .A2(new_n277), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n292), .A3(new_n692), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n292), .B1(new_n876), .B2(new_n692), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n901), .B(new_n903), .C1(KEYINPUT59), .C2(new_n904), .ZN(G1345gat));
  NAND3_X1  g704(.A1(new_n902), .A2(new_n284), .A3(new_n693), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n876), .A2(new_n693), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(new_n284), .ZN(G1346gat));
  NAND3_X1  g707(.A1(new_n880), .A2(new_n285), .A3(new_n851), .ZN(new_n909));
  AOI211_X1 g708(.A(new_n701), .B(new_n866), .C1(new_n868), .C2(new_n875), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n285), .ZN(G1347gat));
  NOR2_X1   g710(.A1(new_n833), .A2(new_n418), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(KEYINPUT121), .Z(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n672), .A3(new_n832), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(G169gat), .B1(new_n915), .B2(new_n554), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n832), .A2(new_n672), .A3(new_n912), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n917), .B(new_n918), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n696), .A2(new_n205), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(G1348gat));
  NAND3_X1  g720(.A1(new_n915), .A2(new_n206), .A3(new_n692), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n919), .A2(new_n692), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(new_n206), .ZN(G1349gat));
  NOR2_X1   g723(.A1(new_n587), .A2(new_n223), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n913), .A2(new_n672), .A3(new_n832), .A4(new_n925), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT123), .Z(new_n927));
  INV_X1    g726(.A(KEYINPUT60), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n917), .A2(KEYINPUT122), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n917), .A2(KEYINPUT122), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n929), .A2(new_n930), .A3(new_n587), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n927), .B(new_n928), .C1(new_n209), .C2(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n209), .B1(new_n919), .B2(new_n693), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n926), .B(KEYINPUT123), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT60), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n932), .A2(new_n935), .ZN(G1350gat));
  OR3_X1    g735(.A1(new_n914), .A2(G190gat), .A3(new_n701), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT61), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n919), .A2(new_n632), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(G190gat), .ZN(new_n940));
  AOI211_X1 g739(.A(KEYINPUT61), .B(new_n210), .C1(new_n919), .C2(new_n632), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(G1351gat));
  NOR2_X1   g741(.A1(new_n434), .A2(new_n418), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n944), .A2(new_n753), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n832), .A2(new_n672), .A3(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n554), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n899), .A2(new_n712), .A3(new_n944), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n554), .A2(G197gat), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(G1352gat));
  XOR2_X1   g750(.A(KEYINPUT124), .B(G204gat), .Z(new_n952));
  AND2_X1   g751(.A1(new_n692), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n832), .A2(new_n672), .A3(new_n945), .A4(new_n953), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n954), .A2(KEYINPUT125), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(KEYINPUT125), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT62), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n944), .A2(new_n712), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n692), .B(new_n959), .C1(new_n897), .C2(new_n898), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n958), .B1(new_n961), .B2(new_n952), .ZN(G1353gat));
  NAND3_X1  g761(.A1(new_n947), .A2(new_n245), .A3(new_n693), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n693), .B(new_n959), .C1(new_n897), .C2(new_n898), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT63), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n245), .B1(KEYINPUT126), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n965), .A2(KEYINPUT126), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n967), .B1(new_n964), .B2(new_n966), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n963), .B1(new_n968), .B2(new_n969), .ZN(G1354gat));
  NAND2_X1  g769(.A1(new_n632), .A2(G218gat), .ZN(new_n971));
  XOR2_X1   g770(.A(new_n971), .B(KEYINPUT127), .Z(new_n972));
  OR2_X1    g771(.A1(new_n946), .A2(new_n701), .ZN(new_n973));
  AOI22_X1  g772(.A1(new_n949), .A2(new_n972), .B1(new_n246), .B2(new_n973), .ZN(G1355gat));
endmodule


