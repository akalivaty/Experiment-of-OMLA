//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT0), .B(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(G143), .B(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  INV_X1    g012(.A(G137), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(G134), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT11), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(G134), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n200), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OAI211_X1 g021(.A(G134), .B(new_n199), .C1(new_n203), .C2(KEYINPUT11), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n198), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n200), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT64), .B(KEYINPUT11), .ZN(new_n211));
  INV_X1    g025(.A(new_n206), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n208), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G131), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n197), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT2), .A2(G113), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT68), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n216), .B(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(KEYINPUT2), .A2(G113), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT67), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n221), .B1(KEYINPUT2), .B2(G113), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  AND2_X1   g038(.A1(KEYINPUT69), .A2(G119), .ZN(new_n225));
  NOR2_X1   g039(.A1(KEYINPUT69), .A2(G119), .ZN(new_n226));
  OAI21_X1  g040(.A(G116), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G116), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G119), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n218), .A2(new_n223), .A3(new_n227), .A4(new_n229), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G128), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n187), .A3(G143), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n189), .B(G146), .C1(new_n234), .C2(KEYINPUT1), .ZN(new_n236));
  OR2_X1    g050(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n235), .B(new_n236), .C1(new_n191), .C2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(G131), .B1(new_n212), .B2(new_n200), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n238), .B(new_n239), .C1(new_n213), .C2(G131), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n215), .A2(new_n233), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT28), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n215), .A2(new_n233), .A3(KEYINPUT28), .A4(new_n240), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n231), .A2(new_n232), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n213), .A2(G131), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n205), .A2(new_n206), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n247), .A2(new_n198), .A3(new_n208), .A4(new_n210), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n246), .A2(new_n248), .B1(new_n193), .B2(new_n196), .ZN(new_n249));
  INV_X1    g063(.A(new_n240), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n245), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n243), .A2(new_n244), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT72), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n254), .B(G101), .ZN(new_n255));
  INV_X1    g069(.A(G237), .ZN(new_n256));
  INV_X1    g070(.A(G953), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n257), .A3(G210), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n255), .B(new_n258), .ZN(new_n259));
  NOR3_X1   g073(.A1(new_n249), .A2(new_n250), .A3(new_n245), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n233), .B1(new_n215), .B2(new_n240), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT28), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n253), .A2(new_n259), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT29), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n259), .B(KEYINPUT70), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(KEYINPUT29), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n215), .A2(KEYINPUT65), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n249), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n240), .A2(KEYINPUT66), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT66), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n248), .A2(new_n273), .A3(new_n238), .A4(new_n239), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n269), .A2(new_n271), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n245), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n243), .A2(new_n244), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n268), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n259), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT30), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n249), .A2(new_n250), .A3(new_n281), .ZN(new_n282));
  AOI211_X1 g096(.A(new_n233), .B(new_n282), .C1(new_n276), .C2(new_n281), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n280), .B1(new_n283), .B2(new_n260), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n266), .A2(G472), .A3(new_n279), .A4(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(G472), .A2(G902), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT73), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT32), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n278), .A2(new_n277), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n267), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n276), .A2(new_n281), .ZN(new_n293));
  INV_X1    g107(.A(new_n282), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n245), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n259), .A3(new_n241), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT31), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n282), .B1(new_n276), .B2(new_n281), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n260), .B1(new_n299), .B2(new_n245), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(KEYINPUT31), .A3(new_n259), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n292), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(G472), .A2(G902), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(KEYINPUT71), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n289), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  NOR4_X1   g119(.A1(new_n283), .A2(new_n297), .A3(new_n280), .A4(new_n260), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT31), .B1(new_n300), .B2(new_n259), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n291), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n304), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(KEYINPUT32), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT73), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n285), .A2(new_n311), .A3(new_n286), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n288), .A2(new_n305), .A3(new_n310), .A4(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT74), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n302), .A2(new_n289), .A3(new_n304), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT32), .B1(new_n308), .B2(new_n309), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n285), .A2(new_n311), .A3(new_n286), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n311), .B1(new_n285), .B2(new_n286), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n318), .A2(new_n321), .A3(KEYINPUT74), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n315), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G125), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(KEYINPUT16), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n324), .A2(KEYINPUT76), .A3(G125), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n330));
  XNOR2_X1  g144(.A(G125), .B(G140), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT16), .ZN(new_n333));
  OAI211_X1 g147(.A(G146), .B(new_n327), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G125), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G140), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n325), .A2(new_n336), .A3(new_n330), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n333), .B1(new_n337), .B2(new_n328), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n187), .B1(new_n338), .B2(new_n326), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n334), .A2(new_n339), .A3(KEYINPUT77), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n341), .B(new_n187), .C1(new_n338), .C2(new_n326), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n256), .A2(new_n257), .A3(G214), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(new_n189), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(KEYINPUT17), .A3(G131), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT91), .ZN(new_n348));
  INV_X1    g162(.A(new_n345), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n198), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n345), .A2(G131), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n352), .A2(KEYINPUT17), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT91), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n343), .A2(new_n355), .A3(new_n346), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n348), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(G113), .B(G122), .ZN(new_n358));
  INV_X1    g172(.A(G104), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n358), .B(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT18), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(new_n198), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n349), .B(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n331), .A2(new_n187), .ZN(new_n364));
  INV_X1    g178(.A(new_n332), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n364), .B1(new_n365), .B2(new_n187), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n357), .A2(new_n360), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT19), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n331), .A2(KEYINPUT90), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT90), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n332), .B1(new_n371), .B2(new_n331), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n370), .B1(new_n372), .B2(new_n369), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n352), .B(new_n334), .C1(new_n373), .C2(G146), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n367), .ZN(new_n375));
  INV_X1    g189(.A(new_n360), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n368), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(G475), .A2(G902), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT20), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT20), .ZN(new_n381));
  INV_X1    g195(.A(new_n379), .ZN(new_n382));
  AOI211_X1 g196(.A(new_n381), .B(new_n382), .C1(new_n368), .C2(new_n377), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n355), .B1(new_n343), .B2(new_n346), .ZN(new_n385));
  INV_X1    g199(.A(new_n346), .ZN(new_n386));
  AOI211_X1 g200(.A(KEYINPUT91), .B(new_n386), .C1(new_n340), .C2(new_n342), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n385), .A2(new_n387), .A3(new_n353), .ZN(new_n388));
  INV_X1    g202(.A(new_n367), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n376), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n368), .ZN(new_n391));
  INV_X1    g205(.A(G902), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G475), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n384), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT14), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT92), .ZN(new_n397));
  INV_X1    g211(.A(G122), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n397), .B1(new_n398), .B2(G116), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n228), .A2(KEYINPUT92), .A3(G122), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n396), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT95), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n228), .A2(G122), .ZN(new_n403));
  OR3_X1    g217(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n399), .A2(new_n396), .A3(new_n400), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n402), .B1(new_n401), .B2(new_n403), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G107), .ZN(new_n408));
  XNOR2_X1  g222(.A(G128), .B(G143), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(KEYINPUT93), .ZN(new_n410));
  INV_X1    g224(.A(G134), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n410), .B(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n403), .B1(new_n399), .B2(new_n400), .ZN(new_n413));
  INV_X1    g227(.A(G107), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  XOR2_X1   g229(.A(new_n415), .B(KEYINPUT94), .Z(new_n416));
  NAND3_X1  g230(.A1(new_n408), .A2(new_n412), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n410), .A2(new_n411), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n409), .A2(KEYINPUT13), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n189), .A2(G128), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n419), .B(G134), .C1(KEYINPUT13), .C2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n413), .A2(new_n414), .ZN(new_n422));
  INV_X1    g236(.A(new_n415), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n418), .B(new_n421), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n417), .A2(new_n424), .ZN(new_n425));
  XOR2_X1   g239(.A(KEYINPUT9), .B(G234), .Z(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(G217), .A3(new_n257), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT96), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT97), .ZN(new_n430));
  INV_X1    g244(.A(new_n428), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n417), .A2(new_n431), .A3(new_n424), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n417), .A2(KEYINPUT97), .A3(new_n431), .A4(new_n424), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n392), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G478), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(KEYINPUT15), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n435), .B(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n395), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n335), .B1(new_n193), .B2(new_n196), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n440), .B1(new_n335), .B2(new_n238), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT88), .ZN(new_n442));
  INV_X1    g256(.A(G224), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(G953), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n441), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n444), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT7), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n445), .B(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n227), .A2(KEYINPUT5), .A3(new_n229), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT69), .B(G119), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT5), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(new_n451), .A3(G116), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(G113), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n232), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT3), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n455), .B1(new_n359), .B2(G107), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n414), .A2(KEYINPUT3), .A3(G104), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G101), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n458), .B(new_n459), .C1(G104), .C2(new_n414), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT84), .B1(new_n414), .B2(G104), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT84), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n359), .A3(G107), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n461), .B(new_n463), .C1(new_n359), .C2(G107), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G101), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n454), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT86), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n460), .A2(new_n465), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(new_n232), .A3(new_n453), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT86), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n454), .A2(new_n471), .A3(new_n466), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n468), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT87), .ZN(new_n474));
  XOR2_X1   g288(.A(G110), .B(G122), .Z(new_n475));
  XOR2_X1   g289(.A(new_n475), .B(KEYINPUT8), .Z(new_n476));
  AND3_X1   g290(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n474), .B1(new_n473), .B2(new_n476), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n448), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT89), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n458), .B1(G104), .B2(new_n414), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G101), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(KEYINPUT4), .A3(new_n460), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT4), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(new_n484), .A3(G101), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n245), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n475), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n487), .A3(new_n470), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT89), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n448), .B(new_n489), .C1(new_n477), .C2(new_n478), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n480), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n486), .A2(new_n470), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n475), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(KEYINPUT6), .A3(new_n488), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n441), .B(new_n444), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n492), .A2(new_n496), .A3(new_n475), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n491), .A2(new_n392), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G210), .B1(G237), .B2(G902), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n491), .A2(new_n392), .A3(new_n500), .A4(new_n498), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(G234), .A2(G237), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n505), .A2(G952), .A3(new_n257), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  XOR2_X1   g321(.A(KEYINPUT21), .B(G898), .Z(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n505), .A2(G902), .A3(G953), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n507), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(G214), .B1(G237), .B2(G902), .ZN(new_n514));
  AND4_X1   g328(.A1(new_n439), .A2(new_n504), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n257), .A2(G221), .A3(G234), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(KEYINPUT22), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(G137), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT23), .ZN(new_n519));
  OAI21_X1  g333(.A(G128), .B1(new_n225), .B2(new_n226), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n234), .A2(G119), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n225), .A2(new_n226), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT23), .B1(new_n523), .B2(new_n234), .ZN(new_n524));
  XOR2_X1   g338(.A(KEYINPUT78), .B(G110), .Z(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n522), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n521), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(new_n450), .B2(G128), .ZN(new_n529));
  XOR2_X1   g343(.A(KEYINPUT24), .B(G110), .Z(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT79), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n519), .B1(new_n450), .B2(G128), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n533), .B(new_n525), .C1(new_n529), .C2(new_n519), .ZN(new_n534));
  OR2_X1    g348(.A1(new_n529), .A2(new_n530), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT79), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n532), .A2(new_n364), .A3(new_n334), .A4(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(KEYINPUT75), .B1(new_n522), .B2(new_n524), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT75), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n540), .B(new_n533), .C1(new_n529), .C2(new_n519), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n541), .A3(G110), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n529), .A2(new_n530), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n340), .A2(new_n542), .A3(new_n342), .A4(new_n543), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n538), .A2(KEYINPUT80), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT80), .B1(new_n538), .B2(new_n544), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n518), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n518), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n538), .A2(new_n544), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT80), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n547), .A2(new_n392), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n555));
  INV_X1    g369(.A(new_n553), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n547), .A2(new_n392), .A3(new_n551), .A4(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(G217), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n559), .B1(G234), .B2(new_n392), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n558), .A2(KEYINPUT82), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT82), .B1(new_n558), .B2(new_n560), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n560), .A2(G902), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n547), .A2(new_n551), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n209), .A2(new_n214), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n469), .A2(new_n238), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n460), .A2(new_n465), .A3(new_n238), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n569), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT12), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n569), .B(KEYINPUT12), .C1(new_n570), .C2(new_n572), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(G110), .B(G140), .ZN(new_n578));
  INV_X1    g392(.A(G227), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(G953), .ZN(new_n580));
  XOR2_X1   g394(.A(new_n578), .B(new_n580), .Z(new_n581));
  NAND3_X1  g395(.A1(new_n483), .A2(new_n197), .A3(new_n485), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n469), .A2(KEYINPUT10), .A3(new_n238), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT10), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n571), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n582), .A2(new_n583), .A3(new_n568), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT85), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n586), .A2(KEYINPUT85), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n577), .B(new_n581), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n586), .A2(KEYINPUT85), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n591), .A2(new_n587), .B1(new_n569), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n590), .B1(new_n593), .B2(new_n581), .ZN(new_n594));
  INV_X1    g408(.A(G469), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(new_n392), .ZN(new_n596));
  NAND2_X1  g410(.A1(G469), .A2(G902), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n592), .A2(new_n569), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n598), .B(new_n581), .C1(new_n588), .C2(new_n589), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n591), .A2(new_n587), .B1(new_n576), .B2(new_n575), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n581), .B(KEYINPUT83), .Z(new_n601));
  OAI211_X1 g415(.A(new_n599), .B(G469), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n596), .A2(new_n597), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(G221), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n426), .B2(new_n392), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n323), .A2(new_n515), .A3(new_n567), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT98), .B(G101), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G3));
  INV_X1    g425(.A(KEYINPUT99), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n504), .B2(new_n514), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n384), .A2(new_n394), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n433), .A2(new_n616), .A3(new_n434), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n429), .A2(KEYINPUT33), .A3(new_n432), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n436), .A2(G902), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT100), .B(G478), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n435), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n615), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n504), .A2(new_n612), .A3(new_n514), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n614), .A2(new_n513), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(G472), .B1(new_n302), .B2(G902), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n308), .A2(new_n309), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n563), .A2(new_n631), .A3(new_n565), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n608), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT34), .B(G104), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT101), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n634), .B(new_n636), .ZN(G6));
  INV_X1    g451(.A(new_n514), .ZN(new_n638));
  AOI211_X1 g452(.A(KEYINPUT99), .B(new_n638), .C1(new_n502), .C2(new_n503), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n613), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n615), .A2(new_n438), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n640), .A2(new_n513), .A3(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n633), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT35), .B(G107), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  NOR2_X1   g460(.A1(new_n548), .A2(KEYINPUT36), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT102), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(new_n549), .Z(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n564), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n607), .B1(new_n563), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n515), .A2(new_n631), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G110), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  INV_X1    g469(.A(G900), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n511), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n506), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n641), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n640), .A2(new_n323), .A3(new_n651), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G128), .ZN(G30));
  XOR2_X1   g476(.A(new_n658), .B(KEYINPUT104), .Z(new_n663));
  XOR2_X1   g477(.A(new_n663), .B(KEYINPUT39), .Z(new_n664));
  OR3_X1    g478(.A1(new_n607), .A2(KEYINPUT40), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n558), .A2(new_n560), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT82), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n558), .A2(KEYINPUT82), .A3(new_n560), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n668), .A2(new_n669), .A3(new_n650), .ZN(new_n670));
  INV_X1    g484(.A(new_n438), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n615), .A2(new_n671), .ZN(new_n672));
  AND4_X1   g486(.A1(new_n514), .A2(new_n665), .A3(new_n670), .A4(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n251), .A2(new_n241), .ZN(new_n674));
  AOI22_X1  g488(.A1(new_n300), .A2(new_n259), .B1(new_n267), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(G472), .B1(new_n675), .B2(G902), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n318), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n504), .B(KEYINPUT38), .ZN(new_n678));
  INV_X1    g492(.A(new_n664), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n608), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n673), .A2(new_n677), .A3(new_n678), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  AND3_X1   g497(.A1(new_n395), .A2(new_n623), .A3(new_n658), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n640), .A2(new_n323), .A3(new_n651), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  NOR3_X1   g500(.A1(new_n613), .A2(new_n639), .A3(new_n512), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n566), .B1(new_n315), .B2(new_n322), .ZN(new_n688));
  INV_X1    g502(.A(new_n596), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n595), .B1(new_n594), .B2(new_n392), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n605), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n687), .A2(new_n688), .A3(new_n625), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT41), .B(G113), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G15));
  NAND4_X1  g510(.A1(new_n687), .A2(new_n688), .A3(new_n642), .A4(new_n693), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G116), .ZN(G18));
  AOI21_X1  g512(.A(new_n670), .B1(new_n315), .B2(new_n322), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n687), .A2(new_n699), .A3(new_n439), .A4(new_n693), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G119), .ZN(G21));
  NAND2_X1  g515(.A1(new_n253), .A2(new_n264), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n298), .A2(new_n301), .B1(new_n267), .B2(new_n702), .ZN(new_n703));
  OR2_X1    g517(.A1(new_n703), .A2(new_n304), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n704), .A2(new_n628), .ZN(new_n705));
  AND4_X1   g519(.A1(new_n513), .A2(new_n563), .A3(new_n705), .A4(new_n565), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n640), .A2(new_n706), .A3(new_n672), .A4(new_n693), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G122), .ZN(G24));
  NAND3_X1  g522(.A1(new_n668), .A2(new_n669), .A3(new_n650), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n684), .A2(new_n709), .A3(new_n705), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n640), .A2(new_n710), .A3(new_n693), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G125), .ZN(G27));
  NAND3_X1  g526(.A1(new_n502), .A2(new_n514), .A3(new_n503), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n603), .A2(KEYINPUT105), .A3(new_n606), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT105), .B1(new_n603), .B2(new_n606), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n323), .A2(new_n567), .A3(new_n684), .A4(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT106), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT42), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n688), .A2(KEYINPUT106), .A3(new_n684), .A4(new_n716), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n310), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n724), .B1(new_n310), .B2(new_n723), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n317), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(KEYINPUT108), .B1(new_n316), .B2(KEYINPUT107), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n310), .A2(new_n723), .A3(new_n724), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n305), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n727), .A2(new_n321), .A3(new_n730), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n731), .A2(new_n567), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(KEYINPUT42), .A3(new_n684), .A4(new_n716), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n722), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G131), .ZN(G33));
  AND3_X1   g549(.A1(new_n688), .A2(new_n660), .A3(new_n716), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n411), .ZN(G36));
  AND2_X1   g551(.A1(new_n368), .A2(new_n377), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n381), .B1(new_n738), .B2(new_n382), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n378), .A2(KEYINPUT20), .A3(new_n379), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n394), .A2(new_n623), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(KEYINPUT109), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n384), .A2(new_n394), .A3(new_n623), .A4(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n709), .A2(new_n630), .A3(new_n744), .A4(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n748));
  OAI21_X1  g562(.A(KEYINPUT110), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n744), .A2(new_n746), .A3(new_n630), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n750), .A2(new_n751), .A3(KEYINPUT44), .A4(new_n709), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n502), .A2(new_n514), .A3(new_n503), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n749), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT111), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n749), .A2(new_n752), .A3(new_n756), .A4(new_n753), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n747), .A2(new_n748), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT112), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n747), .A2(new_n760), .A3(new_n748), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n755), .A2(new_n757), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n599), .B(KEYINPUT45), .C1(new_n600), .C2(new_n601), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(G469), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n597), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT46), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n689), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n770), .A2(KEYINPUT46), .A3(new_n597), .ZN(new_n774));
  AOI211_X1 g588(.A(new_n605), .B(new_n664), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n755), .A2(KEYINPUT113), .A3(new_n757), .A4(new_n762), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n765), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G137), .ZN(G39));
  AOI21_X1  g592(.A(new_n605), .B1(new_n773), .B2(new_n774), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT47), .Z(new_n780));
  NOR4_X1   g594(.A1(new_n780), .A2(new_n615), .A3(new_n624), .A4(new_n659), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n323), .A2(new_n567), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(new_n753), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  NOR2_X1   g598(.A1(new_n678), .A2(new_n638), .ZN(new_n785));
  INV_X1    g599(.A(new_n677), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT49), .ZN(new_n787));
  AOI211_X1 g601(.A(new_n605), .B(new_n741), .C1(new_n691), .C2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n566), .B1(new_n692), .B2(KEYINPUT49), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n785), .A2(new_n786), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n780), .B1(new_n606), .B2(new_n692), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n744), .A2(new_n746), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n507), .A2(new_n567), .A3(new_n794), .A4(new_n705), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n792), .A2(new_n753), .A3(new_n795), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n713), .A2(new_n692), .A3(new_n506), .A4(new_n605), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n797), .A2(new_n567), .A3(new_n786), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(new_n615), .A3(new_n624), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n797), .A2(new_n794), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n709), .A2(new_n705), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n796), .A2(new_n799), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n678), .A2(new_n514), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n795), .A2(new_n693), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT50), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n791), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(G952), .A3(new_n257), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n803), .A2(new_n791), .A3(new_n806), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n661), .A2(new_n685), .A3(new_n711), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n670), .A2(new_n813), .A3(new_n658), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT116), .B1(new_n709), .B2(new_n659), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n814), .A2(new_n608), .A3(new_n815), .A4(new_n677), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n640), .A2(new_n672), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT52), .B1(new_n812), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n323), .A2(new_n567), .A3(new_n693), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n323), .A2(new_n439), .A3(new_n709), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n614), .A2(new_n513), .A3(new_n626), .A4(new_n693), .ZN(new_n822));
  OAI22_X1  g636(.A1(new_n643), .A2(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n614), .A2(new_n626), .A3(new_n672), .A4(new_n693), .ZN(new_n824));
  INV_X1    g638(.A(new_n706), .ZN(new_n825));
  OAI22_X1  g639(.A1(new_n820), .A2(new_n627), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n613), .A2(new_n639), .A3(new_n671), .A4(new_n615), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n709), .A2(new_n659), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n607), .B1(new_n829), .B2(new_n813), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n828), .A2(new_n677), .A3(new_n815), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n709), .A2(new_n608), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n832), .B1(new_n315), .B2(new_n322), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n833), .B(new_n640), .C1(new_n660), .C2(new_n684), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n831), .A2(new_n834), .A3(new_n835), .A4(new_n711), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n734), .A2(new_n819), .A3(new_n827), .A4(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n313), .A2(new_n314), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT74), .B1(new_n318), .B2(new_n321), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n651), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n671), .A2(new_n384), .A3(new_n394), .A4(new_n658), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n753), .A2(new_n843), .A3(KEYINPUT114), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n845), .B1(new_n713), .B2(new_n842), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n838), .B1(new_n841), .B2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n833), .A2(KEYINPUT115), .A3(new_n846), .A4(new_n844), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n736), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n504), .A2(new_n514), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(new_n512), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n641), .B1(new_n615), .B2(new_n624), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n632), .A2(new_n852), .A3(new_n853), .A4(new_n608), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n801), .A2(new_n716), .A3(new_n684), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n609), .A2(new_n854), .A3(new_n652), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n850), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n811), .B1(new_n837), .B2(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n819), .A2(new_n836), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n694), .A2(new_n697), .A3(new_n700), .A4(new_n707), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(new_n722), .B2(new_n733), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n850), .A2(new_n856), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n859), .A2(KEYINPUT53), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT54), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n795), .A2(new_n640), .A3(new_n693), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n734), .A2(new_n819), .A3(new_n827), .A4(new_n836), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n848), .A2(new_n849), .ZN(new_n868));
  INV_X1    g682(.A(new_n736), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n856), .A2(new_n868), .A3(KEYINPUT117), .A4(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n870), .A2(KEYINPUT53), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT117), .B1(new_n850), .B2(new_n856), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n867), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n874), .A2(new_n875), .A3(new_n858), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n810), .A2(new_n865), .A3(new_n866), .A4(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n798), .A2(new_n625), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n732), .A2(new_n800), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT48), .Z(new_n880));
  NOR3_X1   g694(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(G952), .A2(G953), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT118), .Z(new_n883));
  OAI21_X1  g697(.A(new_n790), .B1(new_n881), .B2(new_n883), .ZN(G75));
  AOI21_X1  g698(.A(new_n392), .B1(new_n874), .B2(new_n858), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT56), .B1(new_n885), .B2(G210), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n494), .A2(new_n497), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(new_n495), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT55), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n886), .A2(new_n889), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n257), .A2(G952), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(G51));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n894));
  AOI211_X1 g708(.A(new_n392), .B(new_n770), .C1(new_n874), .C2(new_n858), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n597), .B(KEYINPUT57), .Z(new_n896));
  AND3_X1   g710(.A1(new_n874), .A2(new_n875), .A3(new_n858), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n875), .B1(new_n874), .B2(new_n858), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n895), .B1(new_n899), .B2(new_n594), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n894), .B1(new_n900), .B2(new_n892), .ZN(new_n901));
  INV_X1    g715(.A(new_n892), .ZN(new_n902));
  INV_X1    g716(.A(new_n594), .ZN(new_n903));
  INV_X1    g717(.A(new_n858), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n870), .A2(KEYINPUT53), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n837), .A2(new_n905), .A3(new_n872), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT54), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n876), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n903), .B1(new_n908), .B2(new_n896), .ZN(new_n909));
  OAI211_X1 g723(.A(KEYINPUT119), .B(new_n902), .C1(new_n909), .C2(new_n895), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n901), .A2(new_n910), .ZN(G54));
  NAND3_X1  g725(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n912), .A2(new_n738), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n738), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n913), .A2(new_n914), .A3(new_n892), .ZN(G60));
  INV_X1    g729(.A(KEYINPUT120), .ZN(new_n916));
  NAND2_X1  g730(.A1(G478), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT59), .Z(new_n918));
  AOI21_X1  g732(.A(new_n918), .B1(new_n865), .B2(new_n876), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n617), .A2(new_n618), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n902), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n920), .ZN(new_n922));
  AOI211_X1 g736(.A(new_n922), .B(new_n918), .C1(new_n907), .C2(new_n876), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n916), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n865), .A2(new_n876), .ZN(new_n925));
  INV_X1    g739(.A(new_n918), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n922), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n908), .A2(new_n920), .A3(new_n926), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n928), .A2(KEYINPUT120), .A3(new_n902), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n924), .A2(new_n930), .ZN(G63));
  NAND2_X1  g745(.A1(new_n874), .A2(new_n858), .ZN(new_n932));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT60), .Z(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n547), .A2(new_n551), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n892), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(KEYINPUT61), .B1(new_n937), .B2(KEYINPUT121), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n932), .A2(new_n649), .A3(new_n934), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n937), .B(new_n939), .C1(KEYINPUT121), .C2(KEYINPUT61), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(G66));
  OAI21_X1  g757(.A(G953), .B1(new_n509), .B2(new_n443), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n609), .A2(new_n854), .A3(new_n652), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n860), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n944), .B1(new_n946), .B2(G953), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n887), .B1(G898), .B2(new_n257), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(G69));
  AND3_X1   g763(.A1(new_n661), .A2(new_n685), .A3(new_n711), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n731), .A2(new_n567), .A3(new_n775), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT124), .B1(new_n951), .B2(new_n828), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n731), .A2(new_n567), .A3(new_n775), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n953), .A2(new_n817), .A3(new_n954), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n869), .B(new_n950), .C1(new_n952), .C2(new_n955), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n722), .A2(new_n733), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n777), .A2(new_n958), .A3(new_n783), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n257), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n257), .A2(G900), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT125), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT125), .ZN(new_n964));
  AOI211_X1 g778(.A(new_n964), .B(new_n961), .C1(new_n959), .C2(new_n257), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n299), .B(new_n373), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(KEYINPUT122), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n688), .A2(new_n853), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n969), .A2(new_n680), .A3(new_n713), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n682), .A2(new_n834), .A3(new_n711), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT62), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n950), .A2(KEYINPUT62), .A3(new_n682), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n970), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n777), .A2(new_n783), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n968), .B1(new_n976), .B2(new_n257), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT123), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI211_X1 g793(.A(KEYINPUT123), .B(new_n968), .C1(new_n976), .C2(new_n257), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(G953), .B1(new_n579), .B2(new_n656), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n967), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n982), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n960), .A2(new_n962), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n964), .ZN(new_n986));
  INV_X1    g800(.A(new_n966), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n960), .A2(KEYINPUT125), .A3(new_n962), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n977), .B(new_n978), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n984), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n983), .A2(new_n991), .ZN(G72));
  XOR2_X1   g806(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT127), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(new_n286), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n864), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n284), .A2(new_n296), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n892), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n946), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n995), .B1(new_n976), .B2(new_n999), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n1000), .B(new_n259), .C1(new_n260), .C2(new_n283), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n995), .B1(new_n959), .B2(new_n999), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n1002), .A2(new_n280), .A3(new_n300), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n998), .A2(new_n1001), .A3(new_n1003), .ZN(G57));
endmodule


