

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n349, n350, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n368, n369, n370, n371,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759;

  AND2_X1 U367 ( .A1(n430), .A2(n429), .ZN(n361) );
  NOR2_X2 U368 ( .A1(n562), .A2(n581), .ZN(n706) );
  BUF_X1 U369 ( .A(G113), .Z(n424) );
  XNOR2_X2 U370 ( .A(n487), .B(n486), .ZN(n755) );
  XNOR2_X1 U371 ( .A(n455), .B(n420), .ZN(n716) );
  XNOR2_X1 U372 ( .A(n404), .B(n403), .ZN(n455) );
  INV_X2 U373 ( .A(G116), .ZN(n505) );
  NOR2_X2 U374 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X2 U375 ( .A(G902), .B(KEYINPUT15), .Z(n685) );
  NAND2_X2 U376 ( .A1(n468), .A2(n380), .ZN(n436) );
  XNOR2_X1 U377 ( .A(n373), .B(n354), .ZN(n345) );
  NAND2_X1 U378 ( .A1(n345), .A2(n355), .ZN(n371) );
  INV_X2 U379 ( .A(G113), .ZN(n506) );
  XNOR2_X1 U380 ( .A(n349), .B(n366), .ZN(n365) );
  NAND2_X1 U381 ( .A1(n368), .A2(n361), .ZN(n349) );
  AND2_X2 U382 ( .A1(n756), .A2(n485), .ZN(n483) );
  XNOR2_X2 U383 ( .A(n631), .B(KEYINPUT33), .ZN(n649) );
  NAND2_X2 U384 ( .A1(n350), .A2(n394), .ZN(n488) );
  AND2_X2 U385 ( .A1(n397), .A2(n479), .ZN(n350) );
  XNOR2_X1 U386 ( .A(G119), .B(G110), .ZN(n525) );
  XNOR2_X1 U387 ( .A(G140), .B(G137), .ZN(n576) );
  NAND2_X1 U388 ( .A1(n660), .A2(n636), .ZN(n662) );
  BUF_X1 U389 ( .A(G143), .Z(n700) );
  XOR2_X1 U390 ( .A(KEYINPUT66), .B(KEYINPUT60), .Z(n352) );
  INV_X2 U391 ( .A(G953), .ZN(n731) );
  XOR2_X1 U392 ( .A(n719), .B(n499), .Z(n353) );
  XOR2_X1 U393 ( .A(n384), .B(n715), .Z(n354) );
  AND2_X4 U394 ( .A1(n461), .A2(n436), .ZN(n724) );
  NAND2_X2 U395 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X2 U396 ( .A(G128), .B(G143), .ZN(n476) );
  XNOR2_X2 U397 ( .A(n478), .B(KEYINPUT73), .ZN(n477) );
  NAND2_X1 U398 ( .A1(n644), .A2(n435), .ZN(n487) );
  INV_X2 U399 ( .A(KEYINPUT64), .ZN(n478) );
  AND2_X2 U400 ( .A1(n411), .A2(n432), .ZN(n711) );
  NOR2_X2 U401 ( .A1(n642), .A2(n589), .ZN(n535) );
  XNOR2_X2 U402 ( .A(n629), .B(n514), .ZN(n642) );
  XNOR2_X2 U403 ( .A(n443), .B(n600), .ZN(n753) );
  XNOR2_X2 U404 ( .A(n571), .B(n570), .ZN(n582) );
  XOR2_X2 U405 ( .A(KEYINPUT38), .B(n613), .Z(n651) );
  INV_X2 U406 ( .A(n629), .ZN(n669) );
  AND2_X2 U407 ( .A1(n428), .A2(n427), .ZN(n598) );
  INV_X1 U408 ( .A(n727), .ZN(n355) );
  XOR2_X1 U409 ( .A(G125), .B(G146), .Z(n568) );
  NOR2_X1 U410 ( .A1(n663), .A2(n662), .ZN(n639) );
  XNOR2_X1 U411 ( .A(n410), .B(n472), .ZN(n718) );
  XNOR2_X1 U412 ( .A(n568), .B(n567), .ZN(n414) );
  INV_X1 U413 ( .A(KEYINPUT48), .ZN(n366) );
  NAND2_X1 U414 ( .A1(n395), .A2(n419), .ZN(n394) );
  XOR2_X1 U415 ( .A(KEYINPUT42), .B(n605), .Z(n759) );
  NOR2_X1 U416 ( .A1(n658), .A2(n364), .ZN(n677) );
  XNOR2_X1 U417 ( .A(n362), .B(KEYINPUT107), .ZN(n609) );
  XNOR2_X1 U418 ( .A(n358), .B(KEYINPUT95), .ZN(n672) );
  NAND2_X1 U419 ( .A1(n563), .A2(n706), .ZN(n362) );
  NAND2_X1 U420 ( .A1(n639), .A2(n669), .ZN(n358) );
  XNOR2_X1 U421 ( .A(n584), .B(n583), .ZN(n421) );
  XNOR2_X1 U422 ( .A(n409), .B(KEYINPUT1), .ZN(n663) );
  NOR2_X1 U423 ( .A1(n726), .A2(G902), .ZN(n446) );
  INV_X1 U424 ( .A(n412), .ZN(n403) );
  XNOR2_X1 U425 ( .A(n414), .B(n413), .ZN(n412) );
  XNOR2_X1 U426 ( .A(n376), .B(n569), .ZN(n413) );
  XOR2_X1 U427 ( .A(n566), .B(KEYINPUT16), .Z(n374) );
  INV_X1 U428 ( .A(n689), .ZN(n359) );
  NAND2_X1 U429 ( .A1(G214), .A2(n572), .ZN(n650) );
  XNOR2_X1 U430 ( .A(n568), .B(n441), .ZN(n741) );
  XOR2_X2 U431 ( .A(G110), .B(G104), .Z(n577) );
  XOR2_X1 U432 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n567) );
  XNOR2_X1 U433 ( .A(KEYINPUT22), .B(KEYINPUT67), .ZN(n626) );
  XOR2_X1 U434 ( .A(KEYINPUT85), .B(KEYINPUT72), .Z(n376) );
  INV_X2 U435 ( .A(G122), .ZN(n415) );
  NAND2_X1 U436 ( .A1(n461), .A2(n460), .ZN(n433) );
  XNOR2_X2 U437 ( .A(n463), .B(KEYINPUT70), .ZN(n461) );
  XNOR2_X1 U438 ( .A(n356), .B(n352), .ZN(G60) );
  NAND2_X1 U439 ( .A1(n357), .A2(n355), .ZN(n356) );
  XNOR2_X1 U440 ( .A(n720), .B(n353), .ZN(n357) );
  NOR2_X2 U441 ( .A1(n753), .A2(n759), .ZN(n608) );
  BUF_X2 U442 ( .A(n632), .Z(n640) );
  XNOR2_X1 U443 ( .A(n360), .B(n359), .ZN(G57) );
  NAND2_X1 U444 ( .A1(n416), .A2(n355), .ZN(n360) );
  NAND2_X1 U445 ( .A1(n365), .A2(n616), .ZN(n400) );
  XNOR2_X2 U446 ( .A(n513), .B(G472), .ZN(n629) );
  NAND2_X1 U447 ( .A1(n644), .A2(n643), .ZN(n425) );
  NOR2_X2 U448 ( .A1(n634), .A2(n628), .ZN(n644) );
  XNOR2_X2 U449 ( .A(n363), .B(n390), .ZN(n756) );
  NOR2_X2 U450 ( .A1(n634), .A2(n431), .ZN(n363) );
  INV_X1 U451 ( .A(n649), .ZN(n364) );
  XNOR2_X1 U452 ( .A(n608), .B(n369), .ZN(n368) );
  INV_X1 U453 ( .A(n607), .ZN(n369) );
  XNOR2_X1 U454 ( .A(n371), .B(n370), .ZN(G51) );
  INV_X1 U455 ( .A(KEYINPUT56), .ZN(n370) );
  NAND2_X1 U456 ( .A1(n724), .A2(G210), .ZN(n373) );
  NAND2_X1 U457 ( .A1(n598), .A2(n599), .ZN(n444) );
  XNOR2_X2 U458 ( .A(n444), .B(KEYINPUT39), .ZN(n614) );
  XNOR2_X2 U459 ( .A(n433), .B(n399), .ZN(n398) );
  NOR2_X1 U460 ( .A1(G953), .A2(G237), .ZN(n504) );
  XNOR2_X1 U461 ( .A(n445), .B(n533), .ZN(n439) );
  NOR2_X1 U462 ( .A1(n587), .A2(n375), .ZN(n429) );
  XOR2_X1 U463 ( .A(KEYINPUT5), .B(KEYINPUT68), .Z(n502) );
  XNOR2_X1 U464 ( .A(G137), .B(KEYINPUT94), .ZN(n501) );
  INV_X1 U465 ( .A(KEYINPUT45), .ZN(n493) );
  XOR2_X1 U466 ( .A(KEYINPUT30), .B(n586), .Z(n597) );
  XNOR2_X1 U467 ( .A(n447), .B(n531), .ZN(n726) );
  XNOR2_X1 U468 ( .A(n530), .B(n741), .ZN(n447) );
  XNOR2_X1 U469 ( .A(n556), .B(n442), .ZN(n719) );
  XNOR2_X1 U470 ( .A(n555), .B(n557), .ZN(n442) );
  XNOR2_X1 U471 ( .A(G107), .B(KEYINPUT71), .ZN(n474) );
  NAND2_X1 U472 ( .A1(n481), .A2(n419), .ZN(n480) );
  INV_X1 U473 ( .A(n683), .ZN(n481) );
  INV_X1 U474 ( .A(KEYINPUT79), .ZN(n399) );
  INV_X1 U475 ( .A(KEYINPUT34), .ZN(n422) );
  AND2_X1 U476 ( .A1(n597), .A2(n613), .ZN(n492) );
  INV_X1 U477 ( .A(n585), .ZN(n427) );
  INV_X1 U478 ( .A(n669), .ZN(n438) );
  INV_X1 U479 ( .A(n726), .ZN(n402) );
  XNOR2_X1 U480 ( .A(n606), .B(KEYINPUT46), .ZN(n607) );
  INV_X1 U481 ( .A(n655), .ZN(n452) );
  XNOR2_X1 U482 ( .A(n516), .B(n440), .ZN(n532) );
  XNOR2_X1 U483 ( .A(KEYINPUT90), .B(KEYINPUT20), .ZN(n440) );
  INV_X1 U484 ( .A(KEYINPUT44), .ZN(n484) );
  NAND2_X1 U485 ( .A1(n532), .A2(G217), .ZN(n445) );
  XNOR2_X1 U486 ( .A(G128), .B(KEYINPUT23), .ZN(n526) );
  INV_X1 U487 ( .A(KEYINPUT10), .ZN(n441) );
  XNOR2_X1 U488 ( .A(n449), .B(n448), .ZN(n536) );
  INV_X1 U489 ( .A(KEYINPUT8), .ZN(n448) );
  NAND2_X1 U490 ( .A1(n731), .A2(G234), .ZN(n449) );
  XNOR2_X1 U491 ( .A(G122), .B(n424), .ZN(n547) );
  XNOR2_X1 U492 ( .A(n741), .B(KEYINPUT12), .ZN(n553) );
  INV_X1 U493 ( .A(KEYINPUT97), .ZN(n550) );
  XOR2_X1 U494 ( .A(G131), .B(G140), .Z(n549) );
  XOR2_X1 U495 ( .A(G134), .B(G131), .Z(n740) );
  INV_X1 U496 ( .A(KEYINPUT77), .ZN(n462) );
  INV_X1 U497 ( .A(KEYINPUT74), .ZN(n647) );
  OR2_X1 U498 ( .A1(G902), .A2(G237), .ZN(n572) );
  XNOR2_X1 U499 ( .A(n512), .B(n503), .ZN(n466) );
  XNOR2_X1 U500 ( .A(G116), .B(KEYINPUT100), .ZN(n541) );
  XOR2_X1 U501 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n542) );
  INV_X1 U502 ( .A(KEYINPUT41), .ZN(n434) );
  XNOR2_X1 U503 ( .A(n475), .B(n473), .ZN(n472) );
  XNOR2_X1 U504 ( .A(n577), .B(n474), .ZN(n473) );
  XNOR2_X1 U505 ( .A(n739), .B(n578), .ZN(n475) );
  AND2_X1 U506 ( .A1(n480), .A2(n731), .ZN(n479) );
  INV_X1 U507 ( .A(KEYINPUT35), .ZN(n467) );
  INV_X1 U508 ( .A(KEYINPUT32), .ZN(n390) );
  NAND2_X1 U509 ( .A1(n432), .A2(n638), .ZN(n431) );
  INV_X1 U510 ( .A(n391), .ZN(n709) );
  XNOR2_X1 U511 ( .A(n491), .B(KEYINPUT109), .ZN(n490) );
  INV_X1 U512 ( .A(KEYINPUT105), .ZN(n486) );
  AND2_X1 U513 ( .A1(n438), .A2(n630), .ZN(n435) );
  INV_X1 U514 ( .A(KEYINPUT122), .ZN(n387) );
  INV_X1 U515 ( .A(n635), .ZN(n432) );
  XOR2_X1 U516 ( .A(n596), .B(KEYINPUT47), .Z(n375) );
  AND2_X1 U517 ( .A1(n683), .A2(KEYINPUT119), .ZN(n377) );
  XNOR2_X1 U518 ( .A(KEYINPUT113), .B(KEYINPUT36), .ZN(n378) );
  XNOR2_X1 U519 ( .A(KEYINPUT2), .B(KEYINPUT75), .ZN(n379) );
  XOR2_X1 U520 ( .A(n686), .B(KEYINPUT65), .Z(n380) );
  XOR2_X1 U521 ( .A(n684), .B(KEYINPUT62), .Z(n381) );
  XOR2_X1 U522 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n382) );
  BUF_X1 U523 ( .A(n457), .Z(n383) );
  BUF_X1 U524 ( .A(n716), .Z(n384) );
  BUF_X1 U525 ( .A(n565), .Z(n385) );
  BUF_X1 U526 ( .A(n485), .Z(n386) );
  XNOR2_X1 U527 ( .A(n388), .B(n387), .ZN(G66) );
  NAND2_X1 U528 ( .A1(n401), .A2(n355), .ZN(n388) );
  XNOR2_X1 U529 ( .A(n451), .B(KEYINPUT101), .ZN(n450) );
  BUF_X1 U530 ( .A(n754), .Z(n389) );
  XNOR2_X1 U531 ( .A(n425), .B(KEYINPUT103), .ZN(n754) );
  XNOR2_X1 U532 ( .A(n417), .B(n467), .ZN(n485) );
  XNOR2_X1 U533 ( .A(n423), .B(n422), .ZN(n418) );
  XNOR2_X1 U534 ( .A(n641), .B(n392), .ZN(n391) );
  XOR2_X1 U535 ( .A(KEYINPUT31), .B(KEYINPUT96), .Z(n392) );
  BUF_X1 U536 ( .A(n622), .Z(n393) );
  NAND2_X1 U537 ( .A1(n400), .A2(n379), .ZN(n646) );
  INV_X1 U538 ( .A(n398), .ZN(n395) );
  NAND2_X1 U539 ( .A1(n398), .A2(n377), .ZN(n397) );
  INV_X1 U540 ( .A(n400), .ZN(n469) );
  NAND2_X1 U541 ( .A1(n724), .A2(G475), .ZN(n720) );
  XNOR2_X1 U542 ( .A(n725), .B(n402), .ZN(n401) );
  XNOR2_X1 U543 ( .A(n404), .B(G101), .ZN(n729) );
  XNOR2_X2 U544 ( .A(n405), .B(n374), .ZN(n404) );
  NAND2_X1 U545 ( .A1(n407), .A2(n406), .ZN(n405) );
  NAND2_X1 U546 ( .A1(n565), .A2(n564), .ZN(n406) );
  NAND2_X1 U547 ( .A1(n408), .A2(n577), .ZN(n407) );
  INV_X1 U548 ( .A(n565), .ZN(n408) );
  NOR2_X2 U549 ( .A1(n409), .A2(n662), .ZN(n584) );
  XNOR2_X1 U550 ( .A(n409), .B(KEYINPUT110), .ZN(n592) );
  XNOR2_X2 U551 ( .A(n579), .B(G469), .ZN(n409) );
  XNOR2_X1 U552 ( .A(n410), .B(n466), .ZN(n684) );
  XNOR2_X2 U553 ( .A(n420), .B(n500), .ZN(n410) );
  XNOR2_X1 U554 ( .A(n711), .B(KEYINPUT81), .ZN(n430) );
  XNOR2_X1 U555 ( .A(n575), .B(n378), .ZN(n411) );
  XNOR2_X2 U556 ( .A(n415), .B(G107), .ZN(n566) );
  XNOR2_X1 U557 ( .A(n687), .B(n381), .ZN(n416) );
  NAND2_X1 U558 ( .A1(n418), .A2(n633), .ZN(n417) );
  XNOR2_X2 U559 ( .A(n627), .B(n626), .ZN(n634) );
  INV_X1 U560 ( .A(KEYINPUT119), .ZN(n419) );
  XNOR2_X2 U561 ( .A(n745), .B(G101), .ZN(n420) );
  XNOR2_X1 U562 ( .A(n469), .B(n748), .ZN(n746) );
  AND2_X1 U563 ( .A1(n421), .A2(n438), .ZN(n437) );
  XNOR2_X1 U564 ( .A(n421), .B(KEYINPUT108), .ZN(n428) );
  NAND2_X1 U565 ( .A1(n640), .A2(n649), .ZN(n423) );
  NOR2_X1 U566 ( .A1(n718), .A2(G902), .ZN(n579) );
  XNOR2_X2 U567 ( .A(n426), .B(n493), .ZN(n457) );
  NAND2_X1 U568 ( .A1(n495), .A2(n494), .ZN(n426) );
  NOR2_X2 U569 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X2 U570 ( .A(n623), .B(KEYINPUT0), .ZN(n632) );
  XNOR2_X2 U571 ( .A(n594), .B(KEYINPUT19), .ZN(n622) );
  XNOR2_X2 U572 ( .A(n574), .B(n573), .ZN(n594) );
  AND2_X2 U573 ( .A1(n632), .A2(n625), .ZN(n627) );
  INV_X1 U574 ( .A(n648), .ZN(n675) );
  NAND2_X1 U575 ( .A1(n648), .A2(n604), .ZN(n605) );
  XNOR2_X1 U576 ( .A(n603), .B(n434), .ZN(n648) );
  NAND2_X1 U577 ( .A1(n391), .A2(n454), .ZN(n453) );
  XNOR2_X2 U578 ( .A(n509), .B(n510), .ZN(n565) );
  NOR2_X2 U579 ( .A1(n754), .A2(n450), .ZN(n645) );
  NAND2_X1 U580 ( .A1(n483), .A2(n755), .ZN(n482) );
  INV_X1 U581 ( .A(n383), .ZN(n730) );
  XNOR2_X1 U582 ( .A(n645), .B(KEYINPUT104), .ZN(n494) );
  AND2_X2 U583 ( .A1(n640), .A2(n437), .ZN(n691) );
  XNOR2_X2 U584 ( .A(n439), .B(n446), .ZN(n636) );
  XNOR2_X1 U585 ( .A(n580), .B(n561), .ZN(n588) );
  NAND2_X1 U586 ( .A1(n614), .A2(n706), .ZN(n443) );
  NAND2_X1 U587 ( .A1(n453), .A2(n452), .ZN(n451) );
  INV_X1 U588 ( .A(n691), .ZN(n454) );
  XNOR2_X2 U589 ( .A(n539), .B(KEYINPUT4), .ZN(n745) );
  NAND2_X1 U590 ( .A1(n458), .A2(n456), .ZN(n459) );
  NAND2_X1 U591 ( .A1(n457), .A2(n379), .ZN(n456) );
  XNOR2_X1 U592 ( .A(n646), .B(n462), .ZN(n458) );
  XNOR2_X1 U593 ( .A(n459), .B(n647), .ZN(n460) );
  NAND2_X1 U594 ( .A1(n464), .A2(n469), .ZN(n463) );
  NOR2_X1 U595 ( .A1(n457), .A2(n465), .ZN(n464) );
  INV_X1 U596 ( .A(KEYINPUT2), .ZN(n465) );
  INV_X1 U597 ( .A(n386), .ZN(n757) );
  NAND2_X1 U598 ( .A1(n470), .A2(n469), .ZN(n468) );
  XNOR2_X1 U599 ( .A(n471), .B(KEYINPUT78), .ZN(n470) );
  NOR2_X2 U600 ( .A1(n457), .A2(n515), .ZN(n471) );
  XNOR2_X1 U601 ( .A(n488), .B(n382), .ZN(G75) );
  XNOR2_X1 U602 ( .A(n482), .B(n484), .ZN(n495) );
  XNOR2_X2 U603 ( .A(G119), .B(KEYINPUT3), .ZN(n510) );
  XNOR2_X2 U604 ( .A(n477), .B(n476), .ZN(n539) );
  INV_X1 U605 ( .A(n489), .ZN(n701) );
  NAND2_X1 U606 ( .A1(n490), .A2(n633), .ZN(n489) );
  NAND2_X1 U607 ( .A1(n598), .A2(n492), .ZN(n491) );
  NOR2_X1 U608 ( .A1(n496), .A2(n727), .ZN(G54) );
  XNOR2_X1 U609 ( .A(n498), .B(n497), .ZN(n496) );
  XNOR2_X1 U610 ( .A(n718), .B(n717), .ZN(n497) );
  NAND2_X1 U611 ( .A1(n724), .A2(G469), .ZN(n498) );
  XNOR2_X1 U612 ( .A(KEYINPUT59), .B(KEYINPUT121), .ZN(n499) );
  INV_X1 U613 ( .A(KEYINPUT80), .ZN(n606) );
  XNOR2_X1 U614 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U615 ( .A(n511), .B(n385), .ZN(n512) );
  NOR2_X1 U616 ( .A1(n653), .A2(n624), .ZN(n625) );
  XNOR2_X1 U617 ( .A(n740), .B(G146), .ZN(n500) );
  XNOR2_X1 U618 ( .A(n558), .B(G475), .ZN(n559) );
  INV_X1 U619 ( .A(KEYINPUT93), .ZN(n583) );
  INV_X1 U620 ( .A(KEYINPUT63), .ZN(n688) );
  XNOR2_X1 U621 ( .A(n688), .B(KEYINPUT84), .ZN(n689) );
  NOR2_X1 U622 ( .A1(G952), .A2(n731), .ZN(n727) );
  INV_X1 U623 ( .A(KEYINPUT6), .ZN(n514) );
  XOR2_X1 U624 ( .A(n502), .B(n501), .Z(n503) );
  XOR2_X1 U625 ( .A(KEYINPUT69), .B(n504), .Z(n554) );
  NAND2_X1 U626 ( .A1(n554), .A2(G210), .ZN(n511) );
  NAND2_X1 U627 ( .A1(G113), .A2(n505), .ZN(n508) );
  NAND2_X1 U628 ( .A1(n506), .A2(G116), .ZN(n507) );
  NOR2_X1 U629 ( .A1(n684), .A2(G902), .ZN(n513) );
  XOR2_X1 U630 ( .A(KEYINPUT21), .B(KEYINPUT92), .Z(n518) );
  INV_X1 U631 ( .A(n685), .ZN(n515) );
  NAND2_X1 U632 ( .A1(n515), .A2(G234), .ZN(n516) );
  NAND2_X1 U633 ( .A1(G221), .A2(n532), .ZN(n517) );
  XNOR2_X1 U634 ( .A(n518), .B(n517), .ZN(n660) );
  NAND2_X1 U635 ( .A1(G234), .A2(G237), .ZN(n519) );
  XNOR2_X1 U636 ( .A(n519), .B(KEYINPUT14), .ZN(n520) );
  NAND2_X1 U637 ( .A1(n520), .A2(G952), .ZN(n680) );
  NOR2_X1 U638 ( .A1(G953), .A2(n680), .ZN(n620) );
  NAND2_X1 U639 ( .A1(n520), .A2(G902), .ZN(n521) );
  XOR2_X1 U640 ( .A(KEYINPUT87), .B(n521), .Z(n618) );
  OR2_X1 U641 ( .A1(n618), .A2(n731), .ZN(n522) );
  NOR2_X1 U642 ( .A1(G900), .A2(n522), .ZN(n523) );
  NOR2_X1 U643 ( .A1(n620), .A2(n523), .ZN(n585) );
  INV_X1 U644 ( .A(n576), .ZN(n524) );
  XNOR2_X1 U645 ( .A(n525), .B(n524), .ZN(n529) );
  XOR2_X1 U646 ( .A(KEYINPUT24), .B(KEYINPUT89), .Z(n527) );
  XNOR2_X1 U647 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U648 ( .A(n529), .B(n528), .Z(n531) );
  NAND2_X1 U649 ( .A1(G221), .A2(n536), .ZN(n530) );
  XOR2_X1 U650 ( .A(KEYINPUT25), .B(KEYINPUT91), .Z(n533) );
  NOR2_X1 U651 ( .A1(n585), .A2(n636), .ZN(n534) );
  NAND2_X1 U652 ( .A1(n660), .A2(n534), .ZN(n589) );
  XNOR2_X1 U653 ( .A(n535), .B(KEYINPUT106), .ZN(n563) );
  XOR2_X1 U654 ( .A(n566), .B(G134), .Z(n538) );
  NAND2_X1 U655 ( .A1(G217), .A2(n536), .ZN(n537) );
  XNOR2_X1 U656 ( .A(n538), .B(n537), .ZN(n545) );
  BUF_X1 U657 ( .A(n539), .Z(n540) );
  XNOR2_X1 U658 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U659 ( .A(n540), .B(n543), .Z(n544) );
  XNOR2_X1 U660 ( .A(n545), .B(n544), .ZN(n722) );
  NOR2_X1 U661 ( .A1(G902), .A2(n722), .ZN(n546) );
  XOR2_X1 U662 ( .A(G478), .B(n546), .Z(n581) );
  INV_X1 U663 ( .A(KEYINPUT99), .ZN(n561) );
  XNOR2_X1 U664 ( .A(n547), .B(KEYINPUT11), .ZN(n557) );
  XNOR2_X1 U665 ( .A(G104), .B(n700), .ZN(n548) );
  XNOR2_X1 U666 ( .A(n549), .B(n548), .ZN(n551) );
  XNOR2_X1 U667 ( .A(n553), .B(n552), .ZN(n556) );
  NAND2_X1 U668 ( .A1(n554), .A2(G214), .ZN(n555) );
  NOR2_X1 U669 ( .A1(G902), .A2(n719), .ZN(n560) );
  XNOR2_X1 U670 ( .A(KEYINPUT98), .B(KEYINPUT13), .ZN(n558) );
  XNOR2_X1 U671 ( .A(n560), .B(n559), .ZN(n580) );
  INV_X1 U672 ( .A(n588), .ZN(n562) );
  INV_X1 U673 ( .A(n577), .ZN(n564) );
  NAND2_X1 U674 ( .A1(G224), .A2(n731), .ZN(n569) );
  NOR2_X2 U675 ( .A1(n716), .A2(n685), .ZN(n571) );
  NAND2_X1 U676 ( .A1(G210), .A2(n572), .ZN(n570) );
  NAND2_X1 U677 ( .A1(n582), .A2(n650), .ZN(n574) );
  INV_X1 U678 ( .A(KEYINPUT82), .ZN(n573) );
  NAND2_X1 U679 ( .A1(n609), .A2(n594), .ZN(n575) );
  XNOR2_X1 U680 ( .A(KEYINPUT88), .B(n576), .ZN(n739) );
  NAND2_X1 U681 ( .A1(G227), .A2(n731), .ZN(n578) );
  INV_X1 U682 ( .A(n663), .ZN(n628) );
  XNOR2_X1 U683 ( .A(KEYINPUT83), .B(n628), .ZN(n635) );
  INV_X1 U684 ( .A(n580), .ZN(n602) );
  INV_X1 U685 ( .A(n581), .ZN(n601) );
  NOR2_X1 U686 ( .A1(n602), .A2(n601), .ZN(n633) );
  BUF_X2 U687 ( .A(n582), .Z(n613) );
  NAND2_X1 U688 ( .A1(n669), .A2(n650), .ZN(n586) );
  XNOR2_X1 U689 ( .A(KEYINPUT76), .B(n701), .ZN(n587) );
  NOR2_X1 U690 ( .A1(n601), .A2(n588), .ZN(n708) );
  NOR2_X1 U691 ( .A1(n706), .A2(n708), .ZN(n655) );
  NOR2_X1 U692 ( .A1(n438), .A2(n589), .ZN(n591) );
  XNOR2_X1 U693 ( .A(KEYINPUT111), .B(KEYINPUT28), .ZN(n590) );
  XNOR2_X1 U694 ( .A(n591), .B(n590), .ZN(n593) );
  NOR2_X1 U695 ( .A1(n593), .A2(n592), .ZN(n604) );
  INV_X1 U696 ( .A(n393), .ZN(n595) );
  NAND2_X1 U697 ( .A1(n604), .A2(n595), .ZN(n703) );
  NOR2_X1 U698 ( .A1(n655), .A2(n703), .ZN(n596) );
  XOR2_X1 U699 ( .A(KEYINPUT112), .B(KEYINPUT40), .Z(n600) );
  AND2_X1 U700 ( .A1(n597), .A2(n651), .ZN(n599) );
  NAND2_X1 U701 ( .A1(n651), .A2(n650), .ZN(n654) );
  NAND2_X1 U702 ( .A1(n602), .A2(n601), .ZN(n653) );
  NOR2_X1 U703 ( .A1(n654), .A2(n653), .ZN(n603) );
  NAND2_X1 U704 ( .A1(n609), .A2(n650), .ZN(n610) );
  NOR2_X1 U705 ( .A1(n628), .A2(n610), .ZN(n611) );
  XNOR2_X1 U706 ( .A(n611), .B(KEYINPUT43), .ZN(n612) );
  NOR2_X1 U707 ( .A1(n613), .A2(n612), .ZN(n714) );
  NAND2_X1 U708 ( .A1(n708), .A2(n614), .ZN(n713) );
  INV_X1 U709 ( .A(n713), .ZN(n615) );
  NOR2_X1 U710 ( .A1(n714), .A2(n615), .ZN(n616) );
  INV_X1 U711 ( .A(n636), .ZN(n630) );
  NOR2_X1 U712 ( .A1(G898), .A2(n731), .ZN(n617) );
  XOR2_X1 U713 ( .A(KEYINPUT86), .B(n617), .Z(n728) );
  NOR2_X1 U714 ( .A1(n618), .A2(n728), .ZN(n619) );
  INV_X1 U715 ( .A(n660), .ZN(n624) );
  INV_X1 U716 ( .A(n642), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n639), .A2(n637), .ZN(n631) );
  XNOR2_X1 U718 ( .A(KEYINPUT102), .B(n636), .ZN(n659) );
  NOR2_X1 U719 ( .A1(n637), .A2(n659), .ZN(n638) );
  NAND2_X1 U720 ( .A1(n632), .A2(n672), .ZN(n641) );
  AND2_X1 U721 ( .A1(n659), .A2(n642), .ZN(n643) );
  AND2_X1 U722 ( .A1(n649), .A2(n648), .ZN(n682) );
  NOR2_X1 U723 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U724 ( .A1(n653), .A2(n652), .ZN(n657) );
  NOR2_X1 U725 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U726 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U727 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U728 ( .A(KEYINPUT49), .B(n661), .ZN(n667) );
  XOR2_X1 U729 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n665) );
  NAND2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U731 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U732 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U733 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U734 ( .A(n670), .B(KEYINPUT118), .ZN(n671) );
  NOR2_X1 U735 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U736 ( .A(KEYINPUT51), .B(n673), .Z(n674) );
  NOR2_X1 U737 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U738 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U739 ( .A(n678), .B(KEYINPUT52), .ZN(n679) );
  NOR2_X1 U740 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U741 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U742 ( .A1(n685), .A2(KEYINPUT2), .ZN(n686) );
  NAND2_X1 U743 ( .A1(n724), .A2(G472), .ZN(n687) );
  NAND2_X1 U744 ( .A1(n691), .A2(n706), .ZN(n690) );
  XNOR2_X1 U745 ( .A(n690), .B(G104), .ZN(G6) );
  XNOR2_X1 U746 ( .A(G107), .B(KEYINPUT27), .ZN(n695) );
  XOR2_X1 U747 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n693) );
  NAND2_X1 U748 ( .A1(n691), .A2(n708), .ZN(n692) );
  XNOR2_X1 U749 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U750 ( .A(n695), .B(n694), .ZN(G9) );
  INV_X1 U751 ( .A(n708), .ZN(n696) );
  NOR2_X1 U752 ( .A1(n696), .A2(n703), .ZN(n698) );
  XNOR2_X1 U753 ( .A(KEYINPUT115), .B(KEYINPUT29), .ZN(n697) );
  XNOR2_X1 U754 ( .A(n698), .B(n697), .ZN(n699) );
  XOR2_X1 U755 ( .A(G128), .B(n699), .Z(G30) );
  XOR2_X1 U756 ( .A(n701), .B(n700), .Z(n702) );
  XNOR2_X1 U757 ( .A(KEYINPUT116), .B(n702), .ZN(G45) );
  INV_X1 U758 ( .A(n706), .ZN(n704) );
  NOR2_X1 U759 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U760 ( .A(G146), .B(n705), .Z(G48) );
  NAND2_X1 U761 ( .A1(n709), .A2(n706), .ZN(n707) );
  XNOR2_X1 U762 ( .A(n707), .B(n424), .ZN(G15) );
  NAND2_X1 U763 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U764 ( .A(n710), .B(G116), .ZN(G18) );
  XNOR2_X1 U765 ( .A(n711), .B(G125), .ZN(n712) );
  XNOR2_X1 U766 ( .A(n712), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U767 ( .A(G134), .B(n713), .ZN(G36) );
  XOR2_X1 U768 ( .A(G140), .B(n714), .Z(G42) );
  XOR2_X1 U769 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n715) );
  XOR2_X1 U770 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n717) );
  NAND2_X1 U771 ( .A1(G478), .A2(n724), .ZN(n721) );
  XNOR2_X1 U772 ( .A(n722), .B(n721), .ZN(n723) );
  NOR2_X1 U773 ( .A1(n727), .A2(n723), .ZN(G63) );
  NAND2_X1 U774 ( .A1(G217), .A2(n724), .ZN(n725) );
  NAND2_X1 U775 ( .A1(n729), .A2(n728), .ZN(n738) );
  NAND2_X1 U776 ( .A1(n731), .A2(n730), .ZN(n735) );
  NAND2_X1 U777 ( .A1(G953), .A2(G224), .ZN(n732) );
  XNOR2_X1 U778 ( .A(KEYINPUT61), .B(n732), .ZN(n733) );
  NAND2_X1 U779 ( .A1(n733), .A2(G898), .ZN(n734) );
  NAND2_X1 U780 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U781 ( .A(n736), .B(KEYINPUT123), .ZN(n737) );
  XNOR2_X1 U782 ( .A(n738), .B(n737), .ZN(G69) );
  XOR2_X1 U783 ( .A(KEYINPUT124), .B(n739), .Z(n743) );
  XNOR2_X1 U784 ( .A(n741), .B(n740), .ZN(n742) );
  XNOR2_X1 U785 ( .A(n743), .B(n742), .ZN(n744) );
  XOR2_X1 U786 ( .A(n745), .B(n744), .Z(n748) );
  NOR2_X1 U787 ( .A1(G953), .A2(n746), .ZN(n747) );
  XNOR2_X1 U788 ( .A(n747), .B(KEYINPUT125), .ZN(n752) );
  XNOR2_X1 U789 ( .A(G227), .B(n748), .ZN(n749) );
  NAND2_X1 U790 ( .A1(n749), .A2(G900), .ZN(n750) );
  NAND2_X1 U791 ( .A1(G953), .A2(n750), .ZN(n751) );
  NAND2_X1 U792 ( .A1(n752), .A2(n751), .ZN(G72) );
  XOR2_X1 U793 ( .A(n753), .B(G131), .Z(G33) );
  XOR2_X1 U794 ( .A(n389), .B(G101), .Z(G3) );
  XNOR2_X1 U795 ( .A(n755), .B(G110), .ZN(G12) );
  XNOR2_X1 U796 ( .A(n756), .B(G119), .ZN(G21) );
  XOR2_X1 U797 ( .A(G122), .B(n757), .Z(n758) );
  XNOR2_X1 U798 ( .A(KEYINPUT126), .B(n758), .ZN(G24) );
  XOR2_X1 U799 ( .A(G137), .B(n759), .Z(G39) );
endmodule

