//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  INV_X1    g000(.A(KEYINPUT65), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  AND3_X1   g007(.A1(new_n189), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  OAI22_X1  g008(.A1(new_n189), .A2(new_n193), .B1(new_n191), .B2(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G137), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(KEYINPUT11), .A3(G134), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(G137), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n199), .A2(new_n201), .A3(new_n202), .A4(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n198), .A2(G137), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n200), .A2(G134), .ZN(new_n206));
  OAI21_X1  g020(.A(G131), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n196), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n199), .A2(new_n201), .A3(new_n203), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G131), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n192), .A2(G146), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n190), .A2(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT0), .A2(G128), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(KEYINPUT0), .A2(G128), .ZN(new_n216));
  OAI22_X1  g030(.A1(new_n212), .A2(new_n213), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G143), .B(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(new_n214), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n211), .A2(new_n204), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n187), .B(KEYINPUT30), .C1(new_n209), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n211), .A2(new_n204), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n217), .A2(new_n219), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G128), .ZN(new_n226));
  AOI22_X1  g040(.A1(new_n188), .A2(new_n212), .B1(new_n213), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n218), .A2(new_n189), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(new_n204), .A3(new_n207), .ZN(new_n230));
  OR2_X1    g044(.A1(new_n187), .A2(KEYINPUT30), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n187), .A2(KEYINPUT30), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n224), .A2(new_n230), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n221), .A2(new_n233), .ZN(new_n234));
  OR2_X1    g048(.A1(KEYINPUT2), .A2(G113), .ZN(new_n235));
  NAND3_X1  g049(.A1(KEYINPUT64), .A2(KEYINPUT2), .A3(G113), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT64), .B1(KEYINPUT2), .B2(G113), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n235), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G119), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G116), .ZN(new_n241));
  INV_X1    g055(.A(G116), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G119), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n239), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT2), .A2(G113), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT64), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n236), .ZN(new_n249));
  XNOR2_X1  g063(.A(G116), .B(G119), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n235), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n234), .A2(new_n252), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n245), .A2(new_n251), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n224), .A2(new_n254), .A3(new_n230), .ZN(new_n255));
  INV_X1    g069(.A(G237), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT66), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G237), .ZN(new_n259));
  AOI21_X1  g073(.A(G953), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G210), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G101), .ZN(new_n262));
  INV_X1    g076(.A(G101), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n263), .A3(G210), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n265), .B1(new_n262), .B2(new_n264), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n253), .A2(new_n255), .A3(new_n268), .ZN(new_n269));
  NOR3_X1   g083(.A1(new_n209), .A2(new_n220), .A3(new_n252), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n254), .B1(new_n224), .B2(new_n230), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT28), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT28), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n255), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n268), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n269), .B1(new_n275), .B2(KEYINPUT31), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT31), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n253), .A2(new_n277), .A3(new_n255), .A4(new_n268), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT67), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n270), .B1(new_n234), .B2(new_n252), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT67), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n280), .A2(new_n281), .A3(new_n277), .A4(new_n268), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n276), .A2(new_n279), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G472), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT68), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n283), .A2(new_n288), .A3(new_n284), .A4(new_n285), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT32), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n283), .A2(KEYINPUT32), .A3(new_n284), .A4(new_n285), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n272), .A2(new_n268), .A3(new_n274), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT29), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n294), .B(new_n295), .C1(new_n280), .C2(new_n268), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n296), .B(new_n285), .C1(new_n295), .C2(new_n294), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G472), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n188), .A2(G119), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI211_X1 g118(.A(KEYINPUT71), .B(KEYINPUT23), .C1(new_n188), .C2(G119), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G110), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n240), .A2(G128), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n306), .A2(KEYINPUT73), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(G119), .B(G128), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n310), .A2(KEYINPUT69), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(KEYINPUT69), .ZN(new_n312));
  OR2_X1    g126(.A1(KEYINPUT24), .A2(G110), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT70), .ZN(new_n314));
  NAND2_X1  g128(.A1(KEYINPUT24), .A2(G110), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n314), .B1(new_n313), .B2(new_n315), .ZN(new_n317));
  OAI22_X1  g131(.A1(new_n311), .A2(new_n312), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n303), .B1(new_n240), .B2(G128), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT23), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n302), .A2(new_n303), .A3(new_n301), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n320), .A2(new_n321), .A3(new_n307), .A4(new_n308), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT73), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n309), .A2(new_n318), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT16), .ZN(new_n326));
  INV_X1    g140(.A(G125), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(KEYINPUT72), .A2(G125), .ZN(new_n329));
  INV_X1    g143(.A(G140), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(KEYINPUT72), .A2(G125), .A3(G140), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n328), .B1(new_n333), .B2(new_n326), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G146), .ZN(new_n335));
  XNOR2_X1  g149(.A(G125), .B(G140), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n190), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n325), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n311), .A2(new_n312), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n316), .A2(new_n317), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n306), .A2(new_n308), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G110), .ZN(new_n343));
  INV_X1    g157(.A(new_n335), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n334), .A2(G146), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n341), .B(new_n343), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT22), .B(G137), .ZN(new_n347));
  INV_X1    g161(.A(G953), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(G221), .A3(G234), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n347), .B(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n338), .A2(new_n346), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT75), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT75), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n338), .A2(new_n353), .A3(new_n346), .A4(new_n350), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n338), .A2(new_n346), .ZN(new_n356));
  INV_X1    g170(.A(new_n350), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT74), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT74), .ZN(new_n359));
  AOI211_X1 g173(.A(new_n359), .B(new_n350), .C1(new_n338), .C2(new_n346), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n355), .B(new_n285), .C1(new_n358), .C2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT76), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(KEYINPUT25), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n358), .A2(new_n360), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n366), .A2(new_n285), .A3(new_n355), .A4(new_n363), .ZN(new_n367));
  INV_X1    g181(.A(G217), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n368), .B1(G234), .B2(new_n285), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n365), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(G902), .ZN(new_n371));
  XOR2_X1   g185(.A(new_n371), .B(KEYINPUT77), .Z(new_n372));
  NAND3_X1  g186(.A1(new_n366), .A2(new_n372), .A3(new_n355), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT78), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n370), .A2(new_n373), .A3(KEYINPUT78), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n292), .A2(new_n300), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n377), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT78), .B1(new_n370), .B2(new_n373), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT32), .B1(new_n287), .B2(new_n289), .ZN(new_n383));
  OAI22_X1  g197(.A1(new_n381), .A2(new_n382), .B1(new_n383), .B2(new_n299), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT79), .ZN(new_n385));
  INV_X1    g199(.A(G107), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(G104), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n386), .A2(KEYINPUT3), .A3(G104), .ZN(new_n389));
  AOI21_X1  g203(.A(KEYINPUT3), .B1(new_n386), .B2(G104), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(KEYINPUT80), .A2(KEYINPUT4), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(G101), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT3), .ZN(new_n395));
  INV_X1    g209(.A(G104), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n395), .B1(new_n396), .B2(G107), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n386), .A2(KEYINPUT3), .A3(G104), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n387), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n392), .B1(new_n399), .B2(new_n263), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n399), .A2(new_n263), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n394), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n223), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n388), .B(new_n263), .C1(new_n389), .C2(new_n390), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT81), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n386), .B2(G104), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n386), .A2(G104), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n396), .A2(KEYINPUT81), .A3(G107), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G101), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT82), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n189), .A2(new_n191), .A3(new_n193), .A4(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n213), .A2(new_n226), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n212), .A2(new_n188), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n411), .B1(new_n218), .B2(new_n189), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n404), .B(new_n410), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT10), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n410), .A2(new_n404), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n418), .B1(new_n227), .B2(new_n228), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n403), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  XOR2_X1   g238(.A(new_n222), .B(KEYINPUT83), .Z(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G110), .B(G140), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n348), .A2(G227), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n427), .B(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n423), .A2(KEYINPUT84), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n417), .A2(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT84), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n433), .A3(new_n403), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n431), .A2(new_n222), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT85), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT85), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n431), .A2(new_n437), .A3(new_n222), .A4(new_n434), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n430), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n417), .B1(new_n229), .B2(new_n420), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n222), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT12), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n441), .B(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n429), .B1(new_n443), .B2(new_n426), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n285), .B1(new_n439), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G469), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT86), .ZN(new_n447));
  INV_X1    g261(.A(new_n426), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(new_n436), .B2(new_n438), .ZN(new_n449));
  INV_X1    g263(.A(new_n443), .ZN(new_n450));
  OAI22_X1  g264(.A1(new_n449), .A2(new_n429), .B1(new_n450), .B2(new_n430), .ZN(new_n451));
  XOR2_X1   g265(.A(KEYINPUT87), .B(G469), .Z(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n451), .A2(new_n285), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT86), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n436), .A2(new_n438), .ZN(new_n456));
  INV_X1    g270(.A(new_n430), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n444), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n455), .B(G469), .C1(new_n458), .C2(G902), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n447), .A2(new_n454), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G221), .ZN(new_n461));
  XOR2_X1   g275(.A(KEYINPUT9), .B(G234), .Z(new_n462));
  AOI21_X1  g276(.A(new_n461), .B1(new_n462), .B2(new_n285), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(G214), .B1(G237), .B2(G902), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n348), .A2(G952), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n468), .B1(G234), .B2(G237), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(G898), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT92), .ZN(new_n471));
  AOI211_X1 g285(.A(new_n285), .B(new_n348), .C1(G234), .C2(G237), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT88), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n241), .A2(new_n243), .A3(KEYINPUT5), .ZN(new_n475));
  OAI21_X1  g289(.A(G113), .B1(new_n241), .B2(KEYINPUT5), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G113), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n242), .A2(G119), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT5), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n481), .B(KEYINPUT88), .C1(new_n244), .C2(new_n480), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT89), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n483), .A2(new_n484), .A3(new_n251), .A4(new_n420), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n477), .A2(new_n482), .A3(new_n251), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n410), .A2(new_n404), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT89), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n402), .A2(new_n252), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  XOR2_X1   g304(.A(G110), .B(G122), .Z(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n491), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n485), .A2(new_n488), .A3(new_n493), .A4(new_n489), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(KEYINPUT6), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n229), .A2(new_n327), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n223), .A2(G125), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n348), .A2(G224), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n498), .B(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT6), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n490), .A2(new_n501), .A3(new_n491), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n495), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT7), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n251), .B1(new_n475), .B2(new_n476), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n420), .A2(new_n507), .ZN(new_n508));
  XOR2_X1   g322(.A(new_n491), .B(KEYINPUT8), .Z(new_n509));
  OAI211_X1 g323(.A(new_n508), .B(new_n509), .C1(new_n420), .C2(new_n486), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n496), .A2(new_n497), .A3(new_n504), .A4(new_n499), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n506), .A2(new_n494), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n503), .A2(new_n285), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(G210), .B1(G237), .B2(G902), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n503), .A2(new_n285), .A3(new_n514), .A4(new_n512), .ZN(new_n517));
  AOI211_X1 g331(.A(new_n467), .B(new_n473), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(G128), .B(G143), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT13), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n192), .A2(G128), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n520), .B(G134), .C1(KEYINPUT13), .C2(new_n521), .ZN(new_n522));
  XOR2_X1   g336(.A(G116), .B(G122), .Z(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G107), .ZN(new_n524));
  XNOR2_X1  g338(.A(G116), .B(G122), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n386), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n519), .A2(new_n198), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n522), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n519), .B(new_n198), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n242), .A2(KEYINPUT14), .A3(G122), .ZN(new_n531));
  OAI211_X1 g345(.A(G107), .B(new_n531), .C1(new_n523), .C2(KEYINPUT14), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(new_n526), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n462), .A2(G217), .A3(new_n348), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n534), .A2(new_n535), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(G902), .ZN(new_n539));
  INV_X1    g353(.A(G478), .ZN(new_n540));
  OR2_X1    g354(.A1(new_n540), .A2(KEYINPUT15), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n539), .B(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n257), .A2(new_n259), .ZN(new_n544));
  AND4_X1   g358(.A1(G143), .A2(new_n544), .A3(G214), .A4(new_n348), .ZN(new_n545));
  AOI21_X1  g359(.A(G143), .B1(new_n260), .B2(G214), .ZN(new_n546));
  OAI21_X1  g360(.A(G131), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n258), .A2(G237), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n256), .A2(KEYINPUT66), .ZN(new_n550));
  OAI211_X1 g364(.A(G214), .B(new_n348), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n192), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n260), .A2(G143), .A3(G214), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n202), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n547), .A2(new_n548), .A3(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n344), .A2(new_n345), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n202), .B1(new_n552), .B2(new_n553), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT17), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT18), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n552), .B(new_n553), .C1(new_n560), .C2(new_n202), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n337), .B1(new_n333), .B2(new_n190), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n561), .B(new_n562), .C1(new_n547), .C2(new_n560), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(G113), .B(G122), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(new_n396), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n559), .A2(new_n566), .A3(new_n563), .ZN(new_n569));
  AOI21_X1  g383(.A(G902), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G475), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n559), .A2(new_n566), .A3(new_n563), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n331), .A2(KEYINPUT90), .A3(KEYINPUT19), .A4(new_n332), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT19), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n333), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT90), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n577), .B1(new_n336), .B2(new_n575), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n574), .B(new_n190), .C1(new_n576), .C2(new_n578), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n552), .A2(new_n202), .A3(new_n553), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n335), .B(new_n579), .C1(new_n580), .C2(new_n557), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(new_n563), .A3(KEYINPUT91), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n563), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT91), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n566), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n573), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(G475), .A2(G902), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT20), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n583), .A2(new_n584), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(new_n567), .A3(new_n582), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n569), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT20), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n587), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n572), .B1(new_n589), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n518), .A2(new_n543), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n380), .A2(new_n385), .A3(new_n465), .A4(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(G101), .ZN(G3));
  NAND2_X1  g413(.A1(new_n283), .A2(new_n285), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G472), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n460), .A2(new_n290), .A3(new_n464), .A4(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n538), .A2(KEYINPUT33), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n536), .A2(new_n537), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(G478), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n539), .A2(new_n540), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n540), .A2(new_n285), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n589), .A2(new_n594), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n566), .B1(new_n559), .B2(new_n563), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n285), .B1(new_n573), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(G475), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n611), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT93), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n467), .B1(new_n516), .B2(new_n517), .ZN(new_n618));
  INV_X1    g432(.A(new_n473), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n376), .A2(new_n377), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n603), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT34), .B(G104), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  AOI21_X1  g439(.A(new_n593), .B1(new_n592), .B2(new_n587), .ZN(new_n626));
  AOI211_X1 g440(.A(KEYINPUT20), .B(new_n588), .C1(new_n591), .C2(new_n569), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(KEYINPUT94), .B1(new_n570), .B2(new_n571), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT94), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n614), .A2(new_n630), .A3(G475), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n628), .A2(new_n632), .A3(new_n543), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(KEYINPUT95), .A3(new_n619), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n629), .A2(new_n631), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n635), .A2(new_n542), .A3(new_n612), .A4(new_n619), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT95), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n634), .A2(new_n618), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n603), .A2(new_n639), .A3(new_n622), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  NOR2_X1   g456(.A1(new_n357), .A2(KEYINPUT36), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n356), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n372), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n370), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n454), .A2(new_n459), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n455), .B1(new_n445), .B2(G469), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n464), .B(new_n646), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n290), .A2(new_n601), .ZN(new_n650));
  OR3_X1    g464(.A1(new_n649), .A2(new_n596), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT96), .B(KEYINPUT37), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G110), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n651), .B(new_n653), .ZN(G12));
  NAND2_X1  g468(.A1(new_n292), .A2(new_n300), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n655), .A2(new_n464), .A3(new_n460), .A4(new_n646), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT98), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n516), .A2(new_n517), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n466), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n469), .B(KEYINPUT97), .ZN(new_n660));
  INV_X1    g474(.A(G900), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n472), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n635), .A2(new_n542), .A3(new_n612), .A4(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n657), .B1(new_n659), .B2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n633), .A2(KEYINPUT98), .A3(new_n618), .A4(new_n664), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(KEYINPUT99), .B1(new_n656), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n383), .A2(new_n299), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n649), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT99), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n666), .A2(new_n667), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G128), .ZN(G30));
  XNOR2_X1  g490(.A(new_n663), .B(KEYINPUT39), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n465), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n615), .B1(new_n626), .B2(new_n627), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n680), .A2(new_n542), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n280), .A2(new_n266), .A3(new_n267), .ZN(new_n684));
  OR2_X1    g498(.A1(new_n270), .A2(new_n271), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n285), .B1(new_n685), .B2(new_n268), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  AOI22_X1  g501(.A1(new_n290), .A2(new_n291), .B1(G472), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT100), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n688), .A2(new_n689), .A3(new_n293), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n689), .B1(new_n688), .B2(new_n293), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n646), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n658), .B(KEYINPUT38), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n683), .A2(new_n467), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n192), .ZN(G45));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n616), .B2(new_n664), .ZN(new_n699));
  NOR4_X1   g513(.A1(new_n595), .A2(KEYINPUT101), .A3(new_n611), .A4(new_n663), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(KEYINPUT102), .A3(new_n618), .ZN(new_n702));
  INV_X1    g516(.A(new_n611), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n681), .A2(new_n703), .A3(new_n664), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(KEYINPUT101), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n616), .A2(new_n698), .A3(new_n664), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n706), .A3(new_n618), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT102), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n702), .A2(new_n671), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G146), .ZN(G48));
  INV_X1    g525(.A(KEYINPUT103), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n450), .A2(new_n430), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n432), .A2(new_n433), .A3(new_n403), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n433), .B1(new_n432), .B2(new_n403), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n437), .B1(new_n716), .B2(new_n222), .ZN(new_n717));
  INV_X1    g531(.A(new_n438), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n426), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n429), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n713), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n712), .B1(new_n721), .B2(G902), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n451), .A2(KEYINPUT103), .A3(new_n285), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(G469), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n464), .A3(new_n454), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n621), .A2(new_n726), .A3(new_n378), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT41), .B(G113), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G15));
  NAND3_X1  g543(.A1(new_n726), .A2(new_n639), .A3(new_n378), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G116), .ZN(G18));
  NAND4_X1  g545(.A1(new_n726), .A2(new_n655), .A3(new_n597), .A4(new_n646), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G119), .ZN(G21));
  NAND2_X1  g547(.A1(new_n681), .A2(new_n542), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n601), .A2(KEYINPUT104), .A3(new_n286), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  AOI211_X1 g551(.A(KEYINPUT104), .B(new_n284), .C1(new_n283), .C2(new_n285), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n374), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n726), .A2(new_n518), .A3(new_n735), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  INV_X1    g556(.A(KEYINPUT105), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n699), .A2(new_n700), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT105), .B1(new_n705), .B2(new_n706), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n646), .B1(new_n736), .B2(new_n738), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n725), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n746), .A2(new_n748), .A3(new_n618), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G125), .ZN(G27));
  NOR3_X1   g564(.A1(new_n658), .A2(new_n463), .A3(new_n467), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n454), .A2(new_n446), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n286), .A2(new_n291), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n374), .B1(new_n300), .B2(new_n754), .ZN(new_n755));
  AND4_X1   g569(.A1(KEYINPUT42), .A2(new_n746), .A3(new_n753), .A4(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n746), .A2(KEYINPUT106), .A3(new_n378), .A4(new_n753), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n743), .B1(new_n699), .B2(new_n700), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n705), .A2(new_n706), .A3(KEYINPUT105), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n378), .A2(new_n758), .A3(new_n759), .A4(new_n753), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT106), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n757), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n757), .A2(new_n762), .A3(KEYINPUT107), .A4(new_n763), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n756), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n202), .ZN(G33));
  NAND3_X1  g583(.A1(new_n633), .A2(KEYINPUT108), .A3(new_n664), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT108), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n665), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n378), .A2(new_n753), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G134), .ZN(G36));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n458), .B(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(G469), .B1(new_n776), .B2(G902), .ZN(new_n777));
  XOR2_X1   g591(.A(new_n777), .B(KEYINPUT46), .Z(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n454), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n464), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n677), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n595), .A2(new_n703), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT43), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n650), .A3(new_n646), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n658), .A2(new_n467), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT109), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n785), .B2(new_n786), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT110), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n781), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  INV_X1    g607(.A(KEYINPUT47), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n780), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n779), .A2(KEYINPUT47), .A3(new_n464), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n655), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n622), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n701), .A2(new_n788), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G140), .ZN(G42));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n803));
  INV_X1    g617(.A(new_n649), .ZN(new_n804));
  AND4_X1   g618(.A1(new_n672), .A2(new_n804), .A3(new_n655), .A4(new_n673), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n672), .B1(new_n671), .B2(new_n673), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n710), .B(new_n749), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n659), .A2(new_n734), .ZN(new_n808));
  AND4_X1   g622(.A1(new_n464), .A2(new_n808), .A3(new_n664), .A4(new_n752), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n809), .B(new_n693), .C1(new_n690), .C2(new_n691), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n803), .B1(new_n807), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n744), .A2(new_n745), .A3(new_n659), .ZN(new_n814));
  AOI22_X1  g628(.A1(new_n669), .A2(new_n674), .B1(new_n814), .B2(new_n748), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(KEYINPUT52), .A3(new_n710), .A4(new_n810), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n812), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n813), .B1(new_n812), .B2(new_n816), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n747), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n820), .A2(new_n759), .A3(new_n758), .A4(new_n753), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n821), .A2(new_n773), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n628), .A2(new_n632), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n542), .A2(new_n663), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n671), .A2(new_n823), .A3(new_n788), .A4(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT113), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n598), .A2(new_n651), .A3(new_n730), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n518), .A2(new_n828), .A3(new_n616), .ZN(new_n829));
  INV_X1    g643(.A(new_n616), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT111), .B1(new_n620), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n595), .A2(new_n542), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT112), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n832), .B(new_n833), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n829), .B(new_n831), .C1(new_n834), .C2(new_n620), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n622), .A3(new_n603), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n836), .A2(new_n727), .A3(new_n741), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n825), .A2(KEYINPUT113), .A3(new_n773), .A4(new_n821), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n827), .A2(new_n837), .A3(new_n732), .A4(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n768), .A2(new_n826), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n819), .A2(KEYINPUT53), .A3(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n807), .B2(new_n811), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT115), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n845), .B(new_n842), .C1(new_n807), .C2(new_n811), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n844), .A2(new_n816), .A3(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n840), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n841), .B1(new_n848), .B2(KEYINPUT53), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT54), .ZN(new_n850));
  INV_X1    g664(.A(new_n454), .ZN(new_n851));
  INV_X1    g665(.A(G469), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n451), .A2(new_n285), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n852), .B1(new_n853), .B2(new_n712), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n851), .B1(new_n854), .B2(new_n723), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n463), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n795), .A2(new_n796), .A3(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n784), .A2(new_n660), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n858), .A2(new_n740), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n859), .A2(new_n789), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n859), .A2(new_n726), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n694), .A2(new_n466), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT50), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n855), .A2(new_n751), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n858), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(new_n820), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n862), .A2(KEYINPUT50), .A3(new_n864), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n690), .A2(new_n691), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n873), .A2(new_n622), .A3(new_n469), .A4(new_n866), .ZN(new_n874));
  OR3_X1    g688(.A1(new_n874), .A2(new_n681), .A3(new_n703), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n861), .A2(new_n872), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n468), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n857), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n795), .A2(KEYINPUT117), .A3(new_n796), .A4(new_n856), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(new_n860), .A3(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(KEYINPUT51), .A3(new_n872), .A4(new_n875), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n874), .A2(new_n617), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n878), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n859), .A2(new_n618), .A3(new_n726), .ZN(new_n886));
  INV_X1    g700(.A(new_n818), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n812), .A2(new_n816), .A3(new_n813), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n840), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT53), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n840), .A2(new_n847), .A3(KEYINPUT53), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n850), .A2(new_n885), .A3(new_n886), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n868), .A2(new_n755), .ZN(new_n896));
  XNOR2_X1  g710(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n896), .B(new_n897), .ZN(new_n898));
  OAI22_X1  g712(.A1(new_n895), .A2(new_n898), .B1(G952), .B2(G953), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT49), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n855), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n464), .B(new_n466), .C1(new_n855), .C2(new_n900), .ZN(new_n902));
  OR3_X1    g716(.A1(new_n692), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  OR4_X1    g717(.A1(new_n374), .A2(new_n903), .A3(new_n694), .A4(new_n782), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n899), .A2(new_n904), .ZN(G75));
  AOI21_X1  g719(.A(new_n285), .B1(new_n891), .B2(new_n893), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(G210), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n495), .A2(new_n502), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(new_n500), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT55), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n907), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n911), .B1(new_n907), .B2(new_n908), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n348), .A2(G952), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(G51));
  NAND2_X1  g729(.A1(G469), .A2(G902), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT57), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n916), .A2(KEYINPUT57), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT53), .B1(new_n819), .B2(new_n840), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n840), .A2(KEYINPUT53), .A3(new_n847), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n919), .A2(new_n920), .A3(KEYINPUT54), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n892), .B1(new_n891), .B2(new_n893), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n917), .B(new_n918), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n451), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n906), .A2(G469), .A3(new_n776), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n914), .B1(new_n924), .B2(new_n925), .ZN(G54));
  INV_X1    g740(.A(new_n914), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(new_n586), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n586), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT119), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n928), .A2(KEYINPUT119), .A3(new_n586), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(G60));
  XNOR2_X1  g748(.A(new_n609), .B(KEYINPUT59), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n850), .B2(new_n894), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n604), .A2(new_n606), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT120), .Z(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n927), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n921), .A2(new_n922), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n941), .A2(new_n935), .A3(new_n938), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n940), .A2(new_n942), .ZN(G63));
  NAND2_X1  g757(.A1(G217), .A2(G902), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT60), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n644), .B(new_n946), .C1(new_n919), .C2(new_n920), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n945), .B1(new_n891), .B2(new_n893), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n366), .A2(new_n355), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT122), .Z(new_n950));
  OAI211_X1 g764(.A(new_n947), .B(new_n927), .C1(new_n948), .C2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT121), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n951), .A2(new_n952), .A3(KEYINPUT61), .ZN(new_n953));
  AOI21_X1  g767(.A(KEYINPUT61), .B1(new_n951), .B2(new_n952), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(G66));
  INV_X1    g769(.A(G224), .ZN(new_n956));
  OAI21_X1  g770(.A(G953), .B1(new_n471), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n827), .A2(new_n837), .A3(new_n732), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n959), .B2(G953), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n909), .B1(G898), .B2(new_n348), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT123), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n960), .B(new_n962), .ZN(G69));
  XNOR2_X1  g777(.A(new_n234), .B(KEYINPUT124), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n574), .B1(new_n576), .B2(new_n578), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n964), .B(new_n965), .Z(new_n966));
  INV_X1    g780(.A(new_n807), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n801), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n781), .A2(new_n755), .A3(new_n808), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n792), .A2(new_n969), .A3(new_n773), .ZN(new_n970));
  OR3_X1    g784(.A1(new_n968), .A2(new_n768), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n348), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n348), .B1(G227), .B2(G900), .ZN(new_n973));
  OR2_X1    g787(.A1(KEYINPUT126), .A2(G900), .ZN(new_n974));
  NAND2_X1  g788(.A1(KEYINPUT126), .A2(G900), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n966), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n380), .A2(new_n385), .ZN(new_n978));
  INV_X1    g792(.A(new_n679), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n834), .A2(new_n830), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n978), .A2(new_n979), .A3(new_n788), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n792), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT125), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n696), .A2(new_n807), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT62), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n983), .A2(new_n985), .A3(new_n801), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n973), .B1(new_n986), .B2(new_n348), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n977), .B1(new_n987), .B2(new_n966), .ZN(G72));
  NAND2_X1  g802(.A1(G472), .A2(G902), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT63), .Z(new_n990));
  OAI21_X1  g804(.A(new_n990), .B1(new_n971), .B2(new_n958), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT127), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI211_X1 g807(.A(new_n270), .B(new_n268), .C1(new_n234), .C2(new_n252), .ZN(new_n994));
  OAI211_X1 g808(.A(KEYINPUT127), .B(new_n990), .C1(new_n971), .C2(new_n958), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n990), .B1(new_n986), .B2(new_n958), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n914), .B1(new_n997), .B2(new_n684), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n684), .A2(new_n994), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n849), .A2(new_n990), .A3(new_n999), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n996), .A2(new_n998), .A3(new_n1000), .ZN(G57));
endmodule


