//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n572,
    new_n573, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n586, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n454), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND3_X1   g039(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT68), .B(G2105), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n465), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n474), .A2(G137), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n479), .B1(new_n469), .B2(G2104), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n467), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n480), .A2(new_n481), .A3(new_n470), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n477), .B1(new_n478), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n482), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n464), .A2(KEYINPUT68), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n485), .A2(new_n487), .A3(G137), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n484), .A2(KEYINPUT70), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n476), .A2(new_n483), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G160));
  NOR2_X1   g066(.A1(new_n482), .A2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G136), .ZN(new_n493));
  XOR2_X1   g068(.A(new_n493), .B(KEYINPUT71), .Z(new_n494));
  NAND2_X1  g069(.A1(new_n484), .A2(new_n475), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G112), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n467), .B1(new_n475), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(G100), .A2(G2105), .ZN(new_n499));
  XNOR2_X1  g074(.A(new_n499), .B(KEYINPUT72), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n496), .A2(G124), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n494), .A2(new_n501), .ZN(G162));
  AND2_X1   g077(.A1(new_n481), .A2(new_n470), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n504));
  AND2_X1   g079(.A1(G126), .A2(G2105), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n503), .A2(new_n504), .A3(new_n480), .A4(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n480), .A2(new_n481), .A3(new_n470), .A4(new_n505), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT73), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n485), .A2(new_n487), .A3(G138), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT4), .B1(new_n482), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT3), .B(G2104), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT4), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n474), .A2(new_n512), .A3(new_n513), .A4(G138), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  XOR2_X1   g090(.A(KEYINPUT74), .B(G114), .Z(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G2105), .ZN(new_n517));
  OAI21_X1  g092(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n509), .A2(new_n515), .A3(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(G164));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT5), .B(G543), .Z(new_n524));
  INV_X1    g099(.A(G62), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT5), .B(G543), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT6), .B(G651), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n526), .A2(G651), .B1(new_n529), .B2(G88), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n528), .A2(G50), .A3(G543), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n528), .A2(KEYINPUT75), .A3(G50), .A4(G543), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n530), .A2(new_n531), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n531), .B1(new_n530), .B2(new_n536), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(G303));
  INV_X1    g114(.A(G303), .ZN(G166));
  NAND2_X1  g115(.A1(new_n528), .A2(G89), .ZN(new_n541));
  INV_X1    g116(.A(G63), .ZN(new_n542));
  INV_X1    g117(.A(G651), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(new_n527), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT77), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT7), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n528), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G51), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n547), .A2(new_n548), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n545), .A2(new_n549), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(G168));
  NAND2_X1  g130(.A1(new_n527), .A2(new_n528), .ZN(new_n556));
  INV_X1    g131(.A(G90), .ZN(new_n557));
  INV_X1    g132(.A(G52), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n556), .A2(new_n557), .B1(new_n550), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n543), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n559), .A2(new_n561), .ZN(G171));
  INV_X1    g137(.A(G81), .ZN(new_n563));
  INV_X1    g138(.A(G43), .ZN(new_n564));
  OAI22_X1  g139(.A1(new_n556), .A2(new_n563), .B1(new_n550), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n527), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n566), .A2(new_n543), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT78), .ZN(G153));
  NAND4_X1  g145(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND4_X1  g148(.A1(G319), .A2(G483), .A3(G661), .A4(new_n573), .ZN(G188));
  NAND3_X1  g149(.A1(new_n528), .A2(G53), .A3(G543), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT79), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n529), .A2(G91), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n527), .B(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n579), .B1(new_n582), .B2(new_n543), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n578), .A2(new_n583), .ZN(G299));
  INV_X1    g159(.A(G171), .ZN(G301));
  XNOR2_X1  g160(.A(new_n554), .B(KEYINPUT81), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G286));
  NAND2_X1  g162(.A1(new_n551), .A2(G49), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n529), .A2(G87), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G288));
  INV_X1    g166(.A(G86), .ZN(new_n592));
  INV_X1    g167(.A(G48), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n556), .A2(new_n592), .B1(new_n550), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n527), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n595), .A2(new_n543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n594), .A2(new_n596), .ZN(G305));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  INV_X1    g173(.A(G47), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n556), .A2(new_n598), .B1(new_n550), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n527), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT82), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n581), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n543), .B1(new_n607), .B2(KEYINPUT83), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(KEYINPUT83), .B2(new_n607), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n529), .A2(KEYINPUT10), .A3(G92), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n556), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n610), .A2(new_n613), .B1(G54), .B2(new_n551), .ZN(new_n614));
  AND2_X1   g189(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n606), .B1(new_n615), .B2(G868), .ZN(G284));
  OAI21_X1  g191(.A(new_n606), .B1(new_n615), .B2(G868), .ZN(G321));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  MUX2_X1   g193(.A(G286), .B(G299), .S(new_n618), .Z(G297));
  MUX2_X1   g194(.A(G286), .B(G299), .S(new_n618), .Z(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n615), .B1(new_n621), .B2(G860), .ZN(G148));
  NAND2_X1  g197(.A1(new_n615), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n568), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g201(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n492), .A2(G135), .ZN(new_n631));
  OAI221_X1 g206(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n474), .C2(G111), .ZN(new_n632));
  INV_X1    g207(.A(G123), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n631), .B(new_n632), .C1(new_n495), .C2(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n634), .A2(G2096), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(G2096), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n630), .A2(new_n635), .A3(new_n636), .ZN(G156));
  INV_X1    g212(.A(KEYINPUT14), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n641), .B2(new_n640), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n643), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  AND3_X1   g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(KEYINPUT84), .B(KEYINPUT18), .Z(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  INV_X1    g235(.A(new_n653), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n660), .B1(new_n656), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2096), .B(G2100), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(new_n670), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT20), .Z(new_n674));
  AOI211_X1 g249(.A(new_n672), .B(new_n674), .C1(new_n667), .C2(new_n671), .ZN(new_n675));
  XOR2_X1   g250(.A(G1981), .B(G1986), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT86), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT85), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(G229));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G6), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n594), .A2(new_n596), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(new_n686), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT88), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT32), .B(G1981), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n684), .A2(G22), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G166), .B2(new_n684), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n690), .B1(G1971), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n684), .A2(G23), .ZN(new_n694));
  INV_X1    g269(.A(G288), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n694), .B1(new_n695), .B2(new_n684), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT33), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1976), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n693), .B(new_n698), .C1(G1971), .C2(new_n692), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n699), .A2(KEYINPUT34), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n492), .A2(G131), .ZN(new_n701));
  OAI221_X1 g276(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n474), .C2(G107), .ZN(new_n702));
  INV_X1    g277(.A(G119), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n701), .B(new_n702), .C1(new_n495), .C2(new_n703), .ZN(new_n704));
  MUX2_X1   g279(.A(G25), .B(new_n704), .S(G29), .Z(new_n705));
  XOR2_X1   g280(.A(KEYINPUT35), .B(G1991), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n707), .A2(KEYINPUT87), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(KEYINPUT87), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n684), .A2(G24), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n603), .B2(new_n684), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G1986), .ZN(new_n712));
  NOR3_X1   g287(.A1(new_n708), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n699), .B2(KEYINPUT34), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n700), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT36), .ZN(new_n716));
  NOR2_X1   g291(.A1(G168), .A2(new_n684), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n684), .B2(G21), .ZN(new_n718));
  INV_X1    g293(.A(G1966), .ZN(new_n719));
  INV_X1    g294(.A(G2072), .ZN(new_n720));
  OR2_X1    g295(.A1(G29), .A2(G33), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT25), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n492), .A2(G139), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n512), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n724), .B(new_n725), .C1(new_n474), .C2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n721), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n718), .A2(new_n719), .B1(new_n720), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n720), .B2(new_n729), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT31), .B(G11), .Z(new_n732));
  XOR2_X1   g307(.A(KEYINPUT93), .B(G28), .Z(new_n733));
  OR2_X1    g308(.A1(new_n733), .A2(KEYINPUT30), .ZN(new_n734));
  AOI21_X1  g309(.A(G29), .B1(new_n733), .B2(KEYINPUT30), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n732), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI221_X1 g311(.A(new_n736), .B1(new_n728), .B2(new_n634), .C1(new_n718), .C2(new_n719), .ZN(new_n737));
  NOR2_X1   g312(.A1(G16), .A2(G19), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n568), .B2(G16), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1341), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n684), .A2(G5), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G171), .B2(new_n684), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1961), .ZN(new_n743));
  NOR4_X1   g318(.A1(new_n731), .A2(new_n737), .A3(new_n740), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n728), .A2(G26), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT89), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT28), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n492), .A2(G140), .ZN(new_n748));
  OAI221_X1 g323(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n474), .C2(G116), .ZN(new_n749));
  INV_X1    g324(.A(G128), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n748), .B(new_n749), .C1(new_n495), .C2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n747), .B1(new_n751), .B2(G29), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT90), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G2067), .ZN(new_n754));
  NOR2_X1   g329(.A1(G164), .A2(new_n728), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G27), .B2(new_n728), .ZN(new_n756));
  INV_X1    g331(.A(G2078), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n684), .A2(G20), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT23), .Z(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G299), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT95), .B(G1956), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n758), .B(new_n759), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G34), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n766), .A2(KEYINPUT24), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(KEYINPUT24), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n728), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G160), .B2(new_n728), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2084), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n762), .B2(new_n763), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n744), .A2(new_n754), .A3(new_n765), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n728), .A2(G35), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT94), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G162), .B2(new_n728), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT29), .B(G2090), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(KEYINPUT92), .B1(G29), .B2(G32), .ZN(new_n779));
  NAND3_X1  g354(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT91), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT26), .ZN(new_n782));
  INV_X1    g357(.A(G129), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n495), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n492), .A2(G141), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(G29), .ZN(new_n789));
  MUX2_X1   g364(.A(KEYINPUT92), .B(new_n779), .S(new_n789), .Z(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT27), .B(G1996), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G4), .A2(G16), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n615), .B2(G16), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1348), .ZN(new_n795));
  NOR4_X1   g370(.A1(new_n773), .A2(new_n778), .A3(new_n792), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT96), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n716), .A2(new_n797), .ZN(G311));
  INV_X1    g373(.A(G311), .ZN(G150));
  NAND2_X1  g374(.A1(G80), .A2(G543), .ZN(new_n800));
  INV_X1    g375(.A(G67), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n524), .B2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT97), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n543), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n803), .B2(new_n802), .ZN(new_n805));
  AOI22_X1  g380(.A1(G55), .A2(new_n551), .B1(new_n529), .B2(G93), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n568), .B1(new_n807), .B2(KEYINPUT98), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(KEYINPUT98), .B2(new_n807), .ZN(new_n809));
  INV_X1    g384(.A(new_n568), .ZN(new_n810));
  OR3_X1    g385(.A1(new_n807), .A2(KEYINPUT98), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT38), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n615), .A2(G559), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n815), .A2(KEYINPUT39), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(KEYINPUT39), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n816), .A2(new_n817), .A3(G860), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n807), .A2(G860), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT37), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n818), .A2(new_n820), .ZN(G145));
  NAND2_X1  g396(.A1(new_n727), .A2(KEYINPUT99), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(new_n788), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(new_n751), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(new_n521), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n492), .A2(G142), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT100), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n496), .A2(G130), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n474), .A2(G118), .ZN(new_n829));
  OAI21_X1  g404(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n827), .B(new_n828), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n704), .B(new_n628), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT101), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n825), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n634), .B(new_n490), .ZN(new_n836));
  XNOR2_X1  g411(.A(G162), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n825), .A2(new_n833), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n835), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(G37), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n825), .A2(new_n834), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n837), .B1(new_n835), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT40), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(G395));
  NAND2_X1  g421(.A1(new_n807), .A2(new_n618), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n812), .B(new_n623), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n614), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n578), .A2(new_n583), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n850), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n848), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n853), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT41), .ZN(new_n857));
  NOR3_X1   g432(.A1(new_n856), .A2(new_n857), .A3(new_n851), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT102), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n853), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n849), .A2(KEYINPUT102), .A3(new_n850), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(new_n852), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n858), .B1(new_n857), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n855), .B1(new_n863), .B2(new_n848), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT103), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(G303), .B(new_n695), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n686), .B(new_n603), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT42), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(new_n864), .B2(new_n865), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n866), .B(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n847), .B1(new_n872), .B2(new_n618), .ZN(G295));
  OAI21_X1  g448(.A(new_n847), .B1(new_n872), .B2(new_n618), .ZN(G331));
  NOR2_X1   g449(.A1(G168), .A2(G171), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(new_n586), .B2(G171), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n812), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n812), .A2(new_n876), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n863), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n854), .B1(new_n877), .B2(new_n878), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n869), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(G37), .B1(new_n886), .B2(KEYINPUT104), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n853), .B(new_n852), .C1(new_n879), .C2(new_n857), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n862), .A2(new_n877), .A3(KEYINPUT41), .A4(new_n878), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n869), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n888), .A2(KEYINPUT105), .A3(new_n869), .A4(new_n889), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n884), .A2(new_n895), .A3(new_n885), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n887), .A2(new_n894), .A3(KEYINPUT43), .A4(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n882), .B1(new_n863), .B2(new_n880), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT104), .B1(new_n898), .B2(new_n869), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n869), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n896), .A2(new_n899), .A3(new_n840), .A4(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n897), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT44), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n887), .A2(new_n894), .A3(new_n902), .A4(new_n896), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n901), .A2(KEYINPUT43), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n905), .A2(new_n910), .ZN(G397));
  INV_X1    g486(.A(G1384), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n507), .A2(KEYINPUT73), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n507), .A2(KEYINPUT73), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n520), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n468), .A2(new_n470), .A3(new_n513), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n510), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n503), .A2(G138), .A3(new_n480), .A4(new_n474), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n917), .B1(new_n918), .B2(KEYINPUT4), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n912), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT45), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n476), .A2(G40), .A3(new_n489), .A4(new_n483), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(G1996), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n788), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n928), .A2(KEYINPUT107), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(KEYINPUT107), .ZN(new_n930));
  INV_X1    g505(.A(G2067), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n751), .B(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(new_n925), .B2(new_n788), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n929), .A2(new_n930), .B1(new_n924), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n706), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n704), .A2(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n704), .A2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n924), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G1986), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n603), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g516(.A(new_n941), .B(KEYINPUT106), .Z(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(new_n940), .B2(new_n603), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n924), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n939), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n521), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n923), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT50), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n951), .B1(new_n521), .B2(new_n912), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n950), .A2(G2084), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n921), .A2(G1384), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n923), .B1(new_n521), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(G1966), .B1(new_n922), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(G8), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n554), .A2(KEYINPUT119), .A3(G8), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT119), .B1(new_n554), .B2(G8), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT51), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n957), .A2(new_n963), .A3(KEYINPUT122), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT122), .ZN(new_n965));
  INV_X1    g540(.A(G8), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n954), .B1(new_n915), .B2(new_n919), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n949), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT45), .B1(new_n521), .B2(new_n912), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n719), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n920), .A2(KEYINPUT50), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n923), .B1(new_n521), .B2(new_n947), .ZN(new_n972));
  INV_X1    g547(.A(G2084), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n966), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n965), .B1(new_n975), .B2(new_n962), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n964), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT121), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n960), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  AOI211_X1 g554(.A(KEYINPUT121), .B(new_n966), .C1(new_n970), .C2(new_n974), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT51), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n970), .A2(new_n974), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n958), .A2(new_n959), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n983), .A2(KEYINPUT120), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT120), .B1(new_n983), .B2(new_n984), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT123), .B1(new_n982), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT123), .ZN(new_n990));
  AOI211_X1 g565(.A(new_n990), .B(new_n987), .C1(new_n977), .C2(new_n981), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT62), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n984), .B1(new_n957), .B2(KEYINPUT121), .ZN(new_n993));
  INV_X1    g568(.A(new_n980), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n961), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n964), .A2(new_n976), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n988), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n990), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT62), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n982), .A2(KEYINPUT123), .A3(new_n988), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(G303), .A2(KEYINPUT109), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n530), .A2(new_n536), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT76), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n530), .A2(new_n531), .A3(new_n536), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1004), .A2(new_n1005), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1004), .A2(G8), .A3(new_n1005), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1002), .A2(new_n1008), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G2090), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n971), .A2(new_n972), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1971), .B1(new_n922), .B2(new_n955), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1014), .B1(new_n1015), .B2(KEYINPUT108), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n506), .A2(new_n508), .B1(new_n517), .B2(new_n519), .ZN(new_n1017));
  AOI21_X1  g592(.A(G1384), .B1(new_n1017), .B2(new_n515), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n967), .B(new_n949), .C1(new_n1018), .C2(KEYINPUT45), .ZN(new_n1019));
  INV_X1    g594(.A(G1971), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1019), .A2(KEYINPUT108), .A3(new_n1020), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1012), .B(G8), .C1(new_n1016), .C2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT49), .ZN(new_n1024));
  INV_X1    g599(.A(G1981), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n686), .A2(new_n1025), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n594), .A2(new_n596), .A3(G1981), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1023), .B(new_n1024), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(G305), .A2(G1981), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1027), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1018), .A2(new_n949), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1028), .A2(new_n1032), .A3(G8), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n695), .A2(G1976), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(G8), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT52), .ZN(new_n1037));
  INV_X1    g612(.A(G1976), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT52), .B1(G288), .B2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1033), .A2(G8), .A3(new_n1035), .A4(new_n1039), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1034), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1022), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1020), .B1(new_n968), .B2(new_n969), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n1014), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n966), .B1(new_n1044), .B2(KEYINPUT112), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1043), .A2(new_n1046), .A3(new_n1014), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1012), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n968), .A2(new_n969), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT53), .B1(new_n1049), .B2(new_n757), .ZN(new_n1050));
  INV_X1    g625(.A(G1961), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1051), .B1(new_n950), .B2(new_n952), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n922), .A2(new_n955), .A3(KEYINPUT53), .A4(new_n757), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(G171), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1042), .A2(new_n1048), .A3(new_n1055), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n992), .A2(new_n1001), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1034), .A2(new_n1038), .A3(new_n695), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n1030), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT111), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(KEYINPUT111), .A3(new_n1030), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1061), .A2(G8), .A3(new_n1033), .A4(new_n1062), .ZN(new_n1063));
  OR2_X1    g638(.A1(new_n1016), .A2(new_n1021), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1064), .A2(G8), .A3(new_n1012), .A4(new_n1041), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1042), .A2(new_n1048), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n975), .A2(KEYINPUT113), .A3(new_n586), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT113), .B1(new_n975), .B2(new_n586), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT63), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT63), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1012), .B1(new_n1064), .B2(G8), .ZN(new_n1075));
  OR3_X1    g650(.A1(new_n1074), .A2(new_n1075), .A3(new_n1042), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1066), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  XOR2_X1   g652(.A(KEYINPUT56), .B(G2072), .Z(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT115), .B1(new_n1019), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1078), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n922), .A2(new_n955), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT114), .B(G1956), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n950), .B2(new_n952), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n583), .A2(KEYINPUT57), .A3(new_n577), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1087), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1088));
  AOI21_X1  g663(.A(G1348), .B1(new_n971), .B2(new_n972), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1018), .A2(new_n949), .A3(new_n931), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  OAI22_X1  g667(.A1(new_n1086), .A2(new_n1088), .B1(new_n849), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1083), .A2(new_n1088), .A3(new_n1085), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1092), .A2(KEYINPUT60), .ZN(new_n1096));
  INV_X1    g671(.A(G1348), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n950), .B2(new_n952), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(KEYINPUT60), .A3(new_n1090), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(KEYINPUT118), .A3(new_n615), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT118), .B1(new_n1099), .B2(new_n615), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1098), .A2(new_n849), .A3(KEYINPUT60), .A4(new_n1090), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1104), .B(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1096), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1094), .A2(KEYINPUT61), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT61), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1083), .A2(new_n1088), .A3(new_n1109), .A4(new_n1085), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n810), .A2(KEYINPUT116), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n922), .A2(new_n955), .A3(new_n925), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT58), .B(G1341), .Z(new_n1113));
  NAND2_X1  g688(.A1(new_n1033), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1111), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1108), .A2(new_n1110), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1095), .B1(new_n1107), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(new_n1019), .B2(G2078), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1121), .A2(G301), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1055), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1123), .A2(KEYINPUT124), .A3(new_n1124), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1055), .A2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(KEYINPUT125), .B(G171), .C1(new_n1050), .C2(new_n1054), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1131), .A2(KEYINPUT54), .A3(new_n1122), .A4(new_n1132), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1067), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1119), .A2(new_n1129), .A3(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n989), .A2(new_n991), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1077), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n946), .B1(new_n1057), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT127), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n751), .A2(G2067), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n934), .B2(new_n936), .ZN(new_n1141));
  INV_X1    g716(.A(new_n924), .ZN(new_n1142));
  OR3_X1    g717(.A1(new_n1141), .A2(KEYINPUT126), .A3(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT126), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1144));
  INV_X1    g719(.A(new_n932), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n924), .B1(new_n1145), .B2(new_n927), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n926), .A2(KEYINPUT46), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n926), .A2(KEYINPUT46), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  XOR2_X1   g724(.A(new_n1149), .B(KEYINPUT47), .Z(new_n1150));
  NOR2_X1   g725(.A1(new_n1142), .A2(new_n942), .ZN(new_n1151));
  XOR2_X1   g726(.A(new_n1151), .B(KEYINPUT48), .Z(new_n1152));
  AOI21_X1  g727(.A(new_n1150), .B1(new_n939), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1143), .A2(new_n1144), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1138), .A2(new_n1139), .A3(new_n1155), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT63), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1074), .A2(new_n1075), .A3(new_n1042), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1108), .A2(new_n1110), .A3(new_n1117), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT118), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT60), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1089), .A2(new_n1091), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1162), .B1(new_n1164), .B2(new_n849), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1164), .A2(new_n1105), .A3(new_n849), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1104), .A2(KEYINPUT117), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .A4(new_n1100), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1096), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g745(.A1(new_n1161), .A2(new_n1170), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1127), .A2(new_n1128), .A3(new_n1133), .A4(new_n1067), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n998), .A2(new_n1000), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1160), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n992), .A2(new_n1001), .A3(new_n1056), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n945), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(KEYINPUT127), .B1(new_n1177), .B2(new_n1154), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1156), .A2(new_n1178), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g754(.A(new_n844), .ZN(new_n1181));
  NOR4_X1   g755(.A1(G229), .A2(new_n462), .A3(G401), .A4(G227), .ZN(new_n1182));
  AND3_X1   g756(.A1(new_n1181), .A2(new_n908), .A3(new_n1182), .ZN(G308));
  NAND3_X1  g757(.A1(new_n1181), .A2(new_n908), .A3(new_n1182), .ZN(G225));
endmodule


