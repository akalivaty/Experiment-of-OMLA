//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984, new_n985;
  XNOR2_X1  g000(.A(KEYINPUT96), .B(G64gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G57gat), .ZN(new_n203));
  INV_X1    g002(.A(G64gat), .ZN(new_n204));
  OAI211_X1 g003(.A(new_n203), .B(KEYINPUT97), .C1(G57gat), .C2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G71gat), .A2(G78gat), .ZN(new_n206));
  OR2_X1    g005(.A1(G71gat), .A2(G78gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT9), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n205), .B(new_n209), .C1(KEYINPUT97), .C2(new_n203), .ZN(new_n210));
  XNOR2_X1  g009(.A(G57gat), .B(G64gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n206), .B(new_n207), .C1(new_n211), .C2(new_n208), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT21), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G231gat), .A2(G233gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G127gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G8gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(G15gat), .B(G22gat), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n221), .A2(G1gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n220), .B1(new_n222), .B2(KEYINPUT94), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n221), .B1(new_n224), .B2(G1gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n223), .A2(new_n226), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n227), .B(new_n228), .C1(new_n213), .C2(new_n214), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n219), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n231));
  INV_X1    g030(.A(G155gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(G183gat), .B(G211gat), .Z(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n230), .A2(new_n235), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT93), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n239), .B1(G29gat), .B2(G36gat), .ZN(new_n240));
  INV_X1    g039(.A(G29gat), .ZN(new_n241));
  INV_X1    g040(.A(G36gat), .ZN(new_n242));
  NOR3_X1   g041(.A1(new_n241), .A2(new_n242), .A3(KEYINPUT93), .ZN(new_n243));
  XNOR2_X1  g042(.A(G43gat), .B(G50gat), .ZN(new_n244));
  AOI211_X1 g043(.A(new_n240), .B(new_n243), .C1(KEYINPUT15), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n241), .A2(new_n242), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT14), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n245), .B(new_n247), .C1(KEYINPUT15), .C2(new_n244), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n247), .B1(new_n241), .B2(new_n242), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(KEYINPUT15), .A3(new_n244), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT17), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n248), .A2(KEYINPUT17), .A3(new_n250), .ZN(new_n254));
  NAND2_X1  g053(.A1(G99gat), .A2(G106gat), .ZN(new_n255));
  INV_X1    g054(.A(G85gat), .ZN(new_n256));
  INV_X1    g055(.A(G92gat), .ZN(new_n257));
  AOI22_X1  g056(.A1(KEYINPUT8), .A2(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(new_n256), .B2(new_n257), .ZN(new_n260));
  NAND4_X1  g059(.A1(KEYINPUT100), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G99gat), .B(G106gat), .Z(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n253), .A2(new_n254), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G232gat), .A2(G233gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT98), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT41), .ZN(new_n268));
  XOR2_X1   g067(.A(G190gat), .B(G218gat), .Z(new_n269));
  INV_X1    g068(.A(KEYINPUT101), .ZN(new_n270));
  OAI22_X1  g069(.A1(new_n267), .A2(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n264), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n271), .B1(new_n251), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n265), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n269), .A2(new_n270), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n274), .B(new_n275), .Z(new_n276));
  NAND2_X1  g075(.A1(new_n267), .A2(new_n268), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n277), .B(KEYINPUT99), .Z(new_n278));
  XOR2_X1   g077(.A(G134gat), .B(G162gat), .Z(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT102), .ZN(new_n281));
  OR2_X1    g080(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  OR2_X1    g081(.A1(new_n280), .A2(KEYINPUT102), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n276), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G230gat), .ZN(new_n286));
  INV_X1    g085(.A(G233gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n213), .B(new_n272), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n290), .A2(KEYINPUT10), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n272), .A2(KEYINPUT10), .A3(new_n210), .A4(new_n212), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n288), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n290), .A2(new_n288), .ZN(new_n295));
  XNOR2_X1  g094(.A(G120gat), .B(G148gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(G176gat), .B(G204gat), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n296), .B(new_n297), .Z(new_n298));
  NAND3_X1  g097(.A1(new_n294), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n298), .ZN(new_n300));
  INV_X1    g099(.A(new_n295), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n300), .B1(new_n293), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n238), .A2(new_n285), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT95), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n227), .A2(new_n228), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n307), .B1(new_n252), .B2(new_n251), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n308), .A2(new_n254), .B1(new_n307), .B2(new_n251), .ZN(new_n309));
  NAND2_X1  g108(.A1(G229gat), .A2(G233gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT18), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n309), .A2(KEYINPUT18), .A3(new_n310), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n307), .B(new_n251), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n310), .B(KEYINPUT13), .Z(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n313), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G113gat), .B(G141gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(G169gat), .B(G197gat), .Z(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(KEYINPUT12), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n318), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n313), .A2(new_n314), .A3(new_n317), .A4(new_n324), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT36), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(G169gat), .A2(G176gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT67), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT64), .ZN(new_n335));
  INV_X1    g134(.A(G169gat), .ZN(new_n336));
  INV_X1    g135(.A(G176gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT26), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n330), .A2(KEYINPUT67), .A3(new_n331), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n334), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G183gat), .A2(G190gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n346));
  INV_X1    g145(.A(G183gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT27), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT27), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G183gat), .ZN(new_n350));
  INV_X1    g149(.A(G190gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n348), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT27), .B(G183gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n356), .A2(new_n351), .A3(new_n353), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n346), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n345), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT23), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(G169gat), .B2(G176gat), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n361), .A2(KEYINPUT25), .A3(new_n331), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n338), .A2(new_n340), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n362), .B1(new_n363), .B2(KEYINPUT23), .ZN(new_n364));
  NOR2_X1   g163(.A1(G183gat), .A2(G190gat), .ZN(new_n365));
  AND2_X1   g164(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n365), .B1(new_n366), .B2(G190gat), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(KEYINPUT65), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT24), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n344), .A2(KEYINPUT65), .A3(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n367), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n344), .A2(new_n370), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n347), .A2(new_n351), .ZN(new_n374));
  NAND3_X1  g173(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT23), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n376), .A2(new_n361), .A3(new_n331), .A4(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT25), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n364), .A2(new_n372), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AND2_X1   g179(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n382));
  OAI21_X1  g181(.A(G134gat), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT68), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n218), .ZN(new_n385));
  INV_X1    g184(.A(G134gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G113gat), .B(G120gat), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n383), .B(new_n388), .C1(KEYINPUT1), .C2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G113gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(G120gat), .ZN(new_n392));
  INV_X1    g191(.A(G120gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(G113gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n392), .A2(new_n394), .A3(KEYINPUT69), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT1), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT69), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n397), .A2(new_n391), .A3(G120gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(G127gat), .B(G134gat), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n395), .A2(new_n396), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT70), .B1(new_n390), .B2(new_n400), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n390), .A2(KEYINPUT70), .A3(new_n400), .ZN(new_n402));
  OAI22_X1  g201(.A1(new_n359), .A2(new_n380), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n353), .B1(new_n356), .B2(new_n351), .ZN(new_n404));
  AND4_X1   g203(.A1(new_n351), .A2(new_n348), .A3(new_n350), .A4(new_n353), .ZN(new_n405));
  OAI22_X1  g204(.A1(new_n404), .A2(new_n405), .B1(KEYINPUT66), .B2(KEYINPUT28), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n406), .A2(new_n344), .A3(new_n343), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n400), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT70), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n377), .A2(new_n361), .A3(new_n331), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n379), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n374), .A2(new_n375), .ZN(new_n414));
  INV_X1    g213(.A(new_n369), .ZN(new_n415));
  INV_X1    g214(.A(new_n371), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n362), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n338), .A2(KEYINPUT23), .A3(new_n340), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n413), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n390), .A2(new_n400), .A3(KEYINPUT70), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n407), .A2(new_n410), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n403), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G227gat), .A2(G233gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT33), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(KEYINPUT71), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n427), .A2(KEYINPUT32), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT71), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n425), .B1(new_n403), .B2(new_n423), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n431), .B1(new_n432), .B2(KEYINPUT33), .ZN(new_n433));
  XOR2_X1   g232(.A(G15gat), .B(G43gat), .Z(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(KEYINPUT72), .ZN(new_n435));
  XNOR2_X1  g234(.A(G71gat), .B(G99gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n429), .A2(new_n430), .A3(new_n433), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(KEYINPUT33), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n427), .A2(KEYINPUT32), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n403), .A2(new_n423), .A3(new_n425), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT73), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n443), .B1(new_n441), .B2(new_n442), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n438), .A2(new_n440), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n446), .B1(new_n438), .B2(new_n440), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n329), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT76), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g250(.A(KEYINPUT76), .B(new_n329), .C1(new_n447), .C2(new_n448), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n438), .A2(new_n440), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT75), .B1(new_n444), .B2(new_n445), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n441), .A2(new_n442), .ZN(new_n455));
  INV_X1    g254(.A(new_n443), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT75), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n453), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n438), .A2(new_n440), .A3(new_n446), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(KEYINPUT36), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n451), .A2(new_n452), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(G141gat), .ZN(new_n466));
  INV_X1    g265(.A(G148gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(G141gat), .A2(G148gat), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(G162gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(G155gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n232), .A2(G162gat), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(KEYINPUT83), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT83), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(G162gat), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n232), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT2), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n470), .B(new_n474), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n468), .A2(new_n479), .A3(new_n469), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n472), .A2(new_n473), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  XOR2_X1   g283(.A(G211gat), .B(G218gat), .Z(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT77), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n488));
  OR2_X1    g287(.A1(G197gat), .A2(G204gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(G197gat), .A2(G204gat), .ZN(new_n490));
  AOI211_X1 g289(.A(new_n487), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n490), .ZN(new_n492));
  INV_X1    g291(.A(new_n488), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT77), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n486), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n492), .A2(KEYINPUT77), .A3(new_n493), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n485), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT29), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n484), .B1(new_n498), .B2(KEYINPUT3), .ZN(new_n499));
  XOR2_X1   g298(.A(G197gat), .B(G204gat), .Z(new_n500));
  OAI21_X1  g299(.A(new_n487), .B1(new_n500), .B2(new_n488), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n485), .B1(new_n501), .B2(new_n496), .ZN(new_n502));
  INV_X1    g301(.A(new_n497), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT78), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(KEYINPUT79), .B(KEYINPUT29), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n484), .B2(KEYINPUT3), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT78), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n495), .A2(new_n507), .A3(new_n497), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n504), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G228gat), .A2(G233gat), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n499), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n505), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n513), .B1(new_n495), .B2(new_n497), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n484), .B1(new_n514), .B2(KEYINPUT3), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n495), .A2(new_n497), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n506), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n511), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(G22gat), .B1(new_n512), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT86), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT83), .B(G162gat), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT2), .B1(new_n522), .B2(new_n232), .ZN(new_n523));
  AND4_X1   g322(.A1(new_n468), .A2(new_n472), .A3(new_n473), .A4(new_n469), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n523), .A2(new_n524), .B1(new_n481), .B2(new_n482), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n505), .B1(new_n502), .B2(new_n503), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT3), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n513), .B1(new_n525), .B2(new_n527), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n529), .A2(new_n516), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n510), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G22gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n499), .A2(new_n509), .A3(new_n511), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G78gat), .B(G106gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT31), .B(G50gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n520), .A2(new_n521), .A3(new_n534), .A4(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n534), .A2(KEYINPUT86), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n540), .A2(new_n537), .B1(new_n520), .B2(new_n534), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT5), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n484), .A2(new_n408), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n480), .A2(new_n483), .A3(new_n390), .A4(new_n400), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G225gat), .A2(G233gat), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n543), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n525), .A2(new_n527), .B1(new_n400), .B2(new_n390), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT84), .B1(new_n525), .B2(new_n527), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT84), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n484), .A2(new_n552), .A3(KEYINPUT3), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n410), .A2(KEYINPUT4), .A3(new_n525), .A4(new_n422), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT4), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n548), .B1(new_n545), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n549), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n410), .A2(new_n422), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n556), .B1(new_n560), .B2(new_n484), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n545), .A2(new_n556), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n548), .A2(KEYINPUT5), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(G1gat), .B(G29gat), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT0), .ZN(new_n568));
  XNOR2_X1  g367(.A(G57gat), .B(G85gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT6), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n559), .A2(new_n565), .A3(new_n570), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT85), .ZN(new_n576));
  AND4_X1   g375(.A1(new_n576), .A2(new_n566), .A3(KEYINPUT6), .A4(new_n571), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n570), .B1(new_n559), .B2(new_n565), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n576), .B1(new_n578), .B2(KEYINPUT6), .ZN(new_n579));
  NOR3_X1   g378(.A1(new_n575), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G226gat), .A2(G233gat), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n330), .A2(KEYINPUT67), .A3(new_n331), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT67), .B1(new_n330), .B2(new_n331), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n584), .A2(new_n341), .B1(G183gat), .B2(G190gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n372), .A2(new_n419), .A3(new_n418), .ZN(new_n586));
  AOI22_X1  g385(.A1(new_n585), .A2(new_n406), .B1(new_n586), .B2(new_n413), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n581), .B1(new_n587), .B2(KEYINPUT29), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n588), .B(new_n516), .C1(new_n581), .C2(new_n587), .ZN(new_n589));
  XOR2_X1   g388(.A(G8gat), .B(G36gat), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT81), .ZN(new_n591));
  XNOR2_X1  g390(.A(G64gat), .B(G92gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT80), .B1(new_n587), .B2(new_n581), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT80), .ZN(new_n595));
  INV_X1    g394(.A(new_n581), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n595), .B(new_n596), .C1(new_n359), .C2(new_n380), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n505), .B1(new_n359), .B2(new_n380), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n594), .A2(new_n597), .B1(new_n581), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n504), .A2(new_n508), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n589), .B(new_n593), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT82), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT30), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT30), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n601), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n594), .A2(new_n597), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n598), .A2(new_n581), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n600), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(new_n589), .ZN(new_n612));
  INV_X1    g411(.A(new_n593), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n604), .A2(new_n606), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n542), .B1(new_n580), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n465), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT87), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n465), .A2(KEYINPUT87), .A3(new_n616), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT88), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n572), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n578), .A2(KEYINPUT88), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n548), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n544), .A2(new_n547), .A3(new_n545), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n626), .A2(KEYINPUT39), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT39), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n625), .A2(new_n629), .A3(new_n548), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n570), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT40), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n626), .A2(KEYINPUT39), .A3(new_n627), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n633), .A2(new_n634), .A3(new_n570), .A4(new_n630), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n615), .A2(new_n624), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n540), .A2(new_n537), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n520), .A2(new_n534), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n538), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n577), .A2(new_n579), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n574), .A2(new_n573), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n622), .A2(new_n643), .A3(new_n623), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(new_n644), .A3(new_n601), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n407), .A2(new_n421), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT29), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n596), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n587), .A2(new_n581), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n517), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT89), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT89), .ZN(new_n652));
  OAI211_X1 g451(.A(new_n652), .B(new_n517), .C1(new_n648), .C2(new_n649), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n651), .B(new_n653), .C1(new_n610), .C2(new_n609), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT37), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT37), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n656), .B(new_n589), .C1(new_n599), .C2(new_n600), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n613), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT38), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n655), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n656), .B1(new_n611), .B2(new_n589), .ZN(new_n662));
  OAI21_X1  g461(.A(KEYINPUT38), .B1(new_n662), .B2(new_n658), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n637), .B(new_n641), .C1(new_n645), .C2(new_n664), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n619), .A2(new_n620), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT35), .B1(new_n642), .B2(new_n644), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n604), .A2(new_n606), .A3(new_n614), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n447), .A2(new_n448), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .A4(new_n641), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT90), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n542), .A2(new_n447), .A3(new_n448), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n673), .A2(KEYINPUT90), .A3(new_n668), .A4(new_n667), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT91), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n454), .A2(new_n460), .ZN(new_n676));
  INV_X1    g475(.A(new_n440), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n432), .A2(new_n431), .A3(KEYINPUT33), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT32), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n437), .B1(new_n432), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n677), .B1(new_n681), .B2(new_n433), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n463), .B1(new_n676), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n675), .B1(new_n683), .B2(new_n542), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n580), .A2(new_n615), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n641), .A2(KEYINPUT91), .A3(new_n463), .A4(new_n462), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n672), .A2(new_n674), .B1(new_n687), .B2(KEYINPUT35), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n306), .B(new_n328), .C1(new_n666), .C2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n665), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n690), .B1(new_n617), .B2(new_n618), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n688), .B1(new_n691), .B2(new_n620), .ZN(new_n692));
  INV_X1    g491(.A(new_n328), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT95), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n305), .B1(new_n689), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n580), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT103), .B(G1gat), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1324gat));
  AND2_X1   g497(.A1(new_n695), .A2(new_n615), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT16), .B(G8gat), .Z(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n699), .A2(new_n220), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT42), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(G1325gat));
  INV_X1    g506(.A(G15gat), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n695), .A2(new_n708), .A3(new_n669), .ZN(new_n709));
  INV_X1    g508(.A(new_n465), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n695), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n711), .B2(new_n708), .ZN(G1326gat));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n542), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT43), .B(G22gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1327gat));
  NOR3_X1   g514(.A1(new_n238), .A2(new_n285), .A3(new_n303), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(new_n689), .B2(new_n694), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n718), .A2(new_n241), .A3(new_n580), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(KEYINPUT45), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n719), .A2(KEYINPUT45), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722));
  INV_X1    g521(.A(new_n285), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n465), .A2(new_n665), .A3(new_n616), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n722), .B(new_n723), .C1(new_n688), .C2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n672), .A2(new_n674), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n687), .A2(KEYINPUT35), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n465), .A2(new_n665), .A3(new_n616), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n732), .A2(KEYINPUT105), .A3(new_n722), .A4(new_n723), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n727), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(KEYINPUT44), .B1(new_n692), .B2(new_n285), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n238), .B(KEYINPUT104), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n737), .A2(new_n693), .A3(new_n303), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n580), .ZN(new_n740));
  OAI21_X1  g539(.A(G29gat), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n720), .B1(new_n721), .B2(new_n741), .ZN(G1328gat));
  NAND3_X1  g541(.A1(new_n718), .A2(new_n242), .A3(new_n615), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n743), .A2(KEYINPUT46), .ZN(new_n744));
  OAI21_X1  g543(.A(G36gat), .B1(new_n739), .B2(new_n668), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(KEYINPUT46), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(G1329gat));
  NAND2_X1  g546(.A1(new_n718), .A2(new_n669), .ZN(new_n748));
  INV_X1    g547(.A(G43gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n710), .A2(G43gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n739), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT47), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT47), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n750), .B(new_n754), .C1(new_n739), .C2(new_n751), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(G1330gat));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n641), .A2(new_n757), .A3(G50gat), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT107), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n718), .A2(new_n759), .ZN(new_n760));
  AOI211_X1 g559(.A(KEYINPUT107), .B(new_n717), .C1(new_n689), .C2(new_n694), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT48), .ZN(new_n763));
  OAI211_X1 g562(.A(KEYINPUT106), .B(G50gat), .C1(new_n739), .C2(new_n641), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n763), .B1(new_n762), .B2(new_n764), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(G1331gat));
  NOR2_X1   g566(.A1(new_n304), .A2(new_n328), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(new_n238), .A3(new_n285), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT108), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n730), .B2(new_n731), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n580), .ZN(new_n772));
  XNOR2_X1  g571(.A(KEYINPUT109), .B(G57gat), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1332gat));
  INV_X1    g573(.A(KEYINPUT49), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n771), .B(new_n615), .C1(new_n775), .C2(new_n204), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n204), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1333gat));
  NAND2_X1  g577(.A1(new_n771), .A2(new_n710), .ZN(new_n779));
  INV_X1    g578(.A(new_n669), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n780), .A2(G71gat), .ZN(new_n781));
  AOI22_X1  g580(.A1(new_n779), .A2(G71gat), .B1(new_n771), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g582(.A1(new_n771), .A2(new_n542), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(G78gat), .ZN(G1335gat));
  INV_X1    g584(.A(new_n238), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n768), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n736), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(G85gat), .B1(new_n789), .B2(new_n740), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n732), .A2(new_n693), .A3(new_n786), .A4(new_n723), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n793), .A2(new_n256), .A3(new_n580), .A4(new_n303), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n790), .A2(new_n794), .ZN(G1336gat));
  XOR2_X1   g594(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n796));
  NOR3_X1   g595(.A1(new_n304), .A2(G92gat), .A3(new_n668), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n796), .B1(new_n793), .B2(new_n797), .ZN(new_n798));
  AOI211_X1 g597(.A(new_n668), .B(new_n787), .C1(new_n734), .C2(new_n735), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n257), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n736), .A2(new_n615), .A3(new_n788), .ZN(new_n801));
  XOR2_X1   g600(.A(new_n797), .B(KEYINPUT110), .Z(new_n802));
  AOI22_X1  g601(.A1(new_n801), .A2(G92gat), .B1(new_n793), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n803), .A2(KEYINPUT111), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n793), .A2(new_n802), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(new_n799), .B2(new_n257), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n806), .B1(new_n808), .B2(KEYINPUT52), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n800), .B1(new_n805), .B2(new_n809), .ZN(G1337gat));
  NOR3_X1   g609(.A1(new_n304), .A2(G99gat), .A3(new_n780), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(KEYINPUT114), .Z(new_n812));
  NAND2_X1  g611(.A1(new_n793), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n789), .A2(new_n465), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n814), .A2(KEYINPUT113), .ZN(new_n815));
  OAI21_X1  g614(.A(G99gat), .B1(new_n814), .B2(KEYINPUT113), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n813), .B1(new_n815), .B2(new_n816), .ZN(G1338gat));
  OAI21_X1  g616(.A(G106gat), .B1(new_n789), .B2(new_n641), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT115), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n641), .A2(G106gat), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n793), .A2(new_n303), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(new_n822), .A3(KEYINPUT53), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n818), .B(new_n821), .C1(KEYINPUT115), .C2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(G1339gat));
  NOR2_X1   g625(.A1(new_n305), .A2(new_n328), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n309), .A2(new_n310), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n315), .A2(new_n316), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n323), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n327), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n303), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n291), .A2(new_n292), .A3(new_n288), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n835), .A2(new_n293), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n293), .A2(new_n836), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n300), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n833), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n294), .A2(KEYINPUT54), .A3(new_n834), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n841), .A2(KEYINPUT55), .A3(new_n300), .A4(new_n838), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n840), .A2(new_n299), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n832), .B1(new_n843), .B2(new_n693), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n285), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n285), .B1(new_n831), .B2(new_n847), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n831), .A2(new_n847), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n846), .B1(new_n850), .B2(new_n843), .ZN(new_n851));
  INV_X1    g650(.A(new_n843), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n852), .A2(KEYINPUT117), .A3(new_n849), .A4(new_n848), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n845), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n737), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n827), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n684), .A2(new_n686), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n740), .A2(new_n615), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(G113gat), .B1(new_n860), .B2(new_n328), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n857), .A2(new_n673), .A3(new_n859), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n862), .A2(new_n391), .A3(new_n693), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n861), .A2(new_n863), .ZN(G1340gat));
  AOI21_X1  g663(.A(G120gat), .B1(new_n860), .B2(new_n303), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n862), .A2(new_n393), .A3(new_n304), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(G1341gat));
  NAND3_X1  g666(.A1(new_n860), .A2(new_n218), .A3(new_n238), .ZN(new_n868));
  OAI21_X1  g667(.A(G127gat), .B1(new_n862), .B2(new_n855), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1342gat));
  NOR2_X1   g669(.A1(new_n856), .A2(new_n740), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n285), .A2(G134gat), .A3(new_n615), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n858), .A3(new_n872), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT56), .Z(new_n874));
  OAI21_X1  g673(.A(G134gat), .B1(new_n862), .B2(new_n285), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1343gat));
  NAND2_X1  g675(.A1(new_n465), .A2(new_n859), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n641), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n854), .A2(new_n786), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n879), .B1(new_n880), .B2(new_n827), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n878), .B1(new_n856), .B2(new_n641), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n877), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n466), .B1(new_n883), .B2(new_n328), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n710), .A2(new_n615), .A3(new_n641), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n871), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n328), .A2(new_n466), .ZN(new_n887));
  XOR2_X1   g686(.A(new_n887), .B(KEYINPUT118), .Z(new_n888));
  AND2_X1   g687(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT58), .B1(new_n884), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT58), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n886), .A2(new_n888), .ZN(new_n892));
  AOI211_X1 g691(.A(new_n693), .B(new_n877), .C1(new_n881), .C2(new_n882), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n891), .B(new_n892), .C1(new_n893), .C2(new_n466), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n890), .A2(new_n894), .ZN(G1344gat));
  NAND3_X1  g694(.A1(new_n886), .A2(new_n467), .A3(new_n303), .ZN(new_n896));
  AOI211_X1 g695(.A(KEYINPUT59), .B(new_n467), .C1(new_n883), .C2(new_n303), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT57), .B1(new_n856), .B2(new_n641), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n852), .A2(new_n849), .A3(new_n848), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n238), .B1(new_n845), .B2(new_n900), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n878), .B(new_n542), .C1(new_n901), .C2(new_n827), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n877), .A2(KEYINPUT119), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n304), .B1(new_n877), .B2(KEYINPUT119), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n899), .A2(new_n902), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n898), .B1(new_n905), .B2(G148gat), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n896), .B1(new_n897), .B2(new_n906), .ZN(G1345gat));
  AOI21_X1  g706(.A(new_n232), .B1(new_n883), .B2(new_n737), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n871), .A2(new_n885), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n238), .A2(new_n232), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT120), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n911), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n914));
  AOI211_X1 g713(.A(new_n855), .B(new_n877), .C1(new_n881), .C2(new_n882), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n913), .B(new_n914), .C1(new_n915), .C2(new_n232), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n912), .A2(new_n916), .ZN(G1346gat));
  NAND3_X1  g716(.A1(new_n886), .A2(new_n522), .A3(new_n723), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n883), .A2(new_n723), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n522), .ZN(G1347gat));
  NOR2_X1   g719(.A1(new_n668), .A2(new_n580), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n857), .A2(new_n858), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n328), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n857), .A2(new_n673), .A3(new_n921), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n924), .A2(new_n336), .A3(new_n693), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n923), .A2(new_n925), .ZN(G1348gat));
  NOR2_X1   g725(.A1(new_n304), .A2(G176gat), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n922), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G176gat), .B1(new_n924), .B2(new_n304), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n930), .B(new_n931), .ZN(G1349gat));
  AND2_X1   g731(.A1(new_n238), .A2(new_n356), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n922), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(G183gat), .B1(new_n924), .B2(new_n855), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(KEYINPUT60), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT60), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n934), .A2(new_n935), .A3(new_n936), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1350gat));
  NAND3_X1  g740(.A1(new_n922), .A2(new_n351), .A3(new_n723), .ZN(new_n942));
  OAI21_X1  g741(.A(G190gat), .B1(new_n924), .B2(new_n285), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(G1351gat));
  NAND2_X1  g745(.A1(new_n465), .A2(new_n921), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n856), .A2(new_n641), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(G197gat), .B1(new_n948), .B2(new_n328), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n899), .A2(new_n902), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT123), .ZN(new_n951));
  INV_X1    g750(.A(new_n947), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT123), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n899), .A2(new_n953), .A3(new_n902), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n951), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n328), .A2(G197gat), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n949), .B1(new_n955), .B2(new_n956), .ZN(G1352gat));
  XOR2_X1   g756(.A(KEYINPUT124), .B(G204gat), .Z(new_n958));
  NAND3_X1  g757(.A1(new_n948), .A2(new_n303), .A3(new_n958), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n959), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n963), .B1(new_n959), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n960), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n951), .A2(new_n303), .A3(new_n952), .A4(new_n954), .ZN(new_n967));
  INV_X1    g766(.A(new_n958), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n966), .A2(new_n969), .ZN(G1353gat));
  OAI21_X1  g769(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n786), .A2(new_n947), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n972), .B1(new_n950), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n975), .A2(KEYINPUT126), .A3(KEYINPUT63), .ZN(new_n976));
  NAND2_X1  g775(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n972), .B(new_n977), .C1(new_n950), .C2(new_n974), .ZN(new_n978));
  INV_X1    g777(.A(G211gat), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n948), .A2(new_n979), .A3(new_n238), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n976), .A2(new_n978), .A3(new_n980), .ZN(G1354gat));
  NAND4_X1  g780(.A1(new_n951), .A2(new_n723), .A3(new_n952), .A4(new_n954), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(G218gat), .ZN(new_n983));
  INV_X1    g782(.A(G218gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n948), .A2(new_n984), .A3(new_n723), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n983), .A2(new_n985), .ZN(G1355gat));
endmodule


