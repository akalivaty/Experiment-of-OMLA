//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n624, new_n625,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT66), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT67), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT68), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G238), .A3(G237), .A4(G235), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT70), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT71), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT72), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT72), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n468), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AND3_X1   g051(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n477));
  INV_X1    g052(.A(G137), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n478), .B1(new_n472), .B2(new_n473), .ZN(new_n479));
  XNOR2_X1  g054(.A(KEYINPUT72), .B(G2105), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  OAI221_X1 g058(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n480), .C2(G112), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n472), .A2(new_n473), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n468), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n484), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  NOR2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(KEYINPUT73), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT73), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n486), .A2(new_n493), .A3(new_n464), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n488), .B1(G136), .B2(new_n495), .ZN(G162));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT74), .ZN(new_n499));
  OAI21_X1  g074(.A(G2105), .B1(new_n499), .B2(G114), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(KEYINPUT74), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n498), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g078(.A(G126), .B(G2105), .C1(new_n489), .C2(new_n490), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(G138), .B1(new_n489), .B2(new_n490), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT4), .B1(new_n506), .B2(new_n468), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n486), .A2(new_n480), .A3(new_n508), .A4(G138), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n505), .B1(new_n507), .B2(new_n509), .ZN(G164));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT75), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n511), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n514), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NOR3_X1   g093(.A1(new_n512), .A2(KEYINPUT75), .A3(new_n513), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(G166));
  AND2_X1   g095(.A1(new_n511), .A2(new_n516), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G89), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n511), .A2(KEYINPUT76), .ZN(new_n523));
  OR2_X1    g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT76), .ZN(new_n525));
  NAND2_X1  g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n523), .A2(G63), .A3(G651), .A4(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n522), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT77), .ZN(new_n532));
  AND2_X1   g107(.A1(KEYINPUT6), .A2(G651), .ZN(new_n533));
  NOR2_X1   g108(.A1(KEYINPUT6), .A2(G651), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT6), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(new_n513), .ZN(new_n537));
  NAND2_X1  g112(.A1(KEYINPUT6), .A2(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n537), .A2(KEYINPUT77), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n535), .A2(new_n539), .A3(G543), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT78), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n516), .B2(new_n532), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n544), .A2(KEYINPUT78), .A3(new_n539), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n531), .B1(G51), .B2(new_n546), .ZN(G168));
  NAND2_X1  g122(.A1(G77), .A2(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n523), .A2(new_n527), .ZN(new_n549));
  INV_X1    g124(.A(G64), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g126(.A(KEYINPUT79), .B(G90), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n551), .A2(G651), .B1(new_n521), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n546), .A2(G52), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(G301));
  INV_X1    g130(.A(G301), .ZN(G171));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n549), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n559), .A2(G651), .B1(G81), .B2(new_n521), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n546), .A2(G43), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  NAND4_X1  g143(.A1(new_n535), .A2(new_n539), .A3(G53), .A4(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n544), .A2(new_n571), .A3(G53), .A4(new_n539), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n511), .A2(new_n516), .A3(G91), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n511), .B2(G65), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n574), .B1(new_n577), .B2(new_n513), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n573), .A2(new_n579), .ZN(G299));
  INV_X1    g155(.A(G168), .ZN(G286));
  INV_X1    g156(.A(G166), .ZN(G303));
  NAND2_X1  g157(.A1(new_n521), .A2(G87), .ZN(new_n583));
  INV_X1    g158(.A(G49), .ZN(new_n584));
  AOI21_X1  g159(.A(G74), .B1(new_n523), .B2(new_n527), .ZN(new_n585));
  OAI221_X1 g160(.A(new_n583), .B1(new_n584), .B2(new_n540), .C1(new_n585), .C2(new_n513), .ZN(G288));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n511), .A2(new_n587), .A3(G61), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n587), .B1(new_n511), .B2(G61), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n511), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n595), .A2(new_n517), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT82), .ZN(G305));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n549), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(G85), .B2(new_n521), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n546), .A2(G47), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(new_n546), .A2(G54), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n521), .A2(KEYINPUT10), .A3(G92), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n511), .A2(new_n516), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  INV_X1    g186(.A(new_n511), .ZN(new_n612));
  XNOR2_X1  g187(.A(KEYINPUT83), .B(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n606), .A2(new_n610), .B1(G651), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n605), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G171), .B2(new_n617), .ZN(G284));
  XNOR2_X1  g194(.A(G284), .B(KEYINPUT84), .ZN(G321));
  NAND2_X1  g195(.A1(G299), .A2(new_n617), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G168), .B2(new_n617), .ZN(G297));
  OAI21_X1  g197(.A(new_n621), .B1(G168), .B2(new_n617), .ZN(G280));
  INV_X1    g198(.A(new_n616), .ZN(new_n624));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n562), .A2(new_n617), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n616), .A2(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(new_n617), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g205(.A1(new_n471), .A2(G2105), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n486), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2100), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n495), .A2(G135), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT85), .ZN(new_n637));
  INV_X1    g212(.A(new_n487), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G123), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n480), .A2(G111), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n637), .B(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(G2096), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n635), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n645), .B1(new_n644), .B2(new_n643), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT86), .ZN(G156));
  INV_X1    g222(.A(KEYINPUT14), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(new_n651), .B2(new_n650), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n653), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  AND3_X1   g236(.A1(new_n660), .A2(G14), .A3(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2067), .B(G2678), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT88), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2084), .B(G2090), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT87), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT18), .ZN(new_n670));
  OAI21_X1  g245(.A(KEYINPUT17), .B1(new_n664), .B2(new_n666), .ZN(new_n671));
  AOI22_X1  g246(.A1(new_n671), .A2(new_n668), .B1(new_n664), .B2(new_n666), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n668), .B2(new_n671), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2096), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT20), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n678), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n678), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G229));
  MUX2_X1   g268(.A(G6), .B(G305), .S(G16), .Z(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT32), .B(G1981), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G22), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G166), .B2(new_n698), .ZN(new_n700));
  INV_X1    g275(.A(G1971), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n698), .A2(G23), .ZN(new_n703));
  INV_X1    g278(.A(G288), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(new_n698), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT33), .B(G1976), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  NOR3_X1   g283(.A1(new_n696), .A2(new_n697), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT34), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n698), .A2(G24), .ZN(new_n713));
  INV_X1    g288(.A(G290), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n698), .ZN(new_n715));
  INV_X1    g290(.A(G1986), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G25), .ZN(new_n718));
  OR3_X1    g293(.A1(new_n718), .A2(KEYINPUT89), .A3(G29), .ZN(new_n719));
  OAI21_X1  g294(.A(KEYINPUT89), .B1(new_n718), .B2(G29), .ZN(new_n720));
  OAI221_X1 g295(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n480), .C2(G107), .ZN(new_n721));
  INV_X1    g296(.A(G119), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n487), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G131), .B2(new_n495), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n719), .B(new_n720), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT35), .B(G1991), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n711), .A2(new_n712), .A3(new_n717), .A4(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT36), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n725), .A2(G35), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G162), .B2(new_n725), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT29), .Z(new_n733));
  INV_X1    g308(.A(G2090), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n624), .A2(new_n698), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G4), .B2(new_n698), .ZN(new_n738));
  INV_X1    g313(.A(G1348), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n738), .A2(new_n739), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n735), .A2(new_n736), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n698), .A2(G19), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n563), .B2(new_n698), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(G1341), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n698), .A2(G5), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G171), .B2(new_n698), .ZN(new_n747));
  INV_X1    g322(.A(G1961), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n742), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(G168), .A2(G16), .ZN(new_n752));
  NOR2_X1   g327(.A1(G16), .A2(G21), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(KEYINPUT96), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(KEYINPUT96), .B2(new_n752), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1966), .ZN(new_n756));
  NOR2_X1   g331(.A1(G29), .A2(G33), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n480), .A2(G103), .A3(G2104), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT25), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G139), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n492), .A2(new_n494), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT92), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n486), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n766), .A2(new_n480), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n757), .B1(new_n768), .B2(G29), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(G2072), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT93), .Z(new_n771));
  AND2_X1   g346(.A1(new_n769), .A2(G2072), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n725), .A2(G32), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n495), .A2(G141), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT95), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n638), .A2(G129), .ZN(new_n776));
  NAND3_X1  g351(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT26), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n779), .A2(new_n780), .B1(G105), .B2(new_n631), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n775), .A2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n773), .B1(new_n784), .B2(new_n725), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT27), .B(G1996), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G27), .A2(G29), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G164), .B2(G29), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n643), .A2(G29), .B1(G2078), .B2(new_n789), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n725), .A2(G26), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n495), .A2(G140), .ZN(new_n794));
  NOR2_X1   g369(.A1(G104), .A2(G2105), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT90), .Z(new_n796));
  OAI21_X1  g371(.A(G2104), .B1(new_n480), .B2(G116), .ZN(new_n797));
  INV_X1    g372(.A(G128), .ZN(new_n798));
  OAI22_X1  g373(.A1(new_n796), .A2(new_n797), .B1(new_n798), .B2(new_n487), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n794), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n793), .B1(new_n800), .B2(new_n725), .ZN(new_n801));
  INV_X1    g376(.A(G2067), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n789), .A2(G2078), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT31), .B(G11), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT97), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT30), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n807), .A2(G28), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n725), .B1(new_n807), .B2(G28), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT24), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n725), .B1(new_n810), .B2(G34), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n811), .A2(KEYINPUT94), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(G34), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n811), .B2(KEYINPUT94), .ZN(new_n814));
  OAI22_X1  g389(.A1(new_n482), .A2(new_n725), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(G2084), .ZN(new_n816));
  OAI221_X1 g391(.A(new_n806), .B1(new_n808), .B2(new_n809), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n816), .B2(new_n815), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n790), .A2(new_n803), .A3(new_n804), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n698), .A2(G20), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT23), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n578), .B1(new_n570), .B2(new_n572), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n822), .B2(new_n698), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G1956), .ZN(new_n824));
  NOR4_X1   g399(.A1(new_n772), .A2(new_n787), .A3(new_n819), .A4(new_n824), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n751), .A2(new_n756), .A3(new_n771), .A4(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n730), .A2(new_n826), .ZN(G311));
  INV_X1    g402(.A(G311), .ZN(G150));
  NAND2_X1  g403(.A1(G80), .A2(G543), .ZN(new_n829));
  INV_X1    g404(.A(G67), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n549), .B2(new_n830), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n831), .A2(G651), .B1(G93), .B2(new_n521), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n546), .A2(G55), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(G860), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT37), .Z(new_n836));
  NOR2_X1   g411(.A1(new_n616), .A2(new_n625), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT98), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT38), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n562), .A2(new_n834), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n560), .A2(new_n832), .A3(new_n561), .A4(new_n833), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n839), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n844), .A2(KEYINPUT39), .ZN(new_n845));
  INV_X1    g420(.A(G860), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n844), .B2(KEYINPUT39), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n836), .B1(new_n845), .B2(new_n847), .ZN(G145));
  NAND3_X1  g423(.A1(new_n775), .A2(G164), .A3(new_n782), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(G164), .B1(new_n775), .B2(new_n782), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n800), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n851), .ZN(new_n853));
  INV_X1    g428(.A(new_n800), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n853), .A2(new_n854), .A3(new_n849), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n765), .A2(KEYINPUT100), .A3(new_n767), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT99), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n765), .A2(new_n859), .A3(KEYINPUT100), .A4(new_n767), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n852), .A2(new_n855), .A3(new_n858), .A4(new_n860), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT101), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n862), .A2(new_n866), .A3(new_n863), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n638), .A2(G130), .ZN(new_n868));
  OAI221_X1 g443(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n480), .C2(G118), .ZN(new_n869));
  INV_X1    g444(.A(G142), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n868), .B(new_n869), .C1(new_n762), .C2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n633), .ZN(new_n872));
  INV_X1    g447(.A(new_n724), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n865), .A2(new_n867), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n865), .A2(KEYINPUT102), .A3(new_n867), .A4(new_n874), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n874), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n862), .A2(new_n863), .A3(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(G162), .B(new_n482), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n642), .B(new_n882), .Z(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n879), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n864), .A2(new_n874), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n881), .ZN(new_n889));
  AOI21_X1  g464(.A(G37), .B1(new_n889), .B2(new_n883), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT40), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n885), .B1(new_n877), .B2(new_n878), .ZN(new_n892));
  INV_X1    g467(.A(new_n890), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT40), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n891), .A2(new_n895), .ZN(G395));
  XNOR2_X1  g471(.A(G305), .B(G288), .ZN(new_n897));
  XNOR2_X1  g472(.A(G303), .B(G290), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n897), .B(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT42), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n842), .B(KEYINPUT103), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n628), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n616), .A2(G299), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n605), .A2(new_n822), .A3(new_n615), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT104), .B1(new_n905), .B2(KEYINPUT41), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n907), .B1(new_n903), .B2(new_n904), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n903), .A2(new_n907), .A3(new_n904), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n906), .B1(new_n911), .B2(KEYINPUT104), .ZN(new_n912));
  OR3_X1    g487(.A1(new_n902), .A2(KEYINPUT105), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n905), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n902), .A2(new_n914), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT105), .B1(new_n902), .B2(new_n912), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n900), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND4_X1   g493(.A1(new_n917), .A2(new_n913), .A3(new_n915), .A4(new_n900), .ZN(new_n919));
  OAI21_X1  g494(.A(G868), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n834), .A2(new_n617), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(G295));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n921), .ZN(G331));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n840), .A2(G301), .A3(new_n841), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(G301), .B1(new_n840), .B2(new_n841), .ZN(new_n928));
  OAI21_X1  g503(.A(G286), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n928), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n930), .A2(G168), .A3(new_n926), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n914), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(new_n931), .A3(new_n911), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n899), .ZN(new_n936));
  AOI21_X1  g511(.A(G37), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT106), .B1(new_n932), .B2(new_n912), .ZN(new_n938));
  INV_X1    g513(.A(new_n910), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT104), .B1(new_n939), .B2(new_n908), .ZN(new_n940));
  INV_X1    g515(.A(new_n906), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n942), .A2(new_n943), .A3(new_n931), .A4(new_n929), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n938), .A2(new_n899), .A3(new_n933), .A4(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n925), .B1(new_n937), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n933), .A2(new_n944), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n929), .A2(new_n931), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n943), .B1(new_n948), .B2(new_n942), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n936), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G37), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n950), .A2(new_n925), .A3(new_n951), .A4(new_n945), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n946), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n933), .A2(new_n944), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n899), .B1(new_n955), .B2(new_n938), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n945), .A2(new_n951), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n958), .A2(KEYINPUT108), .A3(new_n925), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n924), .B1(new_n954), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n937), .A2(new_n925), .A3(new_n945), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT107), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT43), .B1(new_n956), .B2(new_n957), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n937), .A2(new_n964), .A3(new_n925), .A4(new_n945), .ZN(new_n965));
  AND4_X1   g540(.A1(new_n924), .A2(new_n962), .A3(new_n963), .A4(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n960), .A2(new_n966), .ZN(G397));
  INV_X1    g542(.A(KEYINPUT120), .ZN(new_n968));
  XNOR2_X1  g543(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(G164), .B2(G1384), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n507), .A2(new_n509), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n503), .A2(new_n504), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1384), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(KEYINPUT45), .A3(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n476), .A2(new_n481), .A3(G40), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT110), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n476), .A2(new_n481), .A3(new_n978), .A4(G40), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n970), .A2(new_n975), .A3(new_n977), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n701), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(G164), .B2(G1384), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n973), .A2(KEYINPUT50), .A3(new_n974), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n977), .A2(new_n734), .A3(new_n979), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(new_n986), .A3(KEYINPUT111), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n981), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT111), .B1(new_n985), .B2(new_n986), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT112), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(G8), .B1(new_n518), .B2(new_n519), .ZN(new_n991));
  XNOR2_X1  g566(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n995));
  OAI211_X1 g570(.A(G8), .B(new_n992), .C1(new_n518), .C2(new_n519), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n995), .B1(new_n994), .B2(new_n996), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT50), .B1(new_n973), .B2(new_n974), .ZN(new_n1001));
  AOI211_X1 g576(.A(new_n982), .B(G1384), .C1(new_n971), .C2(new_n972), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n977), .A2(new_n734), .A3(new_n979), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1000), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1005), .A2(new_n1006), .A3(new_n981), .A4(new_n987), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n990), .A2(G8), .A3(new_n999), .A4(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT49), .ZN(new_n1010));
  INV_X1    g585(.A(G1981), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n594), .A2(new_n1011), .A3(new_n596), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1011), .B1(new_n594), .B2(new_n596), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1010), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1014), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1016), .A2(KEYINPUT49), .A3(new_n1012), .ZN(new_n1017));
  AOI21_X1  g592(.A(G1384), .B1(new_n971), .B2(new_n972), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n977), .A2(new_n1018), .A3(new_n979), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1015), .A2(new_n1017), .A3(G8), .A4(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1976), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1019), .B(G8), .C1(new_n1021), .C2(G288), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT52), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n1026));
  NAND2_X1  g601(.A1(G288), .A2(new_n1021), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI211_X1 g604(.A(KEYINPUT115), .B(KEYINPUT52), .C1(G288), .C2(new_n1021), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1025), .B1(new_n1031), .B2(new_n1022), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1022), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1033), .B(KEYINPUT116), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1024), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1009), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1019), .A2(G8), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1020), .A2(new_n1021), .A3(new_n704), .ZN(new_n1038));
  XOR2_X1   g613(.A(new_n1012), .B(KEYINPUT117), .Z(new_n1039));
  AOI21_X1  g614(.A(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1008), .A2(new_n1035), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n994), .A2(new_n996), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n980), .A2(new_n701), .B1(new_n985), .B2(new_n986), .ZN(new_n1044));
  OAI21_X1  g619(.A(G8), .B1(new_n1044), .B2(KEYINPUT118), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n985), .A2(new_n986), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n981), .A2(KEYINPUT118), .A3(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1043), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT119), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1050), .B(new_n1043), .C1(new_n1045), .C2(new_n1047), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1042), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G1966), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n977), .B(new_n979), .C1(new_n1018), .C2(KEYINPUT45), .ZN(new_n1054));
  NOR3_X1   g629(.A1(G164), .A2(G1384), .A3(new_n969), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1053), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n977), .A2(new_n979), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n985), .A2(new_n816), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G8), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(G286), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT63), .B1(new_n1052), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1007), .A2(G8), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1004), .B1(new_n983), .B2(new_n984), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1064), .A2(KEYINPUT111), .B1(new_n701), .B2(new_n980), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1006), .B1(new_n1065), .B2(new_n1005), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1043), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT63), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1060), .A2(new_n1068), .A3(G286), .ZN(new_n1069));
  AND4_X1   g644(.A1(new_n1008), .A2(new_n1067), .A3(new_n1035), .A4(new_n1069), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n968), .B(new_n1041), .C1(new_n1062), .C2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1008), .A2(new_n1035), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(new_n1073), .A3(new_n1061), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1070), .B1(new_n1074), .B2(new_n1068), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT120), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT126), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n546), .A2(G51), .ZN(new_n1079));
  OAI211_X1 g654(.A(KEYINPUT125), .B(G8), .C1(new_n1079), .C2(new_n531), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT125), .ZN(new_n1081));
  INV_X1    g656(.A(G8), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1081), .B1(G168), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1084), .B1(new_n1059), .B2(G8), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT51), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1078), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1082), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1088));
  OAI211_X1 g663(.A(KEYINPUT126), .B(KEYINPUT51), .C1(new_n1088), .C2(new_n1084), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1060), .B(new_n1086), .C1(new_n1082), .C2(G168), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1087), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1059), .A2(G8), .A3(G286), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n970), .A2(new_n975), .ZN(new_n1094));
  INV_X1    g669(.A(G2078), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1094), .A2(new_n1095), .A3(new_n1057), .ZN(new_n1096));
  XOR2_X1   g671(.A(KEYINPUT127), .B(KEYINPUT53), .Z(new_n1097));
  NAND2_X1  g672(.A1(new_n977), .A2(new_n979), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1098), .B1(new_n983), .B2(new_n984), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1096), .A2(new_n1097), .B1(new_n1100), .B2(new_n748), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1095), .A2(KEYINPUT53), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(G301), .B(KEYINPUT54), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n976), .A2(new_n1103), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1105), .B1(new_n1094), .B2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1104), .A2(new_n1105), .B1(new_n1107), .B2(new_n1101), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1093), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n1110));
  AOI21_X1  g685(.A(G1348), .B1(new_n985), .B2(new_n1057), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1019), .A2(G2067), .ZN(new_n1112));
  NOR4_X1   g687(.A1(new_n1111), .A2(new_n1112), .A3(KEYINPUT60), .A4(new_n616), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n624), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1057), .A2(new_n802), .A3(new_n1018), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1115), .B(new_n616), .C1(new_n1099), .C2(G1348), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1113), .B1(new_n1117), .B2(KEYINPUT60), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n1119));
  NAND3_X1  g694(.A1(G299), .A2(new_n1119), .A3(KEYINPUT57), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n822), .B2(KEYINPUT122), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT56), .B(G2072), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n980), .A2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT121), .B(G1956), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1127), .B1(new_n985), .B2(new_n1057), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1123), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1127), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1003), .B2(new_n1098), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT57), .B1(G299), .B2(new_n1119), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n822), .A2(KEYINPUT122), .A3(new_n1121), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1057), .A2(new_n970), .A3(new_n975), .A4(new_n1124), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1131), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1129), .A2(new_n1136), .A3(KEYINPUT61), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT58), .B(G1341), .Z(new_n1138));
  NAND2_X1  g713(.A1(new_n1019), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(new_n980), .B2(G1996), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n563), .ZN(new_n1141));
  XOR2_X1   g716(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1140), .A2(new_n563), .A3(new_n1142), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1126), .A2(new_n1128), .A3(new_n1123), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1134), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1118), .A2(new_n1137), .A3(new_n1146), .A4(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1148), .A2(new_n1114), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1152), .A2(new_n1149), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1110), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1109), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1151), .A2(new_n1110), .A3(new_n1153), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1093), .A2(KEYINPUT62), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1104), .A2(G171), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1158), .B1(new_n1093), .B2(KEYINPUT62), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1155), .A2(new_n1156), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1052), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1071), .B(new_n1077), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1098), .A2(new_n970), .ZN(new_n1163));
  INV_X1    g738(.A(G1996), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n783), .B(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n800), .B(G2067), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n724), .A2(new_n727), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n724), .A2(new_n727), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(G290), .B(G1986), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1163), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1162), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1163), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1175), .B1(new_n1166), .B2(new_n784), .ZN(new_n1176));
  OAI21_X1  g751(.A(KEYINPUT46), .B1(new_n1175), .B2(G1996), .ZN(new_n1177));
  OR3_X1    g752(.A1(new_n1175), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT47), .ZN(new_n1180));
  AOI22_X1  g755(.A1(new_n1167), .A2(new_n1168), .B1(new_n802), .B2(new_n800), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1181), .A2(new_n1175), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1171), .A2(new_n1163), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n714), .A2(new_n1163), .A3(new_n716), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT48), .ZN(new_n1185));
  AOI211_X1 g760(.A(new_n1180), .B(new_n1182), .C1(new_n1183), .C2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1174), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g762(.A1(new_n887), .A2(new_n890), .ZN(new_n1189));
  NAND3_X1  g763(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n1190));
  NOR4_X1   g764(.A1(G229), .A2(new_n462), .A3(G401), .A4(G227), .ZN(new_n1191));
  AND3_X1   g765(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(G308));
  NAND3_X1  g766(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(G225));
endmodule


