//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 0 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1284, new_n1285,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(new_n202), .A2(new_n203), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G50), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR3_X1   g0013(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  INV_X1    g0015(.A(G1), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n212), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  AOI211_X1 g0022(.A(new_n215), .B(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n214), .B1(new_n223), .B2(KEYINPUT0), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n224), .B1(KEYINPUT0), .B2(new_n223), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT64), .Z(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  INV_X1    g0027(.A(G238), .ZN(new_n228));
  INV_X1    g0028(.A(G87), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n227), .B1(new_n203), .B2(new_n228), .C1(new_n229), .C2(new_n215), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n231));
  INV_X1    g0031(.A(G77), .ZN(new_n232));
  INV_X1    g0032(.A(G244), .ZN(new_n233));
  OAI221_X1 g0033(.A(new_n231), .B1(new_n232), .B2(new_n233), .C1(new_n207), .C2(new_n222), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n218), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT1), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n226), .A2(new_n236), .ZN(G361));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G238), .B(G244), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G232), .ZN(new_n243));
  XOR2_X1   g0043(.A(KEYINPUT2), .B(G226), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT66), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n250), .B(KEYINPUT67), .Z(new_n251));
  NAND2_X1  g0051(.A1(new_n201), .A2(G68), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n203), .A2(G50), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G58), .B(G77), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n251), .B(new_n256), .ZN(G351));
  INV_X1    g0057(.A(KEYINPUT14), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(KEYINPUT73), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(G226), .A3(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(G232), .A3(G1698), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G97), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT72), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n266), .A2(new_n267), .A3(KEYINPUT72), .A4(new_n268), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT13), .ZN(new_n275));
  INV_X1    g0075(.A(G274), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n216), .B1(G41), .B2(G45), .ZN(new_n277));
  NOR3_X1   g0077(.A1(new_n273), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n277), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n278), .B1(G238), .B2(new_n280), .ZN(new_n281));
  AND3_X1   g0081(.A1(new_n274), .A2(new_n275), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n275), .B1(new_n274), .B2(new_n281), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G169), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n259), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(G179), .ZN(new_n287));
  OAI221_X1 g0087(.A(G169), .B1(KEYINPUT73), .B2(new_n258), .C1(new_n282), .C2(new_n283), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n212), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT68), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n290), .B(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G77), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n293), .B1(new_n212), .B2(G68), .C1(new_n201), .C2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n213), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n296), .A2(KEYINPUT11), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G13), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n300), .A2(new_n212), .A3(G1), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  OR3_X1    g0102(.A1(new_n302), .A2(KEYINPUT12), .A3(G68), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT12), .B1(new_n302), .B2(G68), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n301), .A2(new_n298), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n203), .B1(new_n216), .B2(G20), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n303), .A2(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n299), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT11), .B1(new_n296), .B2(new_n298), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT74), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n309), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT74), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n311), .A2(new_n312), .A3(new_n299), .A4(new_n307), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n289), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n283), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n274), .A2(new_n275), .A3(new_n281), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(G190), .A3(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(G200), .B1(new_n282), .B2(new_n283), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n308), .A2(new_n309), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n315), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n305), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT8), .B(G58), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n216), .A2(G20), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n323), .A2(new_n327), .B1(new_n302), .B2(new_n325), .ZN(new_n328));
  AND2_X1   g0128(.A1(KEYINPUT75), .A2(G33), .ZN(new_n329));
  NOR2_X1   g0129(.A1(KEYINPUT75), .A2(G33), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT3), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(new_n212), .A3(new_n262), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT7), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT7), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n331), .A2(new_n334), .A3(new_n212), .A4(new_n262), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(G68), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G58), .A2(G68), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT76), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT76), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n339), .A2(G58), .A3(G68), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n340), .A3(new_n210), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G20), .ZN(new_n342));
  INV_X1    g0142(.A(G159), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n343), .A2(G20), .A3(G33), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT77), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT77), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n342), .A2(new_n348), .A3(new_n345), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n336), .A2(new_n347), .A3(KEYINPUT16), .A4(new_n349), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n350), .A2(new_n298), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT78), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT75), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n261), .ZN(new_n354));
  NAND2_X1  g0154(.A1(KEYINPUT75), .A2(G33), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n260), .A3(new_n355), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n263), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n357));
  AOI21_X1  g0157(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n262), .A2(new_n358), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n356), .A2(new_n357), .B1(new_n359), .B2(new_n334), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n352), .B1(new_n360), .B2(new_n203), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n263), .A2(new_n212), .ZN(new_n362));
  NOR2_X1   g0162(.A1(KEYINPUT3), .A2(G33), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n334), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NOR3_X1   g0164(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT3), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n358), .A2(KEYINPUT7), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n367), .A2(KEYINPUT78), .A3(G68), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n347), .A2(new_n361), .A3(new_n349), .A4(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT16), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n328), .B1(new_n351), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G226), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G1698), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(G223), .B2(G1698), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(new_n262), .B2(new_n331), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n261), .A2(new_n229), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n273), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n278), .B1(G232), .B2(new_n280), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n285), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n378), .A2(new_n379), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n380), .B1(G179), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT18), .B1(new_n372), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n328), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n360), .A2(new_n352), .A3(new_n203), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT78), .B1(new_n367), .B2(G68), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n348), .B1(new_n342), .B2(new_n345), .ZN(new_n388));
  AOI211_X1 g0188(.A(KEYINPUT77), .B(new_n344), .C1(new_n341), .C2(G20), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT16), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n350), .A2(new_n298), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n384), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT18), .ZN(new_n394));
  INV_X1    g0194(.A(new_n382), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G190), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n378), .A2(new_n379), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n381), .B2(G200), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n384), .B(new_n399), .C1(new_n391), .C2(new_n392), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT17), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n371), .A2(new_n298), .A3(new_n350), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n403), .A2(KEYINPUT17), .A3(new_n384), .A4(new_n399), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n383), .A2(new_n396), .A3(new_n402), .A4(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n264), .A2(G222), .A3(new_n265), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n264), .A2(G1698), .ZN(new_n407));
  INV_X1    g0207(.A(G223), .ZN(new_n408));
  OAI221_X1 g0208(.A(new_n406), .B1(new_n232), .B2(new_n264), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n273), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n278), .B1(G226), .B2(new_n280), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  XOR2_X1   g0212(.A(KEYINPUT71), .B(G200), .Z(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n298), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n292), .A2(new_n325), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n294), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n305), .A2(G50), .A3(new_n326), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(G50), .B2(new_n302), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT9), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n410), .A2(G190), .A3(new_n411), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT9), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n418), .B2(new_n420), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n414), .A2(new_n422), .A3(new_n423), .A4(new_n425), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n426), .A2(KEYINPUT10), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(KEYINPUT10), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n324), .A2(new_n295), .B1(new_n212), .B2(new_n232), .ZN(new_n430));
  XNOR2_X1  g0230(.A(KEYINPUT15), .B(G87), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n431), .A2(new_n290), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n298), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT70), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n232), .B1(new_n216), .B2(G20), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n305), .A2(new_n435), .B1(new_n232), .B2(new_n301), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n264), .A2(G232), .A3(new_n265), .ZN(new_n439));
  OAI221_X1 g0239(.A(new_n439), .B1(new_n207), .B2(new_n264), .C1(new_n407), .C2(new_n228), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n273), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n278), .B1(G244), .B2(new_n280), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n413), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n438), .B(new_n444), .C1(new_n397), .C2(new_n443), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n434), .A2(new_n436), .B1(new_n443), .B2(new_n285), .ZN(new_n446));
  INV_X1    g0246(.A(G179), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n441), .A2(new_n447), .A3(new_n442), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n421), .B1(new_n412), .B2(new_n285), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n451), .A2(KEYINPUT69), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n410), .A2(new_n447), .A3(new_n411), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(KEYINPUT69), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n429), .A2(new_n450), .A3(new_n455), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n322), .A2(new_n405), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT23), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(new_n212), .B2(G107), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g0261(.A(KEYINPUT75), .B(G33), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G116), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(new_n463), .B2(G20), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n260), .B1(new_n354), .B2(new_n355), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n212), .B(G87), .C1(new_n465), .C2(new_n363), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT82), .ZN(new_n467));
  AOI21_X1  g0267(.A(G20), .B1(new_n331), .B2(new_n262), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT82), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(new_n469), .A3(G87), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n467), .A2(new_n470), .A3(KEYINPUT22), .ZN(new_n471));
  INV_X1    g0271(.A(new_n264), .ZN(new_n472));
  OR4_X1    g0272(.A1(KEYINPUT22), .A2(new_n472), .A3(G20), .A4(new_n229), .ZN(new_n473));
  AOI211_X1 g0273(.A(KEYINPUT24), .B(new_n464), .C1(new_n471), .C2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT24), .ZN(new_n475));
  OAI21_X1  g0275(.A(KEYINPUT22), .B1(new_n466), .B2(KEYINPUT82), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n469), .B1(new_n468), .B2(G87), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n464), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n298), .B1(new_n474), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n301), .A2(new_n207), .ZN(new_n482));
  OR2_X1    g0282(.A1(new_n482), .A2(KEYINPUT25), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(KEYINPUT25), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n216), .A2(G33), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n305), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n483), .B(new_n484), .C1(new_n486), .C2(new_n207), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n481), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n221), .A2(G1698), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(G250), .B2(G1698), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n491), .B1(new_n262), .B2(new_n331), .ZN(new_n492));
  INV_X1    g0292(.A(G294), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(new_n354), .B2(new_n355), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n273), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n216), .A2(G45), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  OR2_X1    g0297(.A1(KEYINPUT5), .A2(G41), .ZN(new_n498));
  NAND2_X1  g0298(.A1(KEYINPUT5), .A2(G41), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n273), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n273), .A2(new_n276), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n496), .B1(new_n498), .B2(new_n499), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n501), .A2(G264), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n495), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(new_n447), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n495), .A2(new_n504), .A3(KEYINPUT83), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT83), .B1(new_n495), .B2(new_n504), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n506), .B1(new_n509), .B2(G169), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n397), .B1(new_n507), .B2(new_n508), .ZN(new_n512));
  INV_X1    g0312(.A(G200), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n505), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n487), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n489), .A2(new_n511), .B1(new_n481), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n360), .A2(new_n207), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n294), .A2(G77), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G97), .A2(G107), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT6), .B1(new_n208), .B2(new_n519), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n207), .A2(KEYINPUT6), .A3(G97), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n518), .B1(new_n522), .B2(new_n212), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n298), .B1(new_n517), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n301), .A2(KEYINPUT79), .A3(new_n206), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT79), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n302), .B2(G97), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n525), .B(new_n527), .C1(new_n486), .C2(new_n206), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n501), .A2(G257), .B1(new_n502), .B2(new_n503), .ZN(new_n531));
  AND2_X1   g0331(.A1(KEYINPUT4), .A2(G244), .ZN(new_n532));
  AND2_X1   g0332(.A1(KEYINPUT3), .A2(G33), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n265), .B(new_n532), .C1(new_n533), .C2(new_n363), .ZN(new_n534));
  OAI211_X1 g0334(.A(G250), .B(G1698), .C1(new_n533), .C2(new_n363), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G283), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(G244), .B(new_n265), .C1(new_n465), .C2(new_n363), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT4), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n273), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n447), .B(new_n531), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n530), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n531), .B1(new_n540), .B2(new_n541), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT81), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(KEYINPUT81), .B(new_n531), .C1(new_n540), .C2(new_n541), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n543), .B1(new_n548), .B2(new_n285), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n546), .A2(G190), .A3(new_n547), .ZN(new_n550));
  INV_X1    g0350(.A(new_n530), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT80), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n544), .A2(new_n553), .A3(G200), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n553), .B1(new_n544), .B2(G200), .ZN(new_n555));
  OR2_X1    g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n549), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n222), .A2(G1698), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(G257), .B2(G1698), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(new_n262), .B2(new_n331), .ZN(new_n560));
  INV_X1    g0360(.A(G303), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n264), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n273), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n501), .A2(G270), .B1(new_n502), .B2(new_n503), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n563), .A2(new_n564), .A3(G179), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n305), .A2(G116), .A3(new_n485), .ZN(new_n566));
  INV_X1    g0366(.A(G116), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n301), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n297), .A2(new_n213), .B1(G20), .B2(new_n567), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n536), .B(new_n212), .C1(G33), .C2(new_n206), .ZN(new_n570));
  AOI21_X1  g0370(.A(KEYINPUT20), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n569), .A2(KEYINPUT20), .A3(new_n570), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n566), .B(new_n568), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n565), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n563), .A2(new_n564), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n575), .A2(KEYINPUT21), .A3(G169), .A4(new_n573), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n575), .A2(G169), .A3(new_n573), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT21), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n573), .B1(new_n575), .B2(G200), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n397), .B2(new_n575), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n578), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n331), .A2(new_n262), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n228), .A2(G1698), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n585), .A2(new_n586), .B1(G116), .B2(new_n462), .ZN(new_n587));
  OAI211_X1 g0387(.A(G244), .B(G1698), .C1(new_n465), .C2(new_n363), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n541), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n502), .A2(new_n497), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n541), .A2(G250), .A3(new_n496), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n285), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n431), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n594), .A2(new_n302), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n305), .A2(new_n594), .A3(new_n485), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n585), .A2(new_n212), .A3(G68), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT19), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n212), .B1(new_n268), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n229), .A2(new_n206), .A3(new_n207), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n212), .A2(G33), .A3(G97), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n600), .A2(new_n601), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n596), .B(new_n597), .C1(new_n604), .C2(new_n415), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n363), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n606));
  INV_X1    g0406(.A(new_n586), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n463), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI211_X1 g0408(.A(new_n233), .B(new_n265), .C1(new_n331), .C2(new_n262), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n273), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n592), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n447), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n593), .A2(new_n605), .A3(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n413), .B1(new_n589), .B2(new_n592), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n415), .B1(new_n598), .B2(new_n603), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n486), .A2(new_n229), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n615), .A2(new_n595), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n610), .A2(G190), .A3(new_n611), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n614), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n584), .A2(new_n620), .ZN(new_n621));
  AND4_X1   g0421(.A1(new_n457), .A2(new_n516), .A3(new_n557), .A4(new_n621), .ZN(G372));
  INV_X1    g0422(.A(new_n455), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n321), .A2(new_n448), .A3(new_n446), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n315), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n402), .A2(new_n404), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI211_X1 g0427(.A(KEYINPUT18), .B(new_n382), .C1(new_n403), .C2(new_n384), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n394), .B1(new_n393), .B2(new_n395), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT85), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n429), .B(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n623), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n578), .A2(KEYINPUT84), .A3(new_n581), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT84), .ZN(new_n636));
  INV_X1    g0436(.A(new_n581), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n636), .B1(new_n637), .B2(new_n577), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n489), .A2(new_n511), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n481), .A2(new_n515), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n233), .B1(new_n331), .B2(new_n262), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT4), .B1(new_n641), .B2(new_n265), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n273), .B1(new_n642), .B2(new_n537), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT81), .B1(new_n643), .B2(new_n531), .ZN(new_n644));
  INV_X1    g0444(.A(new_n547), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n285), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n543), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n550), .B(new_n551), .C1(new_n555), .C2(new_n554), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n613), .A2(new_n619), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n640), .A2(new_n648), .A3(new_n649), .A4(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n639), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n648), .A2(new_n653), .A3(new_n620), .ZN(new_n654));
  AOI21_X1  g0454(.A(KEYINPUT26), .B1(new_n650), .B2(new_n549), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n613), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n457), .B1(new_n652), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n634), .A2(new_n657), .ZN(G369));
  INV_X1    g0458(.A(G330), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n635), .A2(new_n638), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n216), .A2(new_n212), .A3(G13), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT86), .ZN(new_n663));
  INV_X1    g0463(.A(G213), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(new_n661), .B2(KEYINPUT27), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n573), .ZN(new_n669));
  XOR2_X1   g0469(.A(new_n669), .B(KEYINPUT87), .Z(new_n670));
  OR2_X1    g0470(.A1(new_n660), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n670), .A2(new_n581), .A3(new_n578), .A4(new_n583), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n659), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n489), .A2(new_n668), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n516), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n510), .B1(new_n481), .B2(new_n488), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n668), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n674), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n668), .B1(new_n578), .B2(new_n581), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n516), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n677), .A2(new_n679), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n683), .A2(new_n687), .ZN(G399));
  NOR2_X1   g0488(.A1(new_n220), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n601), .A2(G116), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G1), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n211), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT31), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n610), .A2(new_n611), .ZN(new_n696));
  AOI21_X1  g0496(.A(G179), .B1(new_n495), .B2(new_n504), .ZN(new_n697));
  AND4_X1   g0497(.A1(new_n544), .A2(new_n696), .A3(new_n575), .A4(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n501), .A2(G264), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n495), .A2(new_n699), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n700), .A2(new_n589), .A3(new_n592), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n701), .A2(new_n546), .A3(new_n547), .A4(new_n565), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n698), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n585), .A2(new_n586), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(new_n588), .A3(new_n463), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n592), .B1(new_n706), .B2(new_n273), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n495), .A2(new_n699), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n565), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(KEYINPUT30), .A3(new_n546), .A4(new_n547), .ZN(new_n710));
  AOI211_X1 g0510(.A(new_n695), .B(new_n679), .C1(new_n704), .C2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n565), .A2(new_n707), .A3(new_n708), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n703), .B1(new_n548), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n698), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(new_n710), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(KEYINPUT31), .B1(new_n715), .B2(new_n668), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n516), .A2(new_n557), .A3(new_n621), .A4(new_n679), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n659), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n620), .B1(new_n481), .B2(new_n515), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n578), .A2(new_n581), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n557), .B(new_n720), .C1(new_n677), .C2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n613), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n653), .B1(new_n648), .B2(new_n620), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n650), .A2(new_n549), .A3(KEYINPUT26), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT88), .B1(new_n727), .B2(new_n679), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT88), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n729), .B(new_n668), .C1(new_n722), .C2(new_n726), .ZN(new_n730));
  OAI21_X1  g0530(.A(KEYINPUT29), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n679), .B1(new_n652), .B2(new_n656), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT29), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n719), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n694), .B1(new_n735), .B2(G1), .ZN(G364));
  NAND3_X1  g0536(.A1(new_n671), .A2(new_n659), .A3(new_n672), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n300), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n216), .B1(new_n738), .B2(G45), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n674), .B(new_n737), .C1(new_n689), .C2(new_n740), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT89), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n671), .A2(new_n672), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n689), .A2(new_n740), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT90), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n220), .A2(new_n585), .ZN(new_n749));
  INV_X1    g0549(.A(new_n211), .ZN(new_n750));
  INV_X1    g0550(.A(G45), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n749), .B(new_n752), .C1(new_n751), .C2(new_n256), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n220), .A2(new_n472), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n754), .A2(G355), .B1(new_n567), .B2(new_n220), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n756), .A2(KEYINPUT91), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n213), .B1(G20), .B2(new_n285), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n745), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(new_n756), .B2(KEYINPUT91), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n748), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT92), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n397), .A2(G179), .A3(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n212), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT94), .Z(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n206), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n212), .A2(new_n447), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G200), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT93), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n397), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n768), .B1(G50), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n772), .A2(G190), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n774), .B1(new_n203), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n212), .A2(G179), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G190), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n343), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT32), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n769), .A2(G190), .A3(new_n513), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n472), .B1(new_n784), .B2(G58), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n769), .A2(new_n779), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n782), .B(new_n785), .C1(new_n232), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n413), .A2(new_n778), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n397), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n788), .A2(G190), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n229), .A2(new_n790), .B1(new_n792), .B2(new_n207), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n777), .A2(new_n787), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n780), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n784), .A2(G322), .B1(new_n795), .B2(G329), .ZN(new_n796));
  INV_X1    g0596(.A(G311), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n796), .B(new_n472), .C1(new_n797), .C2(new_n786), .ZN(new_n798));
  INV_X1    g0598(.A(new_n765), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n798), .B1(G294), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT33), .B(G317), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G326), .A2(new_n773), .B1(new_n775), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G283), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n800), .B(new_n802), .C1(new_n803), .C2(new_n792), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n789), .B(KEYINPUT95), .Z(new_n805));
  AOI21_X1  g0605(.A(new_n804), .B1(G303), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n758), .B1(new_n794), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n761), .A2(new_n762), .ZN(new_n808));
  AND4_X1   g0608(.A1(new_n746), .A2(new_n763), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n742), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G396));
  OR2_X1    g0611(.A1(new_n758), .A2(new_n743), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n792), .A2(new_n229), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n784), .A2(G294), .B1(new_n795), .B2(G311), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n814), .B(new_n472), .C1(new_n567), .C2(new_n786), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n768), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(G283), .A2(new_n775), .B1(new_n773), .B2(G303), .ZN(new_n817));
  INV_X1    g0617(.A(new_n805), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n816), .B(new_n817), .C1(new_n207), .C2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n786), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n784), .A2(G143), .B1(new_n820), .B2(G159), .ZN(new_n821));
  INV_X1    g0621(.A(G150), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n776), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G137), .B2(new_n773), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT34), .ZN(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n585), .B1(new_n826), .B2(new_n780), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G58), .B2(new_n799), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n828), .B1(new_n203), .B2(new_n792), .C1(new_n818), .C2(new_n201), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n819), .B1(new_n825), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT96), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n758), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n830), .A2(KEYINPUT96), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n748), .B1(G77), .B2(new_n812), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n437), .A2(new_n668), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n445), .A2(new_n835), .B1(new_n448), .B2(new_n446), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n449), .A2(new_n668), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n834), .B1(new_n743), .B2(new_n839), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n635), .A2(new_n638), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n557), .B(new_n720), .C1(new_n841), .C2(new_n677), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n668), .B1(new_n842), .B2(new_n726), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n838), .ZN(new_n844));
  INV_X1    g0644(.A(new_n836), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT97), .ZN(new_n846));
  INV_X1    g0646(.A(new_n837), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(KEYINPUT97), .B1(new_n836), .B2(new_n837), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n844), .B1(new_n843), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n719), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n747), .B1(new_n851), .B2(new_n852), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n840), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(G384));
  NOR2_X1   g0656(.A1(new_n738), .A2(new_n216), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT40), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n839), .B1(new_n717), .B2(new_n718), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n314), .A2(new_n668), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n315), .A2(new_n321), .A3(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n321), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n314), .B(new_n668), .C1(new_n289), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT16), .B1(new_n390), .B2(new_n336), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n384), .B1(new_n392), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n666), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n405), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n867), .A2(new_n395), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(new_n869), .A3(new_n400), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n393), .A2(new_n395), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n393), .A2(new_n868), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n875), .A2(new_n876), .A3(new_n877), .A4(new_n400), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n871), .A2(new_n879), .A3(KEYINPUT38), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT38), .B1(new_n871), .B2(new_n879), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n858), .B1(new_n865), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n871), .A2(new_n879), .A3(KEYINPUT38), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n875), .A2(new_n876), .A3(new_n400), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(KEYINPUT37), .ZN(new_n886));
  INV_X1    g0686(.A(new_n876), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n878), .A2(new_n886), .B1(new_n405), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n884), .B1(new_n888), .B2(KEYINPUT38), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n889), .A2(KEYINPUT40), .A3(new_n864), .A4(new_n859), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n883), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n716), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n715), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n718), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n457), .A2(new_n894), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n891), .A2(new_n895), .ZN(new_n897));
  NOR3_X1   g0697(.A1(new_n896), .A2(new_n897), .A3(new_n659), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT100), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n886), .A2(new_n878), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n405), .A2(new_n887), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT38), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n880), .A2(new_n903), .A3(KEYINPUT39), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT39), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n874), .A2(new_n878), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n869), .B1(new_n630), .B2(new_n626), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n905), .B1(new_n909), .B2(new_n884), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT99), .B1(new_n904), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT39), .B1(new_n880), .B2(new_n881), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT99), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n884), .B(new_n905), .C1(new_n888), .C2(KEYINPUT38), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n289), .A2(new_n314), .A3(new_n679), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n837), .B1(new_n843), .B2(new_n838), .ZN(new_n920));
  INV_X1    g0720(.A(new_n864), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n920), .A2(new_n882), .A3(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n630), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n922), .B1(new_n923), .B2(new_n666), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n919), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n456), .A2(new_n405), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(new_n315), .A3(new_n321), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n733), .B2(new_n732), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n731), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n634), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n925), .B(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n857), .B1(new_n900), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n900), .B2(new_n931), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT35), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n522), .A2(new_n934), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n213), .A2(new_n212), .A3(new_n567), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT98), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n937), .A2(new_n938), .B1(new_n934), .B2(new_n522), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n938), .B2(new_n937), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT36), .Z(new_n941));
  NAND4_X1  g0741(.A1(new_n750), .A2(G77), .A3(new_n340), .A4(new_n338), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n252), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(G1), .A3(new_n300), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n933), .A2(new_n941), .A3(new_n944), .ZN(G367));
  NOR2_X1   g0745(.A1(new_n786), .A2(new_n803), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n585), .B(new_n946), .C1(G317), .C2(new_n795), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n947), .B1(new_n206), .B2(new_n792), .C1(new_n207), .C2(new_n765), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(G294), .B2(new_n775), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT46), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n805), .B2(G116), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n790), .A2(KEYINPUT46), .A3(new_n567), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n773), .A2(G311), .B1(G303), .B2(new_n784), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT108), .ZN(new_n955));
  INV_X1    g0755(.A(G137), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n786), .A2(new_n201), .B1(new_n780), .B2(new_n956), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n472), .B(new_n957), .C1(G150), .C2(new_n784), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n958), .B1(new_n202), .B2(new_n790), .C1(new_n232), .C2(new_n792), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n766), .A2(G68), .ZN(new_n960));
  INV_X1    g0760(.A(new_n773), .ZN(new_n961));
  INV_X1    g0761(.A(G143), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n960), .B1(new_n961), .B2(new_n962), .C1(new_n343), .C2(new_n776), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n953), .A2(new_n955), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT109), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT47), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n758), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n679), .A2(new_n617), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n613), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n650), .B2(new_n968), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT101), .Z(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n745), .ZN(new_n972));
  INV_X1    g0772(.A(new_n748), .ZN(new_n973));
  INV_X1    g0773(.A(new_n749), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n241), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n759), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(new_n220), .B2(new_n594), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n973), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n967), .A2(new_n972), .A3(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n735), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT44), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n557), .B1(new_n551), .B2(new_n679), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n549), .A2(new_n668), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n981), .B1(new_n687), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n982), .A2(new_n983), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n685), .A2(new_n686), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n986), .A2(KEYINPUT44), .A3(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT45), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n986), .B2(new_n987), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n687), .A2(KEYINPUT45), .A3(new_n984), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n985), .A2(new_n988), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(KEYINPUT104), .ZN(new_n993));
  INV_X1    g0793(.A(new_n681), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n994), .A2(KEYINPUT105), .A3(new_n673), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT105), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n674), .B2(new_n681), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n985), .A2(new_n988), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n990), .A2(new_n991), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT104), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT106), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n1001), .B2(new_n682), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n992), .A2(KEYINPUT106), .A3(new_n683), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n993), .A2(new_n1003), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OR3_X1    g0807(.A1(new_n676), .A2(new_n680), .A3(new_n684), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n685), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(new_n673), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n980), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n689), .B(KEYINPUT41), .Z(new_n1012));
  OAI21_X1  g0812(.A(KEYINPUT107), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1003), .A2(new_n993), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1014), .A2(new_n1015), .A3(new_n735), .A4(new_n1010), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n735), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT107), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1012), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n740), .B1(new_n1013), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n984), .A2(new_n516), .A3(new_n684), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1022), .A2(KEYINPUT42), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n648), .B1(new_n982), .B2(new_n678), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n679), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1022), .A2(KEYINPUT42), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1023), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT102), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n971), .B(KEYINPUT43), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT43), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1029), .A2(new_n1033), .A3(new_n971), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n683), .A2(new_n986), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1035), .A2(KEYINPUT103), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1032), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(KEYINPUT103), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1032), .A2(new_n1034), .A3(KEYINPUT103), .A4(new_n1035), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n979), .B1(new_n1021), .B2(new_n1041), .ZN(G387));
  NAND2_X1  g0842(.A1(new_n681), .A2(new_n745), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n691), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n754), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(G107), .B2(new_n219), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n245), .A2(new_n751), .ZN(new_n1047));
  AOI211_X1 g0847(.A(G45), .B(new_n1044), .C1(G68), .C2(G77), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n324), .A2(G50), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT50), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n974), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1046), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n748), .B1(new_n1052), .B2(new_n976), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT110), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G159), .A2(new_n773), .B1(new_n775), .B2(new_n325), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n786), .A2(new_n203), .B1(new_n780), .B2(new_n822), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n606), .B(new_n1056), .C1(G50), .C2(new_n784), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G77), .A2(new_n789), .B1(new_n791), .B2(G97), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n766), .A2(new_n594), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1055), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n585), .B1(G326), .B2(new_n795), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n790), .A2(new_n493), .B1(new_n803), .B2(new_n765), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n784), .A2(G317), .B1(new_n820), .B2(G303), .ZN(new_n1063));
  INV_X1    g0863(.A(G322), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1063), .B1(new_n961), .B2(new_n1064), .C1(new_n797), .C2(new_n776), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT48), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1062), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n1066), .B2(new_n1065), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT49), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1061), .B1(new_n567), .B2(new_n792), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1060), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1054), .B1(new_n1072), .B2(new_n758), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1010), .A2(new_n740), .B1(new_n1043), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1010), .A2(new_n735), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n689), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1010), .A2(new_n735), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1074), .B1(new_n1076), .B2(new_n1077), .ZN(G393));
  AND2_X1   g0878(.A1(new_n250), .A2(new_n749), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n759), .B1(new_n206), .B2(new_n219), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n748), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n773), .A2(G150), .B1(G159), .B2(new_n784), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT111), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1083), .A2(KEYINPUT51), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(KEYINPUT51), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n585), .B1(new_n962), .B2(new_n780), .C1(new_n324), .C2(new_n786), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1086), .B(new_n813), .C1(G68), .C2(new_n789), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(G50), .A2(new_n775), .B1(new_n766), .B2(G77), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n773), .A2(G317), .B1(G311), .B2(new_n784), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT52), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n472), .B1(new_n780), .B2(new_n1064), .C1(new_n493), .C2(new_n786), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G116), .B2(new_n799), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G107), .A2(new_n791), .B1(new_n789), .B2(G283), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1093), .B(new_n1094), .C1(new_n776), .C2(new_n561), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1089), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1081), .B1(new_n1096), .B2(new_n758), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n745), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1097), .B1(new_n984), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1015), .B1(new_n683), .B2(new_n992), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1099), .B1(new_n1100), .B2(new_n739), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1016), .A2(new_n689), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1075), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(G390));
  NAND2_X1  g0905(.A1(new_n719), .A2(new_n457), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n677), .A2(new_n721), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1107), .A2(new_n651), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n679), .B1(new_n1108), .B2(new_n656), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n729), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n727), .A2(KEYINPUT88), .A3(new_n679), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n733), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n734), .A2(new_n457), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n634), .B(new_n1106), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT112), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n847), .B1(new_n732), .B2(new_n839), .ZN(new_n1117));
  AND4_X1   g0917(.A1(G330), .A2(new_n864), .A3(new_n894), .A4(new_n838), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n864), .B1(new_n719), .B2(new_n838), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n728), .A2(new_n730), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n836), .B1(new_n1121), .B2(new_n847), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n894), .A2(new_n850), .A3(G330), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n921), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n719), .A2(new_n838), .A3(new_n864), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1120), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n929), .A2(KEYINPUT112), .A3(new_n634), .A4(new_n1106), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1116), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n911), .A2(new_n915), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1110), .A2(new_n1111), .A3(new_n847), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1132), .A2(new_n845), .A3(new_n864), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n889), .A2(new_n917), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1131), .A2(new_n1135), .A3(new_n1125), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1125), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1129), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n689), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1131), .A2(new_n1135), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1118), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1131), .A2(new_n1135), .A3(new_n1125), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(KEYINPUT113), .B1(new_n1143), .B2(new_n1129), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT113), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1116), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1139), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1145), .A2(new_n740), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n748), .B1(new_n325), .B2(new_n812), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n789), .A2(G150), .ZN(new_n1152));
  XOR2_X1   g0952(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n1153));
  XNOR2_X1  g0953(.A(new_n1152), .B(new_n1153), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(G128), .A2(new_n773), .B1(new_n766), .B2(G159), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n775), .A2(G137), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT54), .B(G143), .ZN(new_n1157));
  INV_X1    g0957(.A(G125), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n786), .A2(new_n1157), .B1(new_n780), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n264), .B1(new_n783), .B2(new_n826), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1159), .B(new_n1160), .C1(new_n791), .C2(G50), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1161), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n472), .B1(new_n780), .B2(new_n493), .C1(new_n783), .C2(new_n567), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n792), .A2(new_n203), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(G77), .C2(new_n766), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n803), .B2(new_n961), .C1(new_n818), .C2(new_n229), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n775), .A2(G107), .B1(G97), .B2(new_n820), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT115), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1162), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1151), .B1(new_n1169), .B2(new_n758), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n916), .B2(new_n744), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1150), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1149), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(G378));
  OAI21_X1  g0974(.A(new_n747), .B1(G50), .B2(new_n812), .ZN(new_n1175));
  INV_X1    g0975(.A(G41), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n261), .A2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT116), .ZN(new_n1178));
  AOI211_X1 g0978(.A(G50), .B(new_n1178), .C1(new_n1176), .C2(new_n606), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT117), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n960), .B1(new_n961), .B2(new_n567), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n784), .A2(G107), .B1(new_n820), .B2(new_n594), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n803), .B2(new_n780), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G77), .B2(new_n789), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n791), .A2(G58), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1184), .A2(new_n1176), .A3(new_n606), .A4(new_n1185), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1181), .B(new_n1186), .C1(G97), .C2(new_n775), .ZN(new_n1187));
  XOR2_X1   g0987(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n1188));
  OAI21_X1  g0988(.A(new_n1180), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G132), .A2(new_n775), .B1(new_n766), .B2(G150), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n773), .A2(G125), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1157), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n789), .A2(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n784), .A2(G128), .B1(new_n820), .B2(G137), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1191), .A2(new_n1192), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT119), .Z(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n791), .A2(G159), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n795), .A2(G124), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1198), .A2(new_n1199), .A3(new_n1178), .A4(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1190), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1175), .B1(new_n1203), .B2(new_n758), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n421), .A2(new_n666), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n429), .A2(new_n632), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT85), .B1(new_n427), .B2(new_n428), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1205), .B1(new_n1208), .B2(new_n623), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1205), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n633), .A2(new_n455), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1209), .A2(new_n1211), .A3(new_n1213), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1204), .B1(new_n1217), .B2(new_n744), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT120), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n883), .A2(G330), .A3(new_n890), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1217), .A2(new_n883), .A3(G330), .A4(new_n890), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n925), .A2(new_n1225), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n919), .A2(new_n1223), .A3(new_n924), .A4(new_n1224), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1226), .A2(KEYINPUT121), .A3(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n919), .A2(new_n924), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT121), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1228), .A2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1220), .B1(new_n1232), .B2(new_n739), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1116), .A2(new_n1128), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1146), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1237));
  AND4_X1   g1037(.A1(new_n1146), .A2(new_n1147), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1236), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1232), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT57), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1235), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT57), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n689), .B1(new_n1242), .B2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1234), .B1(new_n1241), .B2(new_n1246), .ZN(G375));
  NAND2_X1  g1047(.A1(new_n921), .A2(new_n743), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n748), .B1(G68), .B2(new_n812), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n805), .A2(G97), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n472), .B1(new_n786), .B2(new_n207), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n783), .A2(new_n803), .B1(new_n780), .B2(new_n561), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1251), .B(new_n1252), .C1(new_n791), .C2(G77), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(G116), .A2(new_n775), .B1(new_n773), .B2(G294), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1250), .A2(new_n1059), .A3(new_n1253), .A4(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1185), .A2(new_n585), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n805), .A2(G159), .B1(KEYINPUT122), .B2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(KEYINPUT122), .B2(new_n1256), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(G132), .A2(new_n773), .B1(new_n775), .B2(new_n1193), .ZN(new_n1259));
  INV_X1    g1059(.A(G128), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n786), .A2(new_n822), .B1(new_n780), .B2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(G137), .B2(new_n784), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1259), .B(new_n1262), .C1(new_n201), .C2(new_n767), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1255), .B1(new_n1258), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1249), .B1(new_n1264), .B2(new_n758), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1248), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1127), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1266), .B1(new_n1267), .B2(new_n739), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT123), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT123), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1270), .B(new_n1266), .C1(new_n1267), .C2(new_n739), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1127), .B1(new_n1116), .B2(new_n1128), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1129), .A2(new_n1019), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1272), .B1(new_n1273), .B2(new_n1274), .ZN(G381));
  OR3_X1    g1075(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1276));
  NOR4_X1   g1076(.A1(G387), .A2(G390), .A3(new_n1276), .A4(G381), .ZN(new_n1277));
  XOR2_X1   g1077(.A(new_n1277), .B(KEYINPUT124), .Z(new_n1278));
  AOI21_X1  g1078(.A(new_n690), .B1(new_n1239), .B2(new_n1244), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1243), .B1(new_n1242), .B2(new_n1232), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1233), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1173), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1278), .A2(new_n1282), .ZN(G407));
  INV_X1    g1083(.A(new_n1282), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n667), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G213), .B(new_n1285), .C1(new_n1278), .C2(new_n1282), .ZN(G409));
  XNOR2_X1  g1086(.A(G393), .B(new_n810), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NOR3_X1   g1088(.A1(new_n1011), .A2(KEYINPUT107), .A3(new_n1012), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1018), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n739), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(G390), .B1(new_n1293), .B2(new_n979), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n979), .ZN(new_n1295));
  AOI211_X1 g1095(.A(new_n1295), .B(new_n1104), .C1(new_n1291), .C2(new_n1292), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1288), .B1(new_n1294), .B2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1293), .A2(new_n979), .A3(G390), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G387), .A2(new_n1104), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1287), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n664), .A2(G343), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1227), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n740), .B1(new_n1303), .B2(new_n1229), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1220), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1149), .A2(new_n1172), .A3(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1239), .A2(new_n1019), .A3(new_n1240), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1302), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1273), .B1(KEYINPUT60), .B2(new_n1129), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1235), .A2(KEYINPUT60), .A3(new_n1267), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n689), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1272), .B1(new_n1309), .B2(new_n1311), .ZN(new_n1312));
  AND2_X1   g1112(.A1(new_n1312), .A2(new_n855), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1272), .B(G384), .C1(new_n1309), .C2(new_n1311), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1316));
  OAI211_X1 g1116(.A(new_n1308), .B(new_n1316), .C1(new_n1281), .C2(new_n1173), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT62), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(G375), .A2(G378), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1320), .A2(KEYINPUT62), .A3(new_n1316), .A4(new_n1308), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1319), .A2(KEYINPUT127), .A3(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1312), .A2(new_n855), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT125), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1323), .A2(new_n1324), .A3(new_n1314), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1302), .A2(G2897), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(KEYINPUT125), .B1(new_n1313), .B2(new_n1315), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1323), .A2(new_n1324), .A3(new_n1314), .A4(new_n1326), .ZN(new_n1330));
  AND3_X1   g1130(.A1(new_n1328), .A2(new_n1329), .A3(new_n1330), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1308), .B1(new_n1281), .B2(new_n1173), .ZN(new_n1332));
  AOI21_X1  g1132(.A(KEYINPUT61), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT127), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1317), .A2(new_n1334), .A3(new_n1318), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1333), .A2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1301), .B1(new_n1322), .B2(new_n1336), .ZN(new_n1337));
  OAI211_X1 g1137(.A(new_n689), .B(new_n1138), .C1(new_n1237), .C2(new_n1238), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1172), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1338), .A2(new_n1339), .A3(new_n1220), .A4(new_n1304), .ZN(new_n1340));
  NOR3_X1   g1140(.A1(new_n1242), .A2(new_n1012), .A3(new_n1232), .ZN(new_n1341));
  OAI22_X1  g1141(.A1(new_n1340), .A2(new_n1341), .B1(new_n664), .B2(G343), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1342), .B1(G378), .B2(G375), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1343), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(new_n1316), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT126), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT63), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1345), .B1(new_n1317), .B2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1344), .A2(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1301), .B1(new_n1346), .B2(new_n1317), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1348), .A2(new_n1349), .A3(new_n1333), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1337), .A2(new_n1350), .ZN(G405));
  NAND2_X1  g1151(.A1(new_n1320), .A2(new_n1282), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1352), .A2(new_n1316), .ZN(new_n1353));
  OAI211_X1 g1153(.A(new_n1320), .B(new_n1282), .C1(new_n1313), .C2(new_n1315), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1301), .ZN(new_n1356));
  XNOR2_X1  g1156(.A(new_n1355), .B(new_n1356), .ZN(G402));
endmodule


