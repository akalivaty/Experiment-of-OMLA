//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1299,
    new_n1300;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n202), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n215), .B1(new_n201), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n209), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT64), .Z(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT65), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n203), .A2(G50), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR3_X1   g0026(.A1(new_n225), .A2(new_n207), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n209), .A2(G13), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT0), .Z(new_n230));
  NOR4_X1   g0030(.A1(new_n222), .A2(new_n224), .A3(new_n227), .A4(new_n230), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G58), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT8), .ZN(new_n248));
  OR3_X1    g0048(.A1(new_n248), .A2(new_n201), .A3(KEYINPUT69), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n248), .B1(new_n201), .B2(KEYINPUT69), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G13), .ZN(new_n253));
  NOR3_X1   g0053(.A1(new_n253), .A2(new_n207), .A3(G1), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n207), .A2(G1), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n226), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT68), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n253), .A2(G1), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G20), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n258), .A2(KEYINPUT68), .A3(new_n226), .ZN(new_n264));
  AND3_X1   g0064(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT70), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n261), .A2(new_n264), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT70), .B1(new_n268), .B2(new_n254), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n257), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n256), .B1(new_n270), .B2(new_n251), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT74), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G58), .A2(G68), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n207), .B1(new_n203), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G159), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n273), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(G58), .A2(G68), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G58), .A2(G68), .ZN(new_n281));
  OAI21_X1  g0081(.A(G20), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(KEYINPUT74), .A3(new_n277), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT7), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT3), .B(G33), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n285), .B1(new_n286), .B2(G20), .ZN(new_n287));
  INV_X1    g0087(.A(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT3), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT3), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n202), .B1(new_n287), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n272), .B1(new_n284), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT77), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT77), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n297), .B(new_n272), .C1(new_n284), .C2(new_n294), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  AND3_X1   g0099(.A1(new_n282), .A2(KEYINPUT74), .A3(new_n277), .ZN(new_n300));
  AOI21_X1  g0100(.A(KEYINPUT74), .B1(new_n282), .B2(new_n277), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT75), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT75), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n279), .B2(new_n283), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n286), .A2(new_n285), .A3(G20), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n290), .A2(G33), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n288), .A2(KEYINPUT3), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT73), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT73), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n289), .A2(new_n291), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n207), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n305), .B1(new_n311), .B2(new_n285), .ZN(new_n312));
  OAI22_X1  g0112(.A1(new_n302), .A2(new_n304), .B1(new_n312), .B2(new_n202), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT16), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n259), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n271), .B1(new_n299), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G274), .ZN(new_n317));
  AND2_X1   g0117(.A1(G1), .A2(G13), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G41), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n319), .A2(G1), .A3(G13), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n321), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n323), .B1(new_n216), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G1698), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n286), .A2(G223), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n286), .A2(G1698), .ZN(new_n329));
  INV_X1    g0129(.A(G226), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n328), .B1(new_n288), .B2(new_n212), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n324), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n326), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n333), .A2(G179), .ZN(new_n334));
  INV_X1    g0134(.A(G169), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n316), .A2(new_n338), .A3(KEYINPUT18), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT78), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT78), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n316), .A2(new_n338), .A3(new_n341), .A4(KEYINPUT18), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n316), .A2(new_n338), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT18), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n340), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G190), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n333), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(G200), .B2(new_n333), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n271), .B(new_n349), .C1(new_n299), .C2(new_n315), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT17), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT79), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT79), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n346), .A2(new_n354), .A3(new_n351), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n270), .A2(G50), .ZN(new_n356));
  OAI21_X1  g0156(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n357));
  INV_X1    g0157(.A(G150), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n207), .A2(new_n288), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n207), .A2(G33), .ZN(new_n360));
  OAI221_X1 g0160(.A(new_n357), .B1(new_n358), .B2(new_n359), .C1(new_n251), .C2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G50), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n361), .A2(new_n268), .B1(new_n362), .B2(new_n254), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n356), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n286), .A2(G222), .A3(new_n327), .ZN(new_n365));
  INV_X1    g0165(.A(G77), .ZN(new_n366));
  INV_X1    g0166(.A(G223), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n365), .B1(new_n366), .B2(new_n286), .C1(new_n329), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n332), .ZN(new_n369));
  INV_X1    g0169(.A(new_n323), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n325), .A2(KEYINPUT67), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT67), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n324), .A2(new_n372), .A3(new_n321), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n370), .B1(new_n374), .B2(G226), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n369), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n335), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n364), .B(new_n377), .C1(G179), .C2(new_n376), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G20), .A2(G77), .ZN(new_n379));
  XNOR2_X1  g0179(.A(KEYINPUT15), .B(G87), .ZN(new_n380));
  XNOR2_X1  g0180(.A(KEYINPUT8), .B(G58), .ZN(new_n381));
  OAI221_X1 g0181(.A(new_n379), .B1(new_n380), .B2(new_n360), .C1(new_n359), .C2(new_n381), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n382), .A2(new_n259), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n254), .A2(new_n259), .ZN(new_n384));
  INV_X1    g0184(.A(new_n257), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(G77), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(G77), .B2(new_n263), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n374), .A2(G244), .ZN(new_n389));
  NOR2_X1   g0189(.A1(G232), .A2(G1698), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n327), .A2(G238), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n286), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n392), .B(new_n332), .C1(G107), .C2(new_n286), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n389), .A2(new_n323), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n388), .B1(new_n335), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(G179), .B2(new_n394), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(G200), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n397), .B(new_n388), .C1(new_n347), .C2(new_n394), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n364), .A2(KEYINPUT9), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT9), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n356), .A2(new_n401), .A3(new_n363), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT10), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n376), .A2(new_n347), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n405), .B1(G200), .B2(new_n376), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n403), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n404), .B1(new_n403), .B2(new_n406), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n378), .B(new_n399), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT71), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G97), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(G226), .A2(G1698), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n216), .B2(G1698), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n413), .B1(new_n415), .B2(new_n286), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n411), .B1(new_n416), .B2(new_n324), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n330), .A2(new_n327), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n216), .A2(G1698), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n412), .B1(new_n292), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(KEYINPUT71), .A3(new_n332), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n324), .A2(new_n372), .A3(new_n321), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n372), .B1(new_n324), .B2(new_n321), .ZN(new_n424));
  OAI21_X1  g0224(.A(G238), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n417), .A2(new_n323), .A3(new_n422), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT13), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n370), .B1(new_n374), .B2(G238), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT13), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n428), .A2(new_n429), .A3(new_n422), .A4(new_n417), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n427), .A2(KEYINPUT72), .A3(new_n430), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n417), .A2(new_n422), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT72), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(new_n429), .A4(new_n428), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n431), .A2(G169), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT14), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT14), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n431), .A2(new_n434), .A3(new_n437), .A4(G169), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n427), .A2(G179), .A3(new_n430), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n276), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n366), .B2(new_n360), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n268), .A2(new_n442), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n443), .A2(KEYINPUT11), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n254), .A2(new_n202), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT12), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n443), .A2(KEYINPUT11), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n384), .A2(G68), .A3(new_n385), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n444), .A2(new_n446), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n440), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n431), .A2(G200), .A3(new_n434), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n347), .B1(new_n426), .B2(KEYINPUT13), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n449), .B1(new_n452), .B2(new_n430), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n410), .A2(new_n455), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n353), .A2(new_n355), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT87), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n289), .A2(new_n291), .A3(G264), .A4(G1698), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n289), .A2(new_n291), .A3(G257), .A4(new_n327), .ZN(new_n460));
  INV_X1    g0260(.A(G303), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n459), .B(new_n460), .C1(new_n461), .C2(new_n286), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n332), .ZN(new_n463));
  INV_X1    g0263(.A(G45), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(G1), .ZN(new_n465));
  INV_X1    g0265(.A(G41), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT5), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT81), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(G41), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n320), .A2(new_n465), .A3(new_n467), .A4(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(new_n465), .A3(new_n467), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(G270), .A3(new_n324), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n463), .A2(G179), .A3(new_n471), .A4(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n207), .A2(G116), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n262), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n259), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n263), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n206), .A2(G33), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G116), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n476), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G283), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n482), .B(new_n207), .C1(G33), .C2(new_n217), .ZN(new_n483));
  INV_X1    g0283(.A(new_n475), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n483), .A2(new_n484), .A3(new_n259), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT20), .ZN(new_n486));
  OR2_X1    g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n486), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n481), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n458), .B1(new_n474), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n473), .A2(new_n471), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n491), .B1(new_n332), .B2(new_n462), .ZN(new_n492));
  INV_X1    g0292(.A(new_n480), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n384), .A2(new_n493), .B1(new_n262), .B2(new_n475), .ZN(new_n494));
  INV_X1    g0294(.A(new_n488), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n485), .A2(new_n486), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n492), .A2(new_n497), .A3(KEYINPUT87), .A4(G179), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n490), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n463), .A2(new_n471), .A3(new_n473), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n497), .A2(new_n500), .A3(G169), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT21), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n497), .A2(new_n500), .A3(KEYINPUT21), .A4(G169), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n463), .A2(G190), .A3(new_n471), .A4(new_n473), .ZN(new_n505));
  INV_X1    g0305(.A(G200), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n505), .B(new_n489), .C1(new_n492), .C2(new_n506), .ZN(new_n507));
  AND4_X1   g0307(.A1(new_n499), .A2(new_n503), .A3(new_n504), .A4(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n472), .A2(G264), .A3(new_n324), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT88), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n472), .A2(KEYINPUT88), .A3(G264), .A4(new_n324), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n289), .A2(new_n291), .A3(G250), .A4(new_n327), .ZN(new_n514));
  INV_X1    g0314(.A(G294), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n514), .B1(new_n288), .B2(new_n515), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n292), .A2(new_n218), .A3(new_n327), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n332), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n513), .A2(new_n471), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n335), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n289), .A2(new_n291), .A3(new_n207), .A4(G87), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT22), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT22), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n286), .A2(new_n523), .A3(new_n207), .A4(G87), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT23), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n207), .B2(G107), .ZN(new_n527));
  INV_X1    g0327(.A(G107), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n528), .A2(KEYINPUT23), .A3(G20), .ZN(new_n529));
  INV_X1    g0329(.A(G116), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n288), .A2(new_n530), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n527), .A2(new_n529), .B1(new_n531), .B2(new_n207), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n525), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT24), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT24), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n525), .A2(new_n535), .A3(new_n532), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n477), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n263), .A2(G107), .ZN(new_n538));
  XNOR2_X1  g0338(.A(new_n538), .B(KEYINPUT25), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n261), .A2(new_n263), .A3(new_n264), .A4(new_n479), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n539), .B1(new_n528), .B2(new_n540), .ZN(new_n541));
  OAI221_X1 g0341(.A(new_n520), .B1(G179), .B2(new_n519), .C1(new_n537), .C2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n537), .A2(new_n541), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n519), .A2(new_n506), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n513), .A2(new_n347), .A3(new_n471), .A4(new_n518), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT89), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n543), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n547), .B1(new_n543), .B2(new_n546), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n508), .B(new_n542), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n320), .A2(new_n465), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n213), .B1(new_n206), .B2(G45), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n324), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n211), .A2(new_n327), .ZN(new_n555));
  INV_X1    g0355(.A(G244), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G1698), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n289), .A2(new_n555), .A3(new_n291), .A4(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n531), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n324), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(G169), .B1(new_n554), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n320), .A2(new_n465), .B1(new_n324), .B2(new_n552), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n555), .A2(new_n557), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n531), .B1(new_n563), .B2(new_n286), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n562), .B(G179), .C1(new_n564), .C2(new_n324), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT83), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT85), .ZN(new_n569));
  INV_X1    g0369(.A(new_n380), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n265), .A2(new_n569), .A3(new_n570), .A4(new_n479), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT85), .B1(new_n540), .B2(new_n380), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT19), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n574), .A2(new_n207), .A3(G33), .A4(G97), .ZN(new_n575));
  NOR2_X1   g0375(.A1(G97), .A2(G107), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n576), .A2(new_n212), .B1(new_n412), .B2(new_n207), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n575), .B1(new_n577), .B2(new_n574), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n286), .A2(KEYINPUT84), .A3(new_n207), .A4(G68), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n289), .A2(new_n291), .A3(new_n207), .A4(G68), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT84), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n578), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n583), .A2(new_n259), .B1(new_n254), .B2(new_n380), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n573), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n561), .A2(new_n565), .A3(KEYINPUT83), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n568), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n265), .A2(G87), .A3(new_n479), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n562), .B(G190), .C1(new_n564), .C2(new_n324), .ZN(new_n589));
  OAI21_X1  g0389(.A(G200), .B1(new_n554), .B2(new_n560), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n584), .A2(new_n588), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT86), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n472), .A2(G257), .A3(new_n324), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n289), .A2(new_n291), .A3(G244), .A4(new_n327), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT4), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n286), .A2(KEYINPUT4), .A3(G244), .A4(new_n327), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n286), .A2(G250), .A3(G1698), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n482), .A4(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n595), .B1(new_n601), .B2(new_n332), .ZN(new_n602));
  AOI21_X1  g0402(.A(G169), .B1(new_n602), .B2(new_n471), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT82), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n601), .A2(new_n332), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(new_n594), .A3(new_n471), .ZN(new_n606));
  OAI22_X1  g0406(.A1(new_n603), .A2(new_n604), .B1(G179), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(G179), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n602), .A2(KEYINPUT82), .A3(new_n608), .A4(new_n471), .ZN(new_n609));
  MUX2_X1   g0409(.A(new_n263), .B(new_n540), .S(G97), .Z(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT7), .B1(new_n292), .B2(new_n207), .ZN(new_n611));
  OAI21_X1  g0411(.A(G107), .B1(new_n305), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT6), .ZN(new_n613));
  AND2_X1   g0413(.A1(G97), .A2(G107), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n613), .B1(new_n614), .B2(new_n576), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n528), .A2(KEYINPUT6), .A3(G97), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n617), .A2(G20), .B1(G77), .B2(new_n276), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n477), .B1(new_n612), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT80), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI211_X1 g0421(.A(KEYINPUT80), .B(new_n477), .C1(new_n612), .C2(new_n618), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n610), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n607), .A2(new_n609), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT86), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n587), .A2(new_n625), .A3(new_n591), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n615), .A2(new_n616), .ZN(new_n627));
  OAI22_X1  g0427(.A1(new_n627), .A2(new_n207), .B1(new_n366), .B2(new_n359), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n528), .B1(new_n287), .B2(new_n293), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n259), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT80), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n619), .A2(new_n620), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n606), .A2(G200), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n602), .A2(G190), .A3(new_n471), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n633), .A2(new_n610), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n593), .A2(new_n624), .A3(new_n626), .A4(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n550), .A2(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n457), .A2(new_n638), .ZN(G372));
  INV_X1    g0439(.A(new_n626), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n625), .B1(new_n587), .B2(new_n591), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n640), .A2(new_n624), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g0442(.A(KEYINPUT91), .B(KEYINPUT26), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n607), .A2(new_n609), .A3(new_n623), .ZN(new_n645));
  AND4_X1   g0445(.A1(new_n584), .A2(new_n588), .A3(new_n589), .A4(new_n590), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n573), .A2(new_n584), .B1(new_n561), .B2(new_n565), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT90), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n585), .A2(new_n566), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT90), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(new_n650), .A3(new_n591), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n642), .A2(new_n644), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n542), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n499), .A2(new_n503), .A3(new_n504), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n624), .B(new_n636), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n652), .B1(new_n548), .B2(new_n549), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n649), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n457), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n408), .A2(new_n409), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT17), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n350), .B(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n454), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(new_n396), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n665), .B1(new_n667), .B2(new_n450), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n267), .A2(new_n269), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n385), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n255), .B1(new_n670), .B2(new_n252), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n289), .A2(new_n291), .A3(new_n309), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n309), .B1(new_n289), .B2(new_n291), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n672), .A2(new_n673), .A3(G20), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n293), .B1(new_n674), .B2(KEYINPUT7), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT75), .B1(new_n300), .B2(new_n301), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n279), .A2(new_n283), .A3(new_n303), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n675), .A2(G68), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n477), .B1(new_n678), .B2(KEYINPUT16), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n296), .A2(new_n298), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n671), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n681), .A2(new_n344), .A3(new_n337), .ZN(new_n682));
  AOI21_X1  g0482(.A(KEYINPUT18), .B1(new_n316), .B2(new_n338), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n663), .B1(new_n668), .B2(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n685), .A2(new_n378), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n662), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT92), .ZN(G369));
  NAND2_X1  g0488(.A1(new_n262), .A2(new_n207), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G213), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(G343), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(new_n489), .ZN(new_n696));
  MUX2_X1   g0496(.A(new_n508), .B(new_n657), .S(new_n696), .Z(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  OAI22_X1  g0498(.A1(new_n548), .A2(new_n549), .B1(new_n543), .B2(new_n695), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n542), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n656), .A2(new_n695), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n702), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n657), .A2(new_n695), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n704), .A2(new_n701), .A3(new_n708), .ZN(G399));
  INV_X1    g0509(.A(new_n228), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G41), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n576), .A2(new_n212), .A3(new_n530), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n711), .A2(new_n712), .A3(new_n206), .ZN(new_n713));
  INV_X1    g0513(.A(new_n225), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(new_n711), .ZN(new_n715));
  XOR2_X1   g0515(.A(new_n715), .B(KEYINPUT28), .Z(new_n716));
  INV_X1    g0516(.A(KEYINPUT29), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n717), .B(new_n695), .C1(new_n655), .C2(new_n660), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n550), .A2(new_n637), .A3(new_n694), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n554), .A2(new_n560), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n513), .A2(new_n720), .A3(new_n518), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT94), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n474), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n513), .A2(new_n720), .A3(KEYINPUT94), .A4(new_n518), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n723), .A2(new_n602), .A3(new_n724), .A4(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n724), .A2(new_n602), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n729), .A2(new_n723), .A3(KEYINPUT30), .A4(new_n725), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n720), .A2(G179), .ZN(new_n731));
  AND4_X1   g0531(.A1(new_n606), .A2(new_n519), .A3(new_n500), .A4(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n728), .A2(new_n730), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g0534(.A(KEYINPUT93), .B(KEYINPUT31), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n734), .A2(new_n694), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n732), .B1(new_n726), .B2(new_n727), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n695), .B1(new_n738), .B2(new_n730), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n737), .B1(KEYINPUT31), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(G330), .B1(new_n719), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n660), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n642), .A2(new_n644), .B1(new_n653), .B2(new_n654), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n694), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n718), .B(new_n741), .C1(new_n744), .C2(new_n717), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n716), .B1(new_n746), .B2(G1), .ZN(G364));
  INV_X1    g0547(.A(new_n698), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n253), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n206), .B1(new_n749), .B2(G45), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n711), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G330), .B2(new_n697), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n710), .A2(new_n292), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G355), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(G116), .B2(new_n228), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n672), .A2(new_n673), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n710), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n761), .B1(new_n464), .B2(new_n714), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n243), .A2(new_n464), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n757), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n226), .B1(G20), .B2(new_n335), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n752), .B1(new_n764), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n608), .A2(G200), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT96), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n774), .A2(new_n207), .A3(G190), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n528), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT32), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n207), .A2(G190), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G179), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G159), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n292), .B(new_n777), .C1(new_n778), .C2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n778), .ZN(new_n785));
  NAND3_X1  g0585(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G190), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n786), .A2(new_n347), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n788), .A2(new_n202), .B1(new_n790), .B2(new_n362), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n207), .B1(new_n780), .B2(G190), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n217), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n785), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n774), .A2(new_n207), .A3(new_n347), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G87), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n207), .A2(new_n347), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n608), .A2(G200), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n779), .A2(new_n798), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n799), .A2(new_n201), .B1(new_n800), .B2(new_n366), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT95), .Z(new_n802));
  NAND4_X1  g0602(.A1(new_n784), .A2(new_n794), .A3(new_n796), .A4(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n795), .A2(G303), .B1(new_n775), .B2(G283), .ZN(new_n804));
  INV_X1    g0604(.A(G322), .ZN(new_n805));
  INV_X1    g0605(.A(G311), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n799), .A2(new_n805), .B1(new_n800), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n781), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n286), .B(new_n807), .C1(G329), .C2(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n789), .B(KEYINPUT97), .Z(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G326), .ZN(new_n812));
  INV_X1    g0612(.A(new_n792), .ZN(new_n813));
  XNOR2_X1  g0613(.A(KEYINPUT33), .B(G317), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n813), .A2(G294), .B1(new_n787), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n804), .A2(new_n809), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n803), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n771), .B1(new_n817), .B2(new_n768), .ZN(new_n818));
  INV_X1    g0618(.A(new_n767), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n697), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n754), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  NAND2_X1  g0622(.A1(new_n661), .A2(new_n695), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n396), .A2(new_n694), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n398), .B1(new_n388), .B2(new_n695), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n396), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n823), .B(new_n827), .Z(new_n828));
  AOI21_X1  g0628(.A(new_n752), .B1(new_n828), .B2(new_n741), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n741), .B2(new_n828), .ZN(new_n830));
  INV_X1    g0630(.A(new_n768), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n799), .A2(new_n515), .B1(new_n800), .B2(new_n530), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n286), .B(new_n832), .C1(G311), .C2(new_n808), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n790), .A2(new_n461), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n793), .B(new_n834), .C1(G283), .C2(new_n787), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n795), .A2(G107), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n775), .A2(G87), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n833), .A2(new_n835), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n799), .ZN(new_n839));
  INV_X1    g0639(.A(new_n800), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G143), .A2(new_n839), .B1(new_n840), .B2(G159), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n841), .B1(new_n790), .B2(new_n842), .C1(new_n358), .C2(new_n788), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT34), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  INV_X1    g0646(.A(G132), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n759), .B1(new_n201), .B2(new_n792), .C1(new_n847), .C2(new_n781), .ZN(new_n848));
  OR3_X1    g0648(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n775), .A2(G68), .ZN(new_n850));
  INV_X1    g0650(.A(new_n795), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n851), .B2(new_n362), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT98), .Z(new_n853));
  OAI21_X1  g0653(.A(new_n838), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT99), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n831), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n855), .B2(new_n854), .ZN(new_n857));
  INV_X1    g0657(.A(new_n752), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n768), .A2(new_n765), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n858), .B1(new_n366), .B2(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n857), .B(new_n860), .C1(new_n766), .C2(new_n827), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n830), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(G384));
  NAND2_X1  g0663(.A1(new_n678), .A2(KEYINPUT16), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n313), .A2(new_n272), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n864), .A2(new_n865), .A3(new_n268), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n271), .ZN(new_n867));
  INV_X1    g0667(.A(new_n692), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n346), .B2(new_n351), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n350), .B1(new_n681), .B2(new_n337), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n681), .B2(new_n692), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT101), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT37), .B1(new_n316), .B2(new_n868), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT101), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n877), .A2(new_n878), .A3(new_n350), .A4(new_n343), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n867), .A2(new_n338), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n869), .A2(new_n881), .A3(new_n350), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT37), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n872), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n871), .A2(new_n884), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n876), .A2(new_n879), .B1(new_n882), .B2(KEYINPUT37), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n872), .B1(new_n870), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n734), .A2(new_n694), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n735), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n739), .A2(KEYINPUT31), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n624), .A2(new_n636), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n892), .A2(new_n626), .A3(new_n593), .A4(new_n695), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n889), .B(new_n890), .C1(new_n893), .C2(new_n550), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n449), .A2(new_n694), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n450), .A2(new_n454), .A3(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n449), .B(new_n694), .C1(new_n440), .C2(new_n666), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n894), .A2(new_n898), .A3(new_n827), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT103), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n885), .A2(new_n887), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n899), .A2(new_n900), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT40), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n870), .A2(new_n886), .A3(new_n872), .ZN(new_n906));
  XNOR2_X1  g0706(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n316), .A2(new_n868), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n343), .A2(new_n909), .A3(new_n350), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT37), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n880), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n316), .B(new_n868), .C1(new_n684), .C2(new_n665), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n908), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT104), .B1(new_n906), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT104), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n876), .A2(new_n879), .B1(KEYINPUT37), .B2(new_n910), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n345), .A2(new_n339), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n909), .B1(new_n918), .B2(new_n351), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n907), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n885), .A2(new_n916), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n899), .A2(new_n904), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n915), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n905), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n457), .A2(new_n894), .ZN(new_n925));
  OAI21_X1  g0725(.A(G330), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n924), .B2(new_n925), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT39), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n906), .B2(new_n914), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n450), .A2(new_n694), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n885), .A2(KEYINPUT39), .A3(new_n887), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n885), .A2(new_n887), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n896), .A2(new_n897), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n695), .B(new_n827), .C1(new_n655), .C2(new_n660), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n934), .B1(new_n824), .B2(new_n935), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n933), .A2(new_n936), .B1(new_n684), .B2(new_n692), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n932), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n718), .B1(new_n744), .B2(new_n717), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n457), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n686), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n938), .B(new_n941), .Z(new_n942));
  OAI22_X1  g0742(.A1(new_n927), .A2(new_n942), .B1(new_n206), .B2(new_n749), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n942), .B2(new_n927), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n617), .A2(KEYINPUT35), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n617), .A2(KEYINPUT35), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n226), .A2(new_n207), .A3(new_n530), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT36), .Z(new_n949));
  NOR3_X1   g0749(.A1(new_n225), .A2(new_n366), .A3(new_n280), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n950), .A2(KEYINPUT100), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n950), .A2(KEYINPUT100), .B1(new_n362), .B2(G68), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n206), .B(G13), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  OR3_X1    g0753(.A1(new_n944), .A2(new_n949), .A3(new_n953), .ZN(G367));
  AOI21_X1  g0754(.A(new_n645), .B1(new_n636), .B2(new_n656), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n955), .A2(new_n694), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT42), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n623), .A2(new_n694), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n892), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n645), .A2(new_n694), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n957), .B1(new_n708), .B2(new_n962), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n705), .A2(KEYINPUT42), .A3(new_n707), .A4(new_n961), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n956), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n584), .A2(new_n588), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n694), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n652), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n649), .B2(new_n967), .ZN(new_n969));
  XOR2_X1   g0769(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n970));
  OR3_X1    g0770(.A1(new_n965), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n965), .A2(new_n972), .B1(new_n969), .B2(new_n970), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n703), .A2(new_n961), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n971), .A2(new_n973), .B1(KEYINPUT106), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n974), .A2(KEYINPUT106), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n711), .B(KEYINPUT41), .Z(new_n979));
  AOI21_X1  g0779(.A(new_n961), .B1(new_n708), .B2(new_n701), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT107), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n980), .B1(new_n981), .B2(KEYINPUT44), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(KEYINPUT44), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT108), .Z(new_n984));
  OR2_X1    g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n708), .A2(new_n701), .A3(new_n961), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT45), .Z(new_n987));
  NAND2_X1  g0787(.A1(new_n982), .A2(new_n984), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n703), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n702), .A2(new_n706), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n708), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(new_n748), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n993), .A2(new_n746), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n985), .A2(new_n987), .A3(new_n704), .A4(new_n988), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n990), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n979), .B1(new_n996), .B2(new_n746), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n977), .B(new_n978), .C1(new_n997), .C2(new_n751), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n769), .B1(new_n228), .B2(new_n380), .C1(new_n761), .C2(new_n239), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n999), .A2(new_n752), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n776), .A2(new_n217), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(G283), .A2(new_n840), .B1(new_n808), .B2(G317), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n461), .B2(new_n799), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n759), .B1(G294), .B2(new_n787), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1004), .B(new_n1005), .C1(new_n528), .C2(new_n792), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n795), .A2(G116), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT46), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n1007), .A2(new_n1008), .B1(new_n811), .B2(G311), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n1008), .B2(new_n1007), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n795), .A2(G58), .B1(G137), .B2(new_n808), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT110), .Z(new_n1012));
  OAI22_X1  g0812(.A1(new_n788), .A2(new_n782), .B1(new_n800), .B2(new_n362), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT109), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n286), .B1(new_n792), .B2(new_n202), .C1(new_n358), .C2(new_n799), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n775), .B2(G77), .ZN(new_n1016));
  INV_X1    g0816(.A(G143), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1014), .B(new_n1016), .C1(new_n1017), .C2(new_n810), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n1006), .A2(new_n1010), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT47), .Z(new_n1020));
  OAI221_X1 g0820(.A(new_n1000), .B1(new_n819), .B2(new_n969), .C1(new_n1020), .C2(new_n831), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n998), .A2(new_n1021), .ZN(G387));
  NAND2_X1  g0822(.A1(new_n993), .A2(new_n751), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT111), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n755), .A2(new_n712), .B1(new_n528), .B2(new_n710), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n236), .A2(G45), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n381), .A2(G50), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT50), .ZN(new_n1029));
  AOI211_X1 g0829(.A(G45), .B(new_n712), .C1(G68), .C2(G77), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n761), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1026), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n858), .B1(new_n1033), .B2(new_n769), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n758), .B1(new_n252), .B2(new_n787), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n813), .A2(new_n570), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1035), .B(new_n1036), .C1(new_n782), .C2(new_n790), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n851), .A2(new_n366), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G68), .A2(new_n840), .B1(new_n808), .B2(G150), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n362), .B2(new_n799), .ZN(new_n1040));
  NOR4_X1   g0840(.A1(new_n1037), .A2(new_n1001), .A3(new_n1038), .A4(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(G283), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n851), .A2(new_n515), .B1(new_n1042), .B2(new_n792), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G317), .A2(new_n839), .B1(new_n840), .B2(G303), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n806), .B2(new_n788), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n811), .B2(G322), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1043), .B1(new_n1046), .B2(KEYINPUT48), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT112), .Z(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(KEYINPUT48), .B2(new_n1046), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1050), .A2(KEYINPUT49), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n759), .B1(G326), .B2(new_n808), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n530), .B2(new_n776), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n1050), .B2(KEYINPUT49), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1041), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1034), .B1(new_n705), .B2(new_n819), .C1(new_n1055), .C2(new_n831), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1024), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n711), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n994), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n746), .B2(new_n993), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1057), .A2(new_n1060), .ZN(G393));
  AOI21_X1  g0861(.A(KEYINPUT113), .B1(new_n989), .B2(new_n703), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n990), .A2(new_n995), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1062), .B1(new_n1063), .B2(KEYINPUT113), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n711), .B(new_n996), .C1(new_n1064), .C2(new_n994), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n962), .A2(new_n767), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n769), .B1(new_n217), .B2(new_n228), .C1(new_n761), .C2(new_n246), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n752), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n777), .B1(G283), .B2(new_n795), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n839), .A2(G311), .B1(G317), .B2(new_n789), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT52), .Z(new_n1071));
  OAI21_X1  g0871(.A(new_n292), .B1(new_n800), .B2(new_n515), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G322), .B2(new_n808), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n813), .A2(G116), .B1(G303), .B2(new_n787), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1069), .A2(new_n1071), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n839), .A2(G159), .B1(G150), .B2(new_n789), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT51), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n795), .A2(G68), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n800), .A2(new_n381), .B1(new_n781), .B2(new_n1017), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n758), .A2(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n813), .A2(G77), .B1(G50), .B2(new_n787), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n837), .A2(new_n1078), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1075), .B1(new_n1077), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1068), .B1(new_n1083), .B2(new_n768), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1064), .A2(new_n751), .B1(new_n1066), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1065), .A2(new_n1085), .ZN(G390));
  INV_X1    g0886(.A(new_n859), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n752), .B1(new_n252), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n766), .B1(new_n929), .B2(new_n931), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n795), .A2(G150), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT53), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(KEYINPUT54), .B(G143), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n800), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n286), .B1(new_n799), .B2(new_n847), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1093), .B(new_n1094), .C1(G125), .C2(new_n808), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n788), .A2(new_n842), .B1(new_n792), .B2(new_n782), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(G128), .B2(new_n789), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1095), .B(new_n1097), .C1(new_n362), .C2(new_n776), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n292), .B1(new_n799), .B2(new_n530), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(G294), .B2(new_n808), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n813), .A2(G77), .B1(G283), .B2(new_n789), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n796), .A2(new_n850), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n788), .A2(new_n528), .B1(new_n800), .B2(new_n217), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT117), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n1091), .A2(new_n1098), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1088), .B(new_n1089), .C1(new_n768), .C2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n894), .A2(new_n898), .A3(G330), .A4(new_n827), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n645), .A2(new_n593), .A3(new_n626), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n624), .B1(new_n651), .B2(new_n648), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1109), .A2(new_n643), .B1(new_n1110), .B2(KEYINPUT26), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n695), .B(new_n826), .C1(new_n1111), .C2(new_n660), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n824), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n930), .B1(new_n1113), .B2(new_n898), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n915), .A2(new_n1114), .A3(new_n921), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n935), .A2(new_n824), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n930), .B1(new_n1116), .B2(new_n898), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n929), .B2(new_n931), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1108), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n885), .A2(KEYINPUT39), .A3(new_n887), .ZN(new_n1120));
  AOI21_X1  g0920(.A(KEYINPUT39), .B1(new_n885), .B2(new_n920), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n1120), .A2(new_n1121), .B1(new_n936), .B2(new_n930), .ZN(new_n1122));
  OAI211_X1 g0922(.A(G330), .B(new_n827), .C1(new_n719), .C2(new_n740), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1123), .A2(new_n934), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n915), .A2(new_n1114), .A3(new_n921), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1122), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1119), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1106), .B1(new_n1127), .B2(new_n751), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1123), .A2(new_n934), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(KEYINPUT114), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT114), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1123), .A2(new_n934), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1130), .A2(new_n1107), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n1116), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1113), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n894), .A2(G330), .A3(new_n827), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1124), .B(new_n1135), .C1(new_n1136), .C2(new_n898), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n894), .A2(G330), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n457), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n940), .A2(new_n1140), .A3(new_n686), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT116), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1141), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1119), .A2(new_n1145), .A3(new_n1126), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n711), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n1144), .A2(new_n1127), .B1(new_n1147), .B2(KEYINPUT115), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1147), .A2(KEYINPUT115), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1128), .B1(new_n1148), .B2(new_n1149), .ZN(G378));
  XOR2_X1   g0950(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1151));
  NAND2_X1  g0951(.A1(new_n663), .A2(new_n378), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n364), .A2(new_n868), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT120), .Z(new_n1154));
  NOR2_X1   g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1151), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1157), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1151), .ZN(new_n1160));
  NOR3_X1   g0960(.A1(new_n1159), .A2(new_n1155), .A3(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n923), .A2(G330), .ZN(new_n1163));
  AOI21_X1  g0963(.A(KEYINPUT40), .B1(new_n901), .B2(new_n902), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1162), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n905), .A2(new_n1166), .A3(G330), .A4(new_n923), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n938), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1146), .A2(new_n1142), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n938), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1165), .A2(new_n1167), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT57), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1058), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n1165), .A2(new_n1167), .A3(new_n1171), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1171), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT121), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1178), .A2(new_n1179), .A3(KEYINPUT57), .A4(new_n1170), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1169), .A2(new_n1170), .A3(KEYINPUT57), .A4(new_n1172), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(KEYINPUT121), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1175), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1169), .A2(new_n751), .A3(new_n1172), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n799), .A2(KEYINPUT118), .A3(new_n528), .ZN(new_n1185));
  OAI21_X1  g0985(.A(KEYINPUT118), .B1(new_n799), .B2(new_n528), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n788), .B2(new_n217), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1185), .B(new_n1187), .C1(G116), .C2(new_n789), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n466), .B1(new_n781), .B2(new_n1042), .C1(new_n380), .C2(new_n800), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n759), .B(new_n1189), .C1(G68), .C2(new_n813), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1038), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n775), .A2(G58), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1188), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT58), .ZN(new_n1194));
  AOI21_X1  g0994(.A(G41), .B1(new_n759), .B2(G33), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1092), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n795), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n787), .A2(G132), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G128), .A2(new_n839), .B1(new_n840), .B2(G137), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n813), .A2(G150), .B1(G125), .B2(new_n789), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1201), .A2(KEYINPUT59), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(KEYINPUT59), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n775), .A2(G159), .ZN(new_n1204));
  AOI211_X1 g1004(.A(G33), .B(G41), .C1(new_n808), .C2(G124), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1194), .B1(G50), .B2(new_n1195), .C1(new_n1202), .C2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT119), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n831), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1208), .B2(new_n1207), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n858), .B1(new_n362), .B2(new_n859), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1210), .B(new_n1211), .C1(new_n1162), .C2(new_n766), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1184), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1183), .A2(new_n1213), .ZN(G375));
  NOR2_X1   g1014(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1215));
  OR3_X1    g1015(.A1(new_n1144), .A2(new_n979), .A3(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n934), .A2(new_n765), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n752), .B1(G68), .B2(new_n1087), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n799), .A2(new_n1042), .B1(new_n781), .B2(new_n461), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n286), .B(new_n1219), .C1(G107), .C2(new_n840), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n366), .B2(new_n776), .C1(new_n217), .C2(new_n851), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1036), .B1(new_n790), .B2(new_n515), .C1(new_n530), .C2(new_n788), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G50), .A2(new_n813), .B1(new_n1196), .B2(new_n787), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n759), .B(new_n1223), .C1(new_n847), .C2(new_n790), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n795), .A2(G159), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n839), .A2(G137), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G150), .A2(new_n840), .B1(new_n808), .B2(G128), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1225), .A2(new_n1192), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n1221), .A2(new_n1222), .B1(new_n1224), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1218), .B1(new_n1229), .B2(new_n768), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1138), .A2(new_n751), .B1(new_n1217), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1216), .A2(new_n1231), .ZN(G381));
  NOR2_X1   g1032(.A1(G393), .A2(G396), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n862), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT122), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1235), .A2(new_n1231), .A3(new_n1216), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n998), .A2(new_n1065), .A3(new_n1021), .A4(new_n1085), .ZN(new_n1237));
  OR4_X1    g1037(.A1(G378), .A2(new_n1236), .A3(G375), .A4(new_n1237), .ZN(G407));
  NAND2_X1  g1038(.A1(new_n693), .A2(G213), .ZN(new_n1239));
  OR3_X1    g1039(.A1(G375), .A2(G378), .A3(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(G407), .A2(G213), .A3(new_n1240), .ZN(G409));
  NAND3_X1  g1041(.A1(new_n1183), .A2(G378), .A3(new_n1213), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1184), .B(new_n1212), .C1(new_n1173), .C2(new_n979), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1243), .B(new_n1128), .C1(new_n1149), .C2(new_n1148), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(KEYINPUT123), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1143), .A2(KEYINPUT60), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1215), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1058), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT124), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1215), .A2(KEYINPUT60), .A3(new_n1143), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1250), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1231), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n862), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G384), .B(new_n1231), .C1(new_n1252), .C2(new_n1253), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT123), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1242), .A2(new_n1258), .A3(new_n1244), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1246), .A2(new_n1239), .A3(new_n1257), .A4(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT125), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1259), .A2(new_n1239), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT125), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1262), .A2(new_n1263), .A3(new_n1257), .A4(new_n1246), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT62), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1261), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT61), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n693), .A2(G213), .A3(G2897), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1255), .A2(new_n1256), .A3(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1268), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1245), .A2(new_n1239), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1267), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1265), .B1(new_n1272), .B2(new_n1257), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1266), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G393), .A2(G396), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  OR2_X1    g1078(.A1(new_n1278), .A2(new_n1233), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT127), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G387), .A2(G390), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1281), .A2(new_n1237), .A3(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1279), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1283), .A2(KEYINPUT127), .A3(new_n1284), .ZN(new_n1285));
  OR2_X1    g1085(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1286), .A2(new_n1282), .A3(new_n1237), .A4(new_n1281), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1276), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1261), .A2(new_n1264), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1272), .A2(KEYINPUT63), .A3(new_n1257), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1271), .B1(new_n1262), .B2(new_n1246), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1285), .A2(new_n1267), .A3(new_n1287), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1292), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1289), .A2(new_n1297), .ZN(G405));
  XNOR2_X1  g1098(.A(G375), .B(G378), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1299), .B(new_n1257), .ZN(new_n1300));
  XOR2_X1   g1100(.A(new_n1300), .B(new_n1288), .Z(G402));
endmodule


