//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  OAI21_X1  g035(.A(KEYINPUT67), .B1(new_n460), .B2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n460), .A2(G2104), .ZN(new_n466));
  NAND4_X1  g041(.A1(new_n461), .A2(new_n464), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(new_n466), .A3(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n465), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n463), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NOR3_X1   g051(.A1(new_n469), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT68), .ZN(G160));
  AND4_X1   g053(.A1(G2105), .A2(new_n461), .A3(new_n464), .A4(new_n466), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT69), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(new_n465), .B2(G112), .ZN(new_n482));
  OR3_X1    g057(.A1(KEYINPUT70), .A2(G100), .A3(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(KEYINPUT70), .B1(G100), .B2(G2105), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n467), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G136), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n481), .A2(new_n487), .ZN(G162));
  NOR2_X1   g063(.A1(new_n465), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(new_n479), .B2(G126), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n461), .A2(new_n464), .A3(new_n466), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n470), .A2(new_n466), .ZN(new_n497));
  NOR3_X1   g072(.A1(new_n493), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n492), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  AND2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  OR2_X1    g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n506), .A2(G543), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n508), .A2(G88), .B1(G50), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n503), .A2(new_n504), .ZN(new_n512));
  INV_X1    g087(.A(G62), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G651), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n510), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n515), .A2(new_n516), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(G166));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n509), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n506), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT73), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G51), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n508), .A2(G89), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n532), .B1(new_n505), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n505), .A2(new_n532), .A3(new_n533), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n529), .B(new_n531), .C1(new_n534), .C2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n528), .A2(new_n537), .ZN(G168));
  NAND2_X1  g113(.A1(G77), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G64), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n512), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n508), .A2(G90), .B1(new_n541), .B2(G651), .ZN(new_n542));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n526), .B2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  NAND2_X1  g120(.A1(new_n525), .A2(G43), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G651), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  OAI211_X1 g125(.A(new_n546), .B(new_n549), .C1(new_n550), .C2(new_n507), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g129(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n555));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  OR3_X1    g134(.A1(new_n523), .A2(KEYINPUT9), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT9), .B1(new_n523), .B2(new_n559), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n560), .A2(new_n561), .B1(G91), .B2(new_n508), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n505), .A2(KEYINPUT75), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n512), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n563), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  AND2_X1   g142(.A1(G78), .A2(G543), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n562), .A2(new_n569), .ZN(G299));
  OR2_X1    g145(.A1(new_n528), .A2(new_n537), .ZN(G286));
  INV_X1    g146(.A(G166), .ZN(G303));
  NAND2_X1  g147(.A1(new_n508), .A2(G87), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n509), .A2(G49), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  AOI22_X1  g151(.A1(new_n505), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(new_n548), .ZN(new_n578));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  INV_X1    g154(.A(G48), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n507), .A2(new_n579), .B1(new_n580), .B2(new_n523), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G85), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n584), .A2(new_n548), .B1(new_n585), .B2(new_n507), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(G47), .B2(new_n525), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  AND3_X1   g164(.A1(new_n505), .A2(G92), .A3(new_n506), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT10), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n564), .B2(new_n566), .ZN(new_n593));
  AND2_X1   g168(.A1(G79), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n525), .A2(G54), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n591), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n589), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n589), .B1(new_n598), .B2(G868), .ZN(G321));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(G299), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G168), .B2(new_n601), .ZN(G297));
  OAI21_X1  g178(.A(new_n602), .B1(G168), .B2(new_n601), .ZN(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n598), .B1(new_n605), .B2(G860), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT76), .ZN(G148));
  NOR2_X1   g182(.A1(new_n597), .A2(G559), .ZN(new_n608));
  OR3_X1    g183(.A1(new_n608), .A2(KEYINPUT77), .A3(new_n601), .ZN(new_n609));
  OAI21_X1  g184(.A(KEYINPUT77), .B1(new_n608), .B2(new_n601), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n609), .B(new_n610), .C1(G868), .C2(new_n552), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n497), .A2(new_n474), .ZN(new_n613));
  XNOR2_X1  g188(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT13), .Z(new_n616));
  INV_X1    g191(.A(G2100), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT80), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT82), .B(G2096), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  INV_X1    g196(.A(G111), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G2105), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n479), .A2(G123), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT81), .ZN(new_n625));
  AOI211_X1 g200(.A(new_n623), .B(new_n625), .C1(G135), .C2(new_n486), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n619), .B1(new_n620), .B2(new_n626), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n616), .A2(new_n617), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT79), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n627), .B(new_n629), .C1(new_n620), .C2(new_n626), .ZN(G156));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT84), .B(G2438), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n631), .B(new_n632), .Z(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2430), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT83), .B(KEYINPUT14), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2451), .B(G2454), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n638), .B(new_n642), .Z(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(G14), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n643), .A2(new_n644), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n646), .A2(new_n647), .ZN(G401));
  XOR2_X1   g223(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT86), .ZN(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  INV_X1    g232(.A(new_n649), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n657), .B1(new_n652), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2096), .B(G2100), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(G1971), .B(G1976), .Z(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1956), .B(G2474), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1961), .B(G1966), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n665), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n665), .A2(new_n668), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  OAI221_X1 g249(.A(new_n670), .B1(new_n665), .B2(new_n669), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(G1981), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1986), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT89), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G229));
  NOR2_X1   g259(.A1(G6), .A2(G16), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n582), .B2(G16), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT32), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1981), .ZN(new_n688));
  NAND2_X1  g263(.A1(G166), .A2(G16), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G16), .B2(G22), .ZN(new_n690));
  INV_X1    g265(.A(G1971), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G23), .ZN(new_n695));
  INV_X1    g270(.A(G288), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT33), .B(G1976), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n697), .B(new_n698), .Z(new_n699));
  NOR4_X1   g274(.A1(new_n688), .A2(new_n692), .A3(new_n693), .A4(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT34), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n694), .A2(G24), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n587), .B2(new_n694), .ZN(new_n705));
  INV_X1    g280(.A(G1986), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(G25), .A2(G29), .ZN(new_n708));
  NAND4_X1  g283(.A1(new_n461), .A2(new_n464), .A3(G2105), .A4(new_n466), .ZN(new_n709));
  INV_X1    g284(.A(G119), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n465), .A2(G107), .ZN(new_n711));
  OAI21_X1  g286(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n712));
  OAI22_X1  g287(.A1(new_n709), .A2(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n486), .B2(G131), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n708), .B1(new_n714), .B2(G29), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT35), .B(G1991), .Z(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n715), .A2(new_n717), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n707), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NOR3_X1   g295(.A1(new_n702), .A2(new_n703), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT90), .B(KEYINPUT36), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n723), .A2(KEYINPUT91), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n723), .B(KEYINPUT91), .C1(new_n725), .C2(new_n721), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT31), .B(G11), .ZN(new_n727));
  INV_X1    g302(.A(G28), .ZN(new_n728));
  OR3_X1    g303(.A1(new_n728), .A2(KEYINPUT95), .A3(KEYINPUT30), .ZN(new_n729));
  OAI21_X1  g304(.A(KEYINPUT95), .B1(new_n728), .B2(KEYINPUT30), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT30), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(G28), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n729), .B(new_n730), .C1(new_n733), .C2(KEYINPUT96), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n733), .A2(KEYINPUT96), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n727), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n626), .B2(G29), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT97), .Z(new_n738));
  NOR2_X1   g313(.A1(G168), .A2(new_n694), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n694), .B2(G21), .ZN(new_n740));
  INV_X1    g315(.A(G1966), .ZN(new_n741));
  NAND2_X1  g316(.A1(G301), .A2(G16), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n694), .A2(G5), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n740), .A2(new_n741), .B1(new_n745), .B2(G1961), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n738), .B(new_n746), .C1(new_n741), .C2(new_n740), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT98), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n731), .A2(G35), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G162), .B2(new_n731), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT29), .Z(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(G2090), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT24), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(G34), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(G34), .ZN(new_n756));
  AOI21_X1  g331(.A(G29), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G160), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(G29), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT93), .ZN(new_n760));
  INV_X1    g335(.A(G2084), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n752), .A2(G2090), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n753), .A2(new_n762), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n731), .A2(G33), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT25), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n486), .A2(G139), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n497), .A2(G127), .ZN(new_n770));
  INV_X1    g345(.A(G115), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(new_n463), .ZN(new_n772));
  AOI211_X1 g347(.A(new_n768), .B(new_n769), .C1(G2105), .C2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n766), .B1(new_n773), .B2(new_n731), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2072), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n694), .A2(G4), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n598), .B2(new_n694), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1348), .ZN(new_n778));
  INV_X1    g353(.A(G1961), .ZN(new_n779));
  AOI211_X1 g354(.A(new_n775), .B(new_n778), .C1(new_n779), .C2(new_n744), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n694), .A2(G20), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT23), .Z(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G299), .B2(G16), .ZN(new_n783));
  INV_X1    g358(.A(G1956), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n731), .A2(G26), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT28), .ZN(new_n786));
  INV_X1    g361(.A(G128), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n465), .A2(G116), .ZN(new_n788));
  OAI21_X1  g363(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n789));
  OAI22_X1  g364(.A1(new_n709), .A2(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n486), .B2(G140), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n786), .B1(new_n791), .B2(new_n731), .ZN(new_n792));
  OAI22_X1  g367(.A1(new_n783), .A2(new_n784), .B1(G2067), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n694), .A2(G19), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT92), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n552), .B2(new_n694), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1341), .ZN(new_n797));
  AOI211_X1 g372(.A(new_n793), .B(new_n797), .C1(new_n784), .C2(new_n783), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n731), .A2(G32), .ZN(new_n799));
  INV_X1    g374(.A(G141), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n467), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT94), .Z(new_n802));
  NAND3_X1  g377(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT26), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n805), .A2(new_n806), .B1(G105), .B2(new_n474), .ZN(new_n807));
  INV_X1    g382(.A(G129), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n709), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n802), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n799), .B1(new_n810), .B2(new_n731), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT27), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1996), .ZN(new_n813));
  NOR2_X1   g388(.A1(G27), .A2(G29), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G164), .B2(G29), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT99), .B(G2078), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G2067), .B2(new_n792), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n780), .A2(new_n798), .A3(new_n813), .A4(new_n818), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n748), .A2(new_n765), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n724), .A2(new_n726), .A3(new_n820), .ZN(G150));
  INV_X1    g396(.A(G150), .ZN(G311));
  AND2_X1   g397(.A1(new_n525), .A2(G55), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n824));
  INV_X1    g399(.A(G93), .ZN(new_n825));
  OAI22_X1  g400(.A1(new_n824), .A2(new_n548), .B1(new_n825), .B2(new_n507), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT101), .B(G860), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT37), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n823), .A2(new_n826), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(KEYINPUT100), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT100), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n551), .B1(new_n827), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT38), .Z(new_n836));
  NOR2_X1   g411(.A1(new_n597), .A2(new_n605), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n828), .B1(new_n839), .B2(KEYINPUT39), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n830), .B1(new_n840), .B2(new_n842), .ZN(G145));
  INV_X1    g418(.A(KEYINPUT103), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n773), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n791), .B(new_n501), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n845), .B1(new_n810), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n810), .B2(new_n846), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n773), .A2(new_n844), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n848), .B(new_n849), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n714), .B(new_n615), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n479), .A2(G130), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n465), .A2(G118), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(G142), .B2(new_n486), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n851), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n850), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n850), .A2(new_n858), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(G162), .B(KEYINPUT102), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G160), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n626), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G37), .ZN(new_n866));
  INV_X1    g441(.A(new_n864), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n859), .B2(new_n860), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT104), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n865), .A2(KEYINPUT104), .A3(new_n866), .A4(new_n868), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n871), .A2(KEYINPUT40), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT40), .B1(new_n871), .B2(new_n872), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(G395));
  NAND2_X1  g450(.A1(new_n831), .A2(new_n601), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n597), .B(G299), .Z(new_n877));
  INV_X1    g452(.A(KEYINPUT41), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n835), .B(new_n608), .ZN(new_n880));
  MUX2_X1   g455(.A(new_n877), .B(new_n879), .S(new_n880), .Z(new_n881));
  XNOR2_X1  g456(.A(G290), .B(G166), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n582), .B(G288), .Z(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n884), .B(KEYINPUT42), .Z(new_n885));
  XNOR2_X1  g460(.A(new_n881), .B(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n876), .B1(new_n886), .B2(new_n601), .ZN(G295));
  OAI21_X1  g462(.A(new_n876), .B1(new_n886), .B2(new_n601), .ZN(G331));
  XNOR2_X1  g463(.A(G168), .B(G171), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n835), .B(new_n889), .Z(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n877), .ZN(new_n891));
  INV_X1    g466(.A(new_n884), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n835), .B(new_n889), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n879), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n895), .A2(new_n866), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n891), .A2(new_n894), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n884), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT43), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n895), .A2(new_n866), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n877), .A2(KEYINPUT105), .A3(new_n878), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n893), .B(new_n902), .C1(KEYINPUT105), .C2(new_n879), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n892), .B1(new_n903), .B2(new_n891), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n900), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT44), .B1(new_n899), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n896), .A2(new_n898), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT43), .ZN(new_n908));
  OR3_X1    g483(.A1(new_n900), .A2(KEYINPUT43), .A3(new_n904), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n906), .B1(new_n910), .B2(KEYINPUT44), .ZN(G397));
  OAI21_X1  g486(.A(G8), .B1(new_n528), .B2(new_n537), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n464), .A2(new_n466), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n914), .A2(G137), .A3(new_n465), .A4(new_n461), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n471), .A2(new_n472), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(G2105), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n915), .A2(new_n917), .A3(G40), .A4(new_n475), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT45), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(G1384), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n918), .B1(new_n501), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G1384), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n495), .A2(KEYINPUT4), .B1(new_n497), .B2(new_n498), .ZN(new_n923));
  INV_X1    g498(.A(G126), .ZN(new_n924));
  OAI22_X1  g499(.A1(new_n709), .A2(new_n924), .B1(new_n489), .B2(new_n490), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n922), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n919), .ZN(new_n927));
  AOI21_X1  g502(.A(G1966), .B1(new_n921), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n477), .A2(G40), .A3(new_n761), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT50), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  XOR2_X1   g506(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n932));
  OAI211_X1 g507(.A(new_n922), .B(new_n932), .C1(new_n923), .C2(new_n925), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n929), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n913), .B1(new_n928), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT116), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT119), .ZN(new_n937));
  INV_X1    g512(.A(G8), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT45), .B1(new_n501), .B2(new_n922), .ZN(new_n939));
  INV_X1    g514(.A(G40), .ZN(new_n940));
  NOR4_X1   g515(.A1(new_n469), .A2(new_n473), .A3(new_n940), .A4(new_n476), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n920), .B1(new_n923), .B2(new_n925), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n741), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n918), .A2(G2084), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT50), .B1(new_n501), .B2(new_n922), .ZN(new_n946));
  INV_X1    g521(.A(new_n933), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n938), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT51), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n912), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n937), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(G8), .B1(new_n928), .B2(new_n934), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n953), .A2(KEYINPUT119), .A3(new_n950), .A4(new_n912), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT117), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n912), .B1(new_n949), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n953), .A2(KEYINPUT117), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT51), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT118), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n955), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI211_X1 g536(.A(KEYINPUT118), .B(KEYINPUT51), .C1(new_n957), .C2(new_n958), .ZN(new_n962));
  AOI211_X1 g537(.A(KEYINPUT120), .B(new_n936), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT120), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n959), .A2(new_n960), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n952), .A2(new_n954), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(new_n962), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n936), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT62), .B1(new_n963), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n913), .B1(new_n953), .B2(KEYINPUT117), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n949), .A2(new_n956), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n950), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n966), .B1(new_n973), .B2(KEYINPUT118), .ZN(new_n974));
  INV_X1    g549(.A(new_n962), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n968), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT120), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT62), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n967), .A2(new_n964), .A3(new_n968), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n926), .A2(new_n918), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n981), .A2(new_n938), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1976), .ZN(new_n984));
  NOR2_X1   g559(.A1(G288), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT52), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT52), .B1(G288), .B2(new_n984), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n982), .B(new_n987), .C1(new_n984), .C2(G288), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n582), .A2(new_n676), .ZN(new_n991));
  OAI21_X1  g566(.A(G1981), .B1(new_n578), .B2(new_n581), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n991), .A2(new_n992), .A3(KEYINPUT49), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT49), .B1(new_n991), .B2(new_n992), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n990), .B1(new_n995), .B2(new_n982), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n990), .A3(new_n982), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n989), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(G166), .A2(new_n938), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT55), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n691), .B1(new_n939), .B2(new_n943), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n918), .B1(new_n926), .B2(new_n932), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(KEYINPUT50), .B2(new_n926), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1003), .B1(new_n1005), .B2(G2090), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(G8), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1002), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n918), .B1(new_n931), .B2(new_n933), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1003), .B1(new_n1010), .B2(G2090), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1003), .B(KEYINPUT109), .C1(new_n1010), .C2(G2090), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1013), .A2(new_n1001), .A3(G8), .A4(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n999), .A2(new_n1008), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G2078), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n921), .A2(new_n1017), .A3(new_n927), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT121), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT121), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n921), .A2(new_n1020), .A3(new_n1017), .A4(new_n927), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1019), .A2(KEYINPUT53), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1010), .A2(new_n779), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(G171), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1016), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n970), .A2(new_n980), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT126), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n970), .A2(new_n980), .A3(KEYINPUT126), .A4(new_n1027), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n1009), .A2(G1348), .ZN(new_n1032));
  INV_X1    g607(.A(G2067), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n941), .A2(new_n922), .A3(new_n501), .A4(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n981), .A2(KEYINPUT115), .A3(new_n1033), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n597), .B1(new_n1032), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1041), .B1(new_n562), .B2(new_n569), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1005), .A2(new_n784), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT56), .B(G2072), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n921), .A2(new_n927), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT114), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n921), .A2(new_n1048), .A3(new_n927), .A4(new_n1045), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1043), .A2(new_n1044), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1039), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1044), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1043), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1009), .A2(G1348), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n597), .A2(KEYINPUT60), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1996), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n921), .A2(new_n1060), .A3(new_n927), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT58), .B(G1341), .Z(new_n1062));
  OAI21_X1  g637(.A(new_n1062), .B1(new_n926), .B2(new_n918), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT59), .B1(new_n1064), .B2(new_n552), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n1066));
  AOI211_X1 g641(.A(new_n1066), .B(new_n551), .C1(new_n1061), .C2(new_n1063), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n1059), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1056), .A2(new_n1057), .A3(new_n598), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT60), .B1(new_n1039), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1054), .A2(KEYINPUT61), .A3(new_n1050), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT61), .B1(new_n1054), .B2(new_n1050), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1055), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n942), .A2(KEYINPUT53), .A3(new_n1017), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT122), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n941), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n918), .A2(KEYINPUT122), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n927), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT123), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1077), .A2(new_n927), .A3(KEYINPUT123), .A4(new_n1078), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1075), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(G301), .A3(new_n1024), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1026), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(KEYINPUT124), .A3(new_n1024), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT124), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1018), .A2(new_n1023), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(G1961), .B2(new_n1009), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1089), .B1(new_n1091), .B2(new_n1083), .ZN(new_n1092));
  AOI21_X1  g667(.A(G301), .B1(new_n1088), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1025), .A2(G301), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT54), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1087), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1016), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1074), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1098), .B1(new_n977), .B2(new_n979), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n696), .A2(new_n984), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1100), .B1(new_n997), .B2(new_n998), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n991), .B(KEYINPUT111), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n982), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1015), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n999), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1104), .A2(KEYINPUT112), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT112), .ZN(new_n1108));
  NOR4_X1   g683(.A1(new_n983), .A2(new_n993), .A3(new_n994), .A4(KEYINPUT110), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n984), .B(new_n696), .C1(new_n996), .C2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n983), .B1(new_n1110), .B2(new_n1102), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n986), .B(new_n988), .C1(new_n996), .C2(new_n1109), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1112), .A2(new_n1015), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1108), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1107), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT63), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n949), .A2(G168), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1117), .B(KEYINPUT113), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1116), .B1(new_n1016), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1118), .A2(new_n1116), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1013), .A2(G8), .A3(new_n1014), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n1002), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1120), .A2(new_n1015), .A3(new_n999), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1115), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT125), .B1(new_n1099), .B2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1114), .A2(new_n1107), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n963), .A2(new_n969), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1127), .B(new_n1128), .C1(new_n1129), .C2(new_n1098), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1030), .A2(new_n1031), .A3(new_n1126), .A4(new_n1130), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n927), .A2(G1996), .A3(new_n918), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n810), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n1133), .B(KEYINPUT106), .Z(new_n1134));
  NOR2_X1   g709(.A1(new_n927), .A2(new_n918), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT107), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n791), .B(G2067), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n810), .B2(new_n1060), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1134), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n714), .B(new_n716), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1136), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n587), .B(new_n706), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1135), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1131), .A2(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1132), .B(KEYINPUT46), .Z(new_n1146));
  NAND2_X1  g721(.A1(new_n1137), .A2(new_n810), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1136), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  XOR2_X1   g724(.A(new_n1149), .B(KEYINPUT47), .Z(new_n1150));
  AND2_X1   g725(.A1(new_n1142), .A2(KEYINPUT127), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1142), .A2(KEYINPUT127), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1135), .A2(new_n706), .A3(new_n587), .ZN(new_n1153));
  XOR2_X1   g728(.A(new_n1153), .B(KEYINPUT48), .Z(new_n1154));
  NOR3_X1   g729(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1139), .A2(new_n714), .A3(new_n716), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n791), .A2(new_n1033), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AOI211_X1 g733(.A(new_n1150), .B(new_n1155), .C1(new_n1136), .C2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1145), .A2(new_n1159), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g735(.A(G319), .B1(new_n646), .B2(new_n647), .ZN(new_n1162));
  NOR2_X1   g736(.A1(new_n1162), .A2(G227), .ZN(new_n1163));
  NAND2_X1  g737(.A1(new_n683), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g738(.A(new_n1164), .B1(new_n908), .B2(new_n909), .ZN(new_n1165));
  NAND2_X1  g739(.A1(new_n871), .A2(new_n872), .ZN(new_n1166));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n1166), .ZN(G225));
  INV_X1    g741(.A(G225), .ZN(G308));
endmodule


