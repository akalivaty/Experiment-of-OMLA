//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  AND2_X1   g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G20), .ZN(new_n217));
  INV_X1    g0017(.A(new_n201), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT64), .B(G77), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G116), .A2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n212), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n215), .B1(new_n217), .B2(new_n219), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  XNOR2_X1  g0047(.A(KEYINPUT3), .B(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(G222), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(G1698), .ZN(new_n251));
  INV_X1    g0051(.A(G223), .ZN(new_n252));
  OAI221_X1 g0052(.A(new_n250), .B1(new_n220), .B2(new_n248), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G1), .A2(G13), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n254), .B1(G33), .B2(G41), .ZN(new_n255));
  AND2_X1   g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G41), .ZN(new_n257));
  INV_X1    g0057(.A(G45), .ZN(new_n258));
  AOI21_X1  g0058(.A(G1), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G226), .ZN(new_n261));
  INV_X1    g0061(.A(new_n259), .ZN(new_n262));
  INV_X1    g0062(.A(G274), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n263), .B1(new_n216), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n261), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n256), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n254), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT8), .B(G58), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT67), .ZN(new_n274));
  INV_X1    g0074(.A(G58), .ZN(new_n275));
  OR3_X1    g0075(.A1(new_n275), .A2(KEYINPUT67), .A3(KEYINPUT8), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n210), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n272), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G13), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n285), .A2(new_n210), .A3(G1), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n202), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n271), .B1(new_n209), .B2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n287), .B1(new_n289), .B2(new_n202), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n269), .A2(G200), .B1(new_n291), .B2(KEYINPUT9), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n268), .A2(G190), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n292), .B(new_n293), .C1(KEYINPUT9), .C2(new_n291), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT10), .ZN(new_n295));
  INV_X1    g0095(.A(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT3), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT3), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G33), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n297), .A2(new_n299), .A3(G232), .A4(G1698), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n297), .A2(new_n299), .A3(G226), .A4(new_n249), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G97), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n255), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n260), .A2(G238), .B1(new_n259), .B2(new_n265), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT13), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n306), .B1(new_n304), .B2(new_n305), .ZN(new_n309));
  OAI21_X1  g0109(.A(G169), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT69), .B(KEYINPUT14), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n304), .A2(new_n305), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT13), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n307), .ZN(new_n315));
  INV_X1    g0115(.A(G179), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n310), .A2(new_n312), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(new_n314), .B2(new_n307), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT14), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT68), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT68), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n310), .A2(new_n322), .A3(KEYINPUT14), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n317), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n282), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n325), .A2(new_n202), .B1(new_n210), .B2(G68), .ZN(new_n326));
  INV_X1    g0126(.A(G77), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n279), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n271), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT11), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n286), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n333), .A2(KEYINPUT12), .A3(G68), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT12), .ZN(new_n335));
  INV_X1    g0135(.A(G68), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n335), .B1(new_n286), .B2(new_n336), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n334), .A2(new_n337), .B1(new_n289), .B2(new_n336), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n329), .A2(new_n330), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n332), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n324), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n308), .A2(new_n309), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G190), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n315), .A2(G200), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n343), .A2(new_n344), .A3(new_n340), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n269), .A2(G179), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n268), .A2(G169), .B1(new_n284), .B2(new_n290), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n289), .A2(new_n327), .B1(new_n221), .B2(new_n333), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT15), .B(G87), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n221), .A2(G20), .B1(new_n354), .B2(new_n280), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n325), .B2(new_n273), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n352), .B1(new_n356), .B2(new_n271), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n248), .A2(G232), .A3(new_n249), .ZN(new_n358));
  INV_X1    g0158(.A(G238), .ZN(new_n359));
  OAI221_X1 g0159(.A(new_n358), .B1(new_n206), .B2(new_n248), .C1(new_n251), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n255), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n260), .A2(G244), .B1(new_n259), .B2(new_n265), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n357), .B1(new_n363), .B2(new_n318), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(G179), .B2(new_n363), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(G200), .ZN(new_n366));
  INV_X1    g0166(.A(G190), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n366), .B(new_n357), .C1(new_n367), .C2(new_n363), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n295), .A2(new_n347), .A3(new_n351), .A4(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT17), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n298), .A2(G33), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n296), .A2(KEYINPUT3), .ZN(new_n374));
  OAI211_X1 g0174(.A(KEYINPUT7), .B(new_n210), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT70), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n248), .B2(G20), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n297), .A2(new_n299), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT70), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n379), .A2(new_n380), .A3(KEYINPUT7), .A4(new_n210), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n376), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G68), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n275), .A2(new_n336), .ZN(new_n384));
  OAI21_X1  g0184(.A(G20), .B1(new_n384), .B2(new_n201), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n282), .A2(G159), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n383), .A2(KEYINPUT16), .A3(new_n388), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n248), .A2(new_n377), .A3(G20), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT7), .B1(new_n379), .B2(new_n210), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n388), .B1(new_n392), .B2(new_n336), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n389), .A2(new_n395), .A3(new_n271), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n277), .A2(new_n288), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(new_n277), .B2(new_n333), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n297), .A2(new_n299), .A3(G226), .A4(G1698), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n297), .A2(new_n299), .A3(G223), .A4(new_n249), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G87), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n255), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n260), .A2(G232), .B1(new_n259), .B2(new_n265), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT71), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT71), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G200), .ZN(new_n412));
  INV_X1    g0212(.A(new_n407), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n411), .A2(new_n412), .B1(new_n367), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n372), .B1(new_n400), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(KEYINPUT72), .A2(KEYINPUT18), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n387), .B1(new_n382), .B2(G68), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n272), .B1(new_n417), .B2(KEYINPUT16), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n398), .B1(new_n418), .B2(new_n395), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT71), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT71), .B1(new_n405), .B2(new_n406), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n318), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n413), .A2(new_n316), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n416), .B1(new_n419), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n412), .B1(new_n420), .B2(new_n421), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(G190), .B2(new_n407), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n419), .A2(new_n427), .A3(KEYINPUT17), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n415), .A2(new_n425), .A3(new_n428), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n419), .A2(KEYINPUT18), .A3(new_n424), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT18), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n411), .A2(new_n318), .B1(new_n316), .B2(new_n413), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n431), .B1(new_n400), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT72), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n371), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n359), .A2(G1698), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n438), .A2(new_n297), .A3(new_n299), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT76), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G116), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n297), .A2(new_n299), .A3(G244), .A4(G1698), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n438), .A2(new_n297), .A3(new_n299), .A4(KEYINPUT76), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n441), .A2(new_n442), .A3(new_n443), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n255), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n258), .A2(G1), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n265), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n216), .A2(new_n264), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n209), .A2(G45), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(G250), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n446), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n318), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n452), .B1(new_n445), .B2(new_n255), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n316), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n248), .A2(new_n210), .A3(G68), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT19), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n210), .B1(new_n302), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(G87), .B2(new_n207), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n459), .B1(new_n279), .B2(new_n205), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n458), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n463), .A2(new_n271), .B1(new_n286), .B2(new_n353), .ZN(new_n464));
  XOR2_X1   g0264(.A(new_n353), .B(KEYINPUT77), .Z(new_n465));
  NAND2_X1  g0265(.A1(new_n209), .A2(G33), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n333), .A2(new_n272), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n455), .A2(new_n457), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(G87), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n464), .B(new_n471), .C1(new_n456), .C2(new_n412), .ZN(new_n472));
  OR2_X1    g0272(.A1(new_n472), .A2(KEYINPUT78), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n454), .A2(new_n367), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n474), .B1(new_n472), .B2(KEYINPUT78), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n470), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  OR2_X1    g0276(.A1(KEYINPUT5), .A2(G41), .ZN(new_n477));
  NAND2_X1  g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n450), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n265), .ZN(new_n480));
  INV_X1    g0280(.A(new_n478), .ZN(new_n481));
  NOR2_X1   g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n447), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n449), .ZN(new_n484));
  INV_X1    g0284(.A(G257), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n480), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n297), .A2(new_n299), .A3(G244), .A4(new_n249), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n248), .A2(KEYINPUT4), .A3(G244), .A4(new_n249), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G283), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n248), .A2(G250), .A3(G1698), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n489), .A2(new_n490), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n486), .B1(new_n255), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n316), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n378), .A2(new_n375), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n496), .A2(G107), .B1(G77), .B2(new_n282), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G97), .A2(G107), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT6), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT73), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT73), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT6), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT74), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(G97), .B1(new_n500), .B2(new_n502), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n207), .B(new_n498), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n207), .A2(new_n498), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n506), .A2(G20), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n272), .B1(new_n497), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n286), .A2(new_n205), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n333), .A2(new_n272), .A3(new_n466), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(new_n205), .ZN(new_n514));
  OAI221_X1 g0314(.A(new_n495), .B1(G169), .B2(new_n494), .C1(new_n511), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n493), .A2(new_n255), .ZN(new_n516));
  INV_X1    g0316(.A(new_n486), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G200), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n497), .A2(new_n510), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n271), .ZN(new_n521));
  INV_X1    g0321(.A(new_n514), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n494), .A2(G190), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n519), .A2(new_n521), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT75), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n515), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n476), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT80), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(G294), .ZN(new_n529));
  INV_X1    g0329(.A(G294), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(KEYINPUT80), .ZN(new_n531));
  OAI21_X1  g0331(.A(G33), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n297), .A2(new_n299), .A3(G257), .A4(G1698), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n297), .A2(new_n299), .A3(G250), .A4(new_n249), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n255), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n479), .A2(new_n255), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G264), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n538), .A3(new_n480), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n412), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n255), .A2(new_n535), .B1(new_n537), .B2(G264), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(new_n367), .A3(new_n480), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n542), .A3(KEYINPUT81), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT81), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n539), .A2(new_n544), .A3(new_n412), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n297), .A2(new_n299), .A3(new_n210), .A4(G87), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT22), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT22), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n248), .A2(new_n548), .A3(new_n210), .A4(G87), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT24), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n442), .A2(G20), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT23), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n210), .B2(G107), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n552), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n550), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n551), .B1(new_n550), .B2(new_n556), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n271), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n286), .A2(new_n206), .ZN(new_n560));
  XOR2_X1   g0360(.A(KEYINPUT79), .B(KEYINPUT25), .Z(new_n561));
  XNOR2_X1  g0361(.A(new_n560), .B(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n562), .B1(G107), .B2(new_n467), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n543), .A2(new_n545), .A3(new_n559), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n559), .A2(new_n563), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n539), .A2(G179), .ZN(new_n566));
  AOI21_X1  g0366(.A(G169), .B1(new_n541), .B2(new_n480), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n515), .A2(new_n524), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n570), .B1(KEYINPUT75), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT21), .ZN(new_n573));
  INV_X1    g0373(.A(G116), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n270), .A2(new_n254), .B1(G20), .B2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n491), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n575), .A2(KEYINPUT20), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(KEYINPUT20), .B1(new_n575), .B2(new_n576), .ZN(new_n578));
  OR2_X1    g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n286), .A2(new_n574), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n467), .A2(G116), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n483), .A2(G270), .A3(new_n449), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n480), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n297), .A2(new_n299), .A3(G264), .A4(G1698), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n297), .A2(new_n299), .A3(G257), .A4(new_n249), .ZN(new_n588));
  INV_X1    g0388(.A(G303), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n587), .B(new_n588), .C1(new_n589), .C2(new_n248), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n255), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G169), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n573), .B1(new_n583), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n582), .B1(G200), .B2(new_n592), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n367), .B2(new_n592), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n586), .A2(new_n591), .A3(G179), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n582), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n582), .A2(new_n592), .A3(KEYINPUT21), .A4(G169), .ZN(new_n599));
  AND4_X1   g0399(.A1(new_n594), .A2(new_n596), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n527), .A2(new_n572), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n437), .A2(new_n601), .ZN(G372));
  NOR2_X1   g0402(.A1(new_n430), .A2(new_n433), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n346), .A2(new_n365), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n341), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n415), .B(new_n428), .C1(new_n605), .C2(KEYINPUT83), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n605), .A2(KEYINPUT83), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n603), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n350), .B1(new_n608), .B2(new_n295), .ZN(new_n609));
  INV_X1    g0409(.A(new_n515), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n476), .A2(KEYINPUT26), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n472), .ZN(new_n612));
  INV_X1    g0412(.A(new_n474), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n454), .A2(new_n318), .B1(new_n464), .B2(new_n468), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n612), .A2(new_n613), .B1(new_n614), .B2(new_n457), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT26), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n611), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n470), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n515), .A2(new_n524), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n621), .A2(new_n564), .A3(new_n615), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n594), .A2(new_n598), .A3(new_n599), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT82), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n569), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n565), .A2(new_n568), .A3(KEYINPUT82), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n620), .B1(new_n622), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n436), .B1(new_n619), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n609), .A2(new_n629), .ZN(G369));
  NAND3_X1  g0430(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n631), .A2(KEYINPUT27), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(KEYINPUT27), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(G213), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(G343), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n583), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n623), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n623), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n596), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n639), .B1(new_n641), .B2(new_n638), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G330), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n565), .A2(new_n636), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n564), .A2(new_n569), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT84), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT84), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n564), .A2(new_n569), .A3(new_n644), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n569), .A2(new_n637), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n643), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n626), .ZN(new_n654));
  AOI21_X1  g0454(.A(KEYINPUT82), .B1(new_n565), .B2(new_n568), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n654), .A2(new_n655), .A3(new_n636), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n623), .A2(new_n637), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n656), .B1(new_n649), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n653), .A2(new_n659), .ZN(G399));
  INV_X1    g0460(.A(new_n213), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(G41), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(G1), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n219), .B2(new_n663), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT28), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT88), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n456), .A2(new_n541), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n516), .A2(KEYINPUT30), .A3(new_n517), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n669), .A2(new_n670), .A3(KEYINPUT85), .A4(new_n597), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT85), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n585), .B1(new_n255), .B2(new_n590), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n673), .A2(new_n456), .A3(G179), .A4(new_n541), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n494), .A2(KEYINPUT30), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n673), .A2(new_n456), .A3(G179), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n494), .B1(new_n541), .B2(new_n480), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n671), .A2(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT30), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n674), .B2(new_n518), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(KEYINPUT31), .A3(new_n636), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n671), .A2(new_n676), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n681), .A2(KEYINPUT86), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n678), .A2(new_n677), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n597), .A2(new_n541), .A3(new_n494), .A4(new_n456), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT86), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(new_n688), .A3(new_n680), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n684), .A2(new_n685), .A3(new_n686), .A4(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT31), .B1(new_n690), .B2(new_n636), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT87), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n683), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AOI211_X1 g0493(.A(KEYINPUT87), .B(KEYINPUT31), .C1(new_n690), .C2(new_n636), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n668), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n689), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n688), .B1(new_n687), .B2(new_n680), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n637), .B1(new_n698), .B2(new_n679), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT87), .B1(new_n699), .B2(KEYINPUT31), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n691), .A2(new_n692), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n700), .A2(new_n701), .A3(KEYINPUT88), .A4(new_n683), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n527), .A2(new_n572), .A3(new_n600), .A4(new_n637), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n695), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT89), .ZN(new_n706));
  AND4_X1   g0506(.A1(new_n564), .A2(new_n615), .A3(new_n515), .A4(new_n524), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n640), .B1(new_n654), .B2(new_n655), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n470), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n611), .A2(new_n618), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n636), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n706), .B1(new_n711), .B2(KEYINPUT29), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n637), .B1(new_n619), .B2(new_n628), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT29), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(KEYINPUT89), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n569), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n707), .B1(new_n716), .B2(new_n623), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n476), .A2(new_n617), .A3(new_n610), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n470), .B1(new_n616), .B2(KEYINPUT26), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n720), .A2(KEYINPUT29), .A3(new_n637), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n712), .A2(new_n715), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n705), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n667), .B1(new_n724), .B2(G1), .ZN(G364));
  AOI21_X1  g0525(.A(new_n254), .B1(G20), .B2(new_n318), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n210), .A2(new_n316), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n729), .A2(G190), .A3(G200), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n731), .A2(KEYINPUT91), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(KEYINPUT91), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n221), .ZN(new_n736));
  NOR4_X1   g0536(.A1(new_n210), .A2(new_n412), .A3(G179), .A4(G190), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n206), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n728), .A2(G190), .A3(new_n412), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n379), .B1(new_n742), .B2(G58), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G179), .A2(G200), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(G20), .A3(new_n367), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G159), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n728), .A2(G200), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n367), .ZN(new_n749));
  AOI22_X1  g0549(.A1(KEYINPUT32), .A2(new_n747), .B1(new_n749), .B2(G50), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n736), .A2(new_n740), .A3(new_n743), .A4(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n748), .A2(G190), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n210), .B1(new_n744), .B2(G190), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n752), .A2(G68), .B1(G97), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G87), .ZN(new_n756));
  NOR4_X1   g0556(.A1(new_n210), .A2(new_n367), .A3(new_n412), .A4(G179), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n755), .B1(KEYINPUT32), .B2(new_n747), .C1(new_n756), .C2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G317), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(KEYINPUT33), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n760), .A2(KEYINPUT33), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n752), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n529), .A2(new_n531), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n763), .B1(new_n589), .B2(new_n758), .C1(new_n764), .C2(new_n753), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n730), .A2(G311), .B1(new_n742), .B2(G322), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n749), .A2(G326), .B1(G283), .B2(new_n737), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n248), .B1(new_n746), .B2(G329), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n751), .A2(new_n759), .B1(new_n765), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT92), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n727), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n771), .B2(new_n770), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n285), .A2(G20), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n209), .B1(new_n774), .B2(G45), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n662), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n213), .A2(new_n248), .ZN(new_n778));
  INV_X1    g0578(.A(G355), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n778), .A2(new_n779), .B1(G116), .B2(new_n213), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n661), .A2(new_n248), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n219), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n782), .B1(new_n258), .B2(new_n783), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n246), .A2(new_n258), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n780), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G13), .A2(G33), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(G20), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n726), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n777), .B1(new_n786), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT90), .ZN(new_n793));
  INV_X1    g0593(.A(new_n789), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n773), .B(new_n793), .C1(new_n642), .C2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n642), .A2(G330), .ZN(new_n796));
  INV_X1    g0596(.A(new_n777), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n643), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n795), .B1(new_n796), .B2(new_n798), .ZN(G396));
  INV_X1    g0599(.A(new_n705), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n368), .B1(new_n357), .B2(new_n637), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n365), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n365), .B2(new_n636), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT93), .ZN(new_n804));
  MUX2_X1   g0604(.A(new_n804), .B(new_n803), .S(new_n711), .Z(new_n805));
  NOR2_X1   g0605(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n806), .A2(KEYINPUT94), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(KEYINPUT94), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n777), .B1(new_n800), .B2(new_n805), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n726), .A2(new_n787), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n797), .B1(new_n327), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n752), .ZN(new_n813));
  INV_X1    g0613(.A(G283), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n813), .A2(new_n814), .B1(new_n206), .B2(new_n758), .ZN(new_n815));
  INV_X1    g0615(.A(G311), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n379), .B1(new_n745), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G294), .B2(new_n742), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n754), .A2(G97), .B1(new_n737), .B2(G87), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n818), .B(new_n819), .C1(new_n734), .C2(new_n574), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n815), .B(new_n820), .C1(G303), .C2(new_n749), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n379), .B1(new_n746), .B2(G132), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n275), .B2(new_n753), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n758), .A2(new_n202), .B1(new_n738), .B2(new_n336), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G137), .A2(new_n749), .B1(new_n742), .B2(G143), .ZN(new_n825));
  INV_X1    g0625(.A(G150), .ZN(new_n826));
  INV_X1    g0626(.A(G159), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n825), .B1(new_n826), .B2(new_n813), .C1(new_n734), .C2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT34), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n823), .B(new_n824), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n821), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n803), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n812), .B1(new_n832), .B2(new_n727), .C1(new_n833), .C2(new_n788), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n810), .A2(new_n834), .ZN(G384));
  NOR3_X1   g0635(.A1(new_n219), .A2(new_n220), .A3(new_n384), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n202), .B2(G68), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n837), .A2(new_n209), .A3(G13), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT96), .Z(new_n839));
  NOR2_X1   g0639(.A1(new_n217), .A2(new_n574), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n506), .A2(new_n509), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT35), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n842), .B2(new_n841), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT95), .Z(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n839), .B1(new_n846), .B2(KEYINPUT36), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n341), .A2(new_n637), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n417), .A2(KEYINPUT16), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n398), .B1(new_n850), .B2(new_n418), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n851), .A2(new_n634), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT72), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT18), .B1(new_n419), .B2(new_n424), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n400), .A2(new_n431), .A3(new_n432), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n415), .A2(new_n425), .A3(new_n428), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n852), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n634), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n422), .B2(new_n423), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n851), .A2(new_n860), .B1(new_n400), .B2(new_n414), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n400), .A2(new_n432), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n400), .A2(new_n859), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n419), .A2(new_n427), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n863), .A2(new_n864), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n858), .A2(KEYINPUT38), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT38), .B1(new_n858), .B2(new_n868), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT39), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT98), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n858), .A2(KEYINPUT38), .A3(new_n868), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT39), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT37), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n415), .A2(new_n854), .A3(new_n855), .A4(new_n428), .ZN(new_n877));
  INV_X1    g0677(.A(new_n864), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n876), .A2(new_n867), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n873), .B(new_n874), .C1(KEYINPUT38), .C2(new_n879), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n871), .A2(new_n872), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n872), .B1(new_n871), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n849), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n365), .A2(new_n636), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n884), .B(KEYINPUT97), .Z(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n713), .B2(new_n803), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n340), .A2(new_n637), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n345), .B(new_n889), .C1(new_n324), .C2(new_n340), .ZN(new_n890));
  INV_X1    g0690(.A(new_n340), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n319), .A2(new_n311), .B1(new_n342), .B2(G179), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n319), .A2(KEYINPUT68), .A3(new_n320), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n322), .B1(new_n310), .B2(KEYINPUT14), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n891), .B(new_n636), .C1(new_n895), .C2(new_n346), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n887), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n869), .A2(new_n870), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n898), .A2(new_n899), .B1(new_n603), .B2(new_n859), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n883), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n436), .A2(new_n712), .A3(new_n715), .A4(new_n721), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n609), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n902), .B(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n897), .A2(new_n833), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT40), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n690), .A2(new_n636), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n909), .A2(KEYINPUT99), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT99), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n690), .B2(new_n636), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n910), .A2(KEYINPUT31), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n690), .A2(KEYINPUT31), .A3(new_n636), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n703), .A2(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n907), .B(new_n908), .C1(new_n913), .C2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n916), .A2(new_n899), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n703), .A2(new_n914), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n912), .A2(KEYINPUT31), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n699), .A2(new_n911), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n906), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n873), .B1(KEYINPUT38), .B2(new_n879), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n908), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n913), .A2(new_n915), .ZN(new_n926));
  OR3_X1    g0726(.A1(new_n925), .A2(new_n437), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n925), .B1(new_n437), .B2(new_n926), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n927), .A2(new_n928), .A3(G330), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n905), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n209), .B2(new_n774), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n905), .A2(new_n929), .ZN(new_n932));
  OAI221_X1 g0732(.A(new_n847), .B1(KEYINPUT36), .B2(new_n846), .C1(new_n931), .C2(new_n932), .ZN(G367));
  NAND2_X1  g0733(.A1(new_n757), .A2(G116), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT46), .Z(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n735), .B2(G283), .ZN(new_n936));
  INV_X1    g0736(.A(new_n749), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n937), .A2(new_n816), .B1(new_n589), .B2(new_n741), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT107), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n379), .B1(new_n745), .B2(new_n760), .C1(new_n813), .C2(new_n764), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n738), .A2(new_n205), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(G107), .B2(new_n754), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n936), .A2(new_n939), .A3(new_n941), .A4(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT108), .ZN(new_n945));
  INV_X1    g0745(.A(G137), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n248), .B1(new_n745), .B2(new_n946), .C1(new_n741), .C2(new_n826), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n813), .A2(new_n827), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n947), .B(new_n948), .C1(G143), .C2(new_n749), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n753), .A2(new_n336), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n738), .A2(new_n220), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n950), .B(new_n951), .C1(G58), .C2(new_n757), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n949), .B(new_n952), .C1(new_n202), .C2(new_n734), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n945), .A2(new_n953), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n954), .A2(KEYINPUT47), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(KEYINPUT47), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n955), .A2(new_n726), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n781), .A2(new_n239), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n791), .B1(new_n661), .B2(new_n354), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n797), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n464), .A2(new_n471), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n636), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n615), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n620), .B2(new_n962), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n957), .B(new_n960), .C1(new_n794), .C2(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n966));
  OAI21_X1  g0766(.A(new_n636), .B1(new_n511), .B2(new_n514), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n621), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT100), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n515), .B2(new_n637), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n494), .A2(G169), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(new_n521), .B2(new_n522), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n972), .A2(KEYINPUT100), .A3(new_n495), .A4(new_n636), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n968), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n966), .B1(new_n659), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n657), .B1(new_n646), .B2(new_n648), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n621), .A2(new_n967), .B1(new_n970), .B2(new_n973), .ZN(new_n978));
  INV_X1    g0778(.A(new_n966), .ZN(new_n979));
  NOR4_X1   g0779(.A1(new_n977), .A2(new_n978), .A3(new_n656), .A4(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT44), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n659), .B2(new_n975), .ZN(new_n983));
  OAI211_X1 g0783(.A(KEYINPUT44), .B(new_n978), .C1(new_n977), .C2(new_n656), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n653), .B1(new_n981), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n981), .A2(new_n653), .A3(new_n985), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(KEYINPUT106), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT106), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n981), .A2(new_n985), .A3(new_n989), .A4(new_n653), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n986), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n651), .A2(new_n657), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n649), .A2(new_n658), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n643), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n992), .A2(new_n643), .A3(new_n993), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n705), .A2(new_n722), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(KEYINPUT105), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT105), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n705), .A2(new_n722), .A3(new_n998), .A4(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n991), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n724), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n662), .B(KEYINPUT41), .Z(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n776), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n515), .B1(new_n978), .B2(new_n569), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n637), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n977), .A2(new_n975), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(KEYINPUT42), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT101), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1009), .A2(new_n1011), .A3(KEYINPUT101), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1014), .B(new_n1015), .C1(KEYINPUT42), .C2(new_n1010), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT103), .Z(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1016), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n652), .A2(new_n975), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT102), .Z(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1022), .A2(new_n1026), .A3(new_n1023), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n965), .B1(new_n1007), .B2(new_n1030), .ZN(G387));
  INV_X1    g0831(.A(new_n998), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n723), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n662), .B(KEYINPUT110), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n999), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n651), .A2(new_n789), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n778), .A2(new_n664), .B1(G107), .B2(new_n213), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n236), .A2(G45), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n664), .ZN(new_n1039));
  AOI211_X1 g0839(.A(G45), .B(new_n1039), .C1(G68), .C2(G77), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n273), .A2(G50), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT50), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n782), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1037), .B1(new_n1038), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n777), .B1(new_n1044), .B2(new_n791), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT109), .Z(new_n1046));
  AOI22_X1  g0846(.A1(G311), .A2(new_n752), .B1(new_n742), .B2(G317), .ZN(new_n1047));
  INV_X1    g0847(.A(G322), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1047), .B1(new_n1048), .B2(new_n937), .C1(new_n734), .C2(new_n589), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT48), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n758), .A2(new_n764), .B1(new_n814), .B2(new_n753), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n1050), .B2(new_n1049), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT49), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n738), .A2(new_n574), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n248), .B(new_n1058), .C1(G326), .C2(new_n746), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1056), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n731), .A2(new_n336), .B1(new_n202), .B2(new_n741), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n379), .B(new_n1061), .C1(G150), .C2(new_n746), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n758), .A2(new_n220), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n942), .B(new_n1063), .C1(new_n749), .C2(G159), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n278), .A2(new_n752), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n465), .A2(new_n754), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1062), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1060), .A2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1036), .B(new_n1046), .C1(new_n1068), .C2(new_n727), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1035), .B(new_n1069), .C1(new_n775), .C2(new_n1032), .ZN(G393));
  AOI22_X1  g0870(.A1(G317), .A2(new_n749), .B1(new_n742), .B2(G311), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT52), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n379), .B1(new_n745), .B2(new_n1048), .C1(new_n731), .C2(new_n530), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n740), .B1(new_n589), .B2(new_n813), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n758), .A2(new_n814), .B1(new_n574), .B2(new_n753), .ZN(new_n1075));
  OR4_X1    g0875(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n813), .A2(new_n202), .B1(new_n753), .B2(new_n327), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n379), .B(new_n1077), .C1(G87), .C2(new_n737), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n757), .A2(G68), .B1(new_n746), .B2(G143), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT112), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1078), .B(new_n1080), .C1(new_n273), .C2(new_n734), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G150), .A2(new_n749), .B1(new_n742), .B2(G159), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT51), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1076), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n726), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n781), .A2(new_n243), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n791), .B1(G97), .B2(new_n661), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n797), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n789), .B2(new_n978), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n983), .A2(new_n984), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n656), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n993), .A2(new_n1092), .A3(new_n975), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n979), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n659), .A2(new_n975), .A3(new_n966), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n652), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT111), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n986), .A2(KEYINPUT111), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1099), .A2(new_n1100), .B1(new_n988), .B2(new_n990), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1090), .B1(new_n1101), .B2(new_n776), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n999), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1034), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1003), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1102), .B1(new_n1104), .B2(new_n1105), .ZN(G390));
  NAND2_X1  g0906(.A1(new_n876), .A2(new_n867), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n877), .A2(new_n878), .ZN(new_n1108));
  AOI21_X1  g0908(.A(KEYINPUT38), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n869), .A2(KEYINPUT39), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT38), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n852), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n429), .B2(new_n434), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n862), .A2(new_n867), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1111), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n874), .B1(new_n1115), .B2(new_n873), .ZN(new_n1116));
  OAI21_X1  g0916(.A(KEYINPUT98), .B1(new_n1110), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n871), .A2(new_n872), .A3(new_n880), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n885), .B1(new_n711), .B2(new_n833), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n890), .A2(new_n896), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n848), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1117), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n720), .A2(new_n637), .A3(new_n833), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n886), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n897), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n848), .B(KEYINPUT113), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1125), .A2(new_n923), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(G330), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n926), .A2(new_n1129), .A3(new_n906), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n704), .A2(G330), .A3(new_n833), .A4(new_n897), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1122), .A2(new_n1127), .A3(new_n1132), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n776), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1117), .A2(new_n1118), .A3(new_n787), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n811), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n777), .B1(new_n278), .B2(new_n1137), .ZN(new_n1138));
  XOR2_X1   g0938(.A(KEYINPUT54), .B(G143), .Z(new_n1139));
  NAND2_X1  g0939(.A1(new_n735), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n757), .A2(G150), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT53), .Z(new_n1142));
  OAI22_X1  g0942(.A1(new_n738), .A2(new_n202), .B1(new_n827), .B2(new_n753), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n813), .A2(new_n946), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(G128), .C2(new_n749), .ZN(new_n1145));
  INV_X1    g0945(.A(G125), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n248), .B1(new_n745), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(G132), .B2(new_n742), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1140), .A2(new_n1142), .A3(new_n1145), .A4(new_n1148), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n734), .A2(new_n205), .B1(new_n206), .B2(new_n813), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(KEYINPUT114), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n937), .A2(new_n814), .B1(new_n753), .B2(new_n327), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n758), .A2(new_n756), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n738), .A2(new_n336), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n379), .B1(new_n745), .B2(new_n530), .C1(new_n741), .C2(new_n574), .ZN(new_n1155));
  NOR4_X1   g0955(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1151), .A2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1150), .A2(KEYINPUT114), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1149), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1138), .B1(new_n1159), .B2(new_n726), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1136), .A2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n926), .A2(new_n1129), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n436), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1163), .A2(new_n609), .A3(new_n903), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n704), .A2(G330), .A3(new_n833), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n1120), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1130), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n887), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n804), .B(G330), .C1(new_n913), .C2(new_n915), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1124), .B1(new_n1170), .B2(new_n1120), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n1132), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1164), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1134), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1164), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1130), .B1(new_n1165), .B2(new_n1120), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1172), .B1(new_n1176), .B2(new_n1119), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1131), .A2(new_n1133), .A3(new_n1175), .A4(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n1034), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1135), .B(new_n1161), .C1(new_n1174), .C2(new_n1179), .ZN(G378));
  NAND2_X1  g0980(.A1(new_n295), .A2(new_n351), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n291), .A2(new_n634), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1181), .B(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1183), .B(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n848), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n907), .B1(new_n913), .B2(new_n915), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n869), .A2(new_n1109), .ZN(new_n1189));
  OAI21_X1  g0989(.A(KEYINPUT40), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1115), .A2(new_n873), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n922), .A2(new_n908), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1129), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1187), .A2(new_n1193), .A3(new_n900), .ZN(new_n1194));
  OAI21_X1  g0994(.A(G330), .B1(new_n917), .B2(new_n924), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n883), .B2(new_n901), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1186), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1193), .B1(new_n1187), .B2(new_n900), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n883), .A2(new_n901), .A3(new_n1195), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1198), .A2(new_n1199), .A3(new_n1185), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n776), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n248), .A2(G41), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n937), .A2(new_n574), .B1(new_n275), .B2(new_n738), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G97), .B2(new_n752), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n465), .A2(new_n730), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1203), .B1(new_n814), .B2(new_n745), .C1(new_n206), .C2(new_n741), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1209), .A2(new_n950), .A3(new_n1063), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1207), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT58), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1205), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n1212), .B2(new_n1211), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n757), .A2(new_n1139), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1215), .A2(KEYINPUT115), .B1(new_n742), .B2(G128), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(KEYINPUT115), .B2(new_n1215), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT116), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n731), .A2(new_n946), .B1(new_n937), .B2(new_n1146), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n752), .A2(G132), .B1(G150), .B2(new_n754), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1218), .A2(new_n1219), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1224));
  AOI211_X1 g1024(.A(G33), .B(G41), .C1(new_n746), .C2(G124), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n827), .B2(new_n738), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1223), .B2(KEYINPUT59), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1214), .B1(new_n1224), .B2(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1228), .A2(new_n727), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT117), .Z(new_n1230));
  AOI211_X1 g1030(.A(new_n797), .B(new_n1230), .C1(new_n202), .C2(new_n811), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1185), .A2(new_n787), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1202), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1034), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1200), .A2(new_n1197), .B1(new_n1178), .B2(new_n1175), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1235), .B1(new_n1236), .B2(KEYINPUT57), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1178), .A2(new_n1175), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT57), .B1(new_n1201), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1234), .B1(new_n1237), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(G375));
  NAND2_X1  g1042(.A1(new_n1120), .A2(new_n787), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n777), .B1(G68), .B2(new_n1137), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n758), .A2(new_n827), .B1(new_n202), .B2(new_n753), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G132), .B2(new_n749), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n379), .B1(new_n746), .B2(G128), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n730), .A2(G150), .B1(new_n742), .B2(G137), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n752), .A2(new_n1139), .B1(G58), .B2(new_n737), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n735), .A2(G107), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n741), .A2(new_n814), .B1(new_n589), .B2(new_n745), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(G294), .B2(new_n749), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n752), .A2(G116), .B1(G97), .B2(new_n757), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1251), .A2(new_n1066), .A3(new_n1253), .A4(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n248), .B1(new_n737), .B2(G77), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(KEYINPUT119), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1250), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1244), .B1(new_n1258), .B2(new_n726), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT120), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1177), .A2(new_n776), .B1(new_n1243), .B2(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1169), .A2(KEYINPUT118), .A3(new_n1164), .A4(new_n1172), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1164), .B(new_n1172), .C1(new_n1176), .C2(new_n1119), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT118), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1262), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1177), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1006), .B1(new_n1267), .B2(new_n1164), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1261), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1269), .B(KEYINPUT121), .ZN(G381));
  NOR3_X1   g1070(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1271));
  INV_X1    g1071(.A(G390), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NOR4_X1   g1073(.A1(G381), .A2(G387), .A3(G378), .A4(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1241), .ZN(G407));
  INV_X1    g1075(.A(G378), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n635), .A2(G213), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1241), .A2(new_n1276), .A3(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(G407), .A2(G213), .A3(new_n1279), .ZN(G409));
  AOI22_X1  g1080(.A1(new_n1201), .A2(new_n776), .B1(new_n1232), .B2(new_n1231), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1201), .A2(new_n1238), .A3(KEYINPUT57), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1034), .ZN(new_n1283));
  OAI211_X1 g1083(.A(G378), .B(new_n1281), .C1(new_n1283), .C2(new_n1239), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1236), .A2(new_n1006), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1281), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1276), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1284), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT60), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1289), .B1(new_n1177), .B2(new_n1175), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1266), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT122), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1267), .A2(new_n1292), .A3(KEYINPUT60), .A4(new_n1164), .ZN(new_n1293));
  OAI21_X1  g1093(.A(KEYINPUT122), .B1(new_n1263), .B2(new_n1289), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n1034), .A3(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1261), .B1(new_n1291), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT123), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G384), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(G384), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT123), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1296), .A2(new_n1298), .A3(new_n1300), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1265), .B(new_n1262), .C1(new_n1173), .C2(new_n1289), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1302), .A2(new_n1034), .A3(new_n1293), .A4(new_n1294), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1303), .A2(KEYINPUT123), .A3(new_n1299), .A4(new_n1261), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1301), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1288), .A2(new_n1277), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(KEYINPUT62), .ZN(new_n1307));
  AOI21_X1  g1107(.A(G378), .B1(new_n1281), .B2(new_n1285), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1308), .B1(new_n1241), .B2(G378), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1278), .A2(G2897), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1301), .A2(new_n1304), .A3(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1310), .B1(new_n1301), .B2(new_n1304), .ZN(new_n1312));
  OAI22_X1  g1112(.A1(new_n1309), .A2(new_n1278), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT61), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1278), .B1(new_n1284), .B2(new_n1287), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1315), .A2(new_n1316), .A3(new_n1305), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1307), .A2(new_n1313), .A3(new_n1314), .A4(new_n1317), .ZN(new_n1318));
  OAI211_X1 g1118(.A(new_n965), .B(G390), .C1(new_n1007), .C2(new_n1030), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(KEYINPUT124), .ZN(new_n1320));
  XOR2_X1   g1120(.A(G393), .B(G396), .Z(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(G387), .A2(new_n1272), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1319), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1320), .A2(new_n1323), .A3(new_n1319), .A4(new_n1321), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1318), .A2(new_n1327), .ZN(new_n1328));
  AND4_X1   g1128(.A1(KEYINPUT63), .A2(new_n1288), .A3(new_n1277), .A4(new_n1305), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT63), .B1(new_n1315), .B2(new_n1305), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1325), .A2(new_n1314), .A3(new_n1326), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(new_n1332), .B(KEYINPUT125), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1331), .A2(new_n1333), .A3(new_n1313), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1328), .A2(new_n1334), .ZN(G405));
  NAND3_X1  g1135(.A1(new_n1327), .A2(KEYINPUT126), .A3(new_n1305), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1305), .A2(KEYINPUT126), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1337), .A2(new_n1326), .A3(new_n1325), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1336), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(G375), .A2(new_n1276), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(new_n1284), .ZN(new_n1341));
  XNOR2_X1  g1141(.A(new_n1339), .B(new_n1341), .ZN(G402));
endmodule


